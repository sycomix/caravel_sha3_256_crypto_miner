magic
tech sky130A
magscale 1 2
timestamp 1608616637
<< locali >>
rect 180993 699227 181027 699669
rect 190193 699227 190227 699669
rect 190745 699227 190779 699669
rect 199853 699227 199887 699669
rect 200129 699159 200163 699737
rect 200313 699227 200347 699669
rect 209513 699227 209547 699669
rect 209697 699159 209731 699737
rect 210065 699227 210099 699669
rect 219173 699227 219207 699669
rect 219449 699159 219483 699737
rect 219633 699227 219667 699669
rect 228833 699227 228867 699669
rect 229017 699159 229051 699737
rect 229385 699227 229419 699669
rect 233249 699227 233283 699941
rect 241437 699771 241471 701641
rect 292221 700077 292531 700111
rect 277961 699771 277995 699805
rect 277961 699737 278145 699771
rect 292221 699703 292255 700077
rect 292497 700043 292531 700077
rect 292405 699703 292439 700009
rect 306389 699941 306883 699975
rect 301973 699873 302157 699907
rect 301973 699703 302007 699873
rect 306389 699771 306423 699941
rect 306849 699907 306883 699941
rect 292405 699669 292497 699703
rect 292589 699669 292773 699703
rect 292589 699431 292623 699669
rect 302065 699431 302099 699669
rect 306481 699227 306515 699669
rect 239321 699193 239505 699227
rect 239321 699159 239355 699193
rect 264989 699159 265023 699193
rect 264989 699125 265173 699159
rect 306389 698887 306423 699193
rect 306665 699159 306699 699669
rect 306757 699159 306791 699873
rect 318809 699703 318843 699873
rect 321511 699737 321569 699771
rect 325341 699227 325375 699669
rect 325433 699159 325467 699873
rect 331229 699839 331263 700213
rect 336013 699771 336047 700213
rect 338129 699771 338163 700213
rect 347697 699839 347731 700213
rect 325985 699227 326019 699669
rect 354321 699227 354355 699669
rect 325617 698887 325651 699193
rect 354413 699159 354447 699737
rect 354781 699431 354815 699669
rect 364165 699431 364199 699669
rect 364257 699431 364291 699737
rect 373733 699737 373951 699771
rect 373733 699703 373767 699737
rect 373825 699499 373859 699669
rect 373917 699499 373951 699737
rect 340739 699125 340831 699159
rect 306389 698853 306481 698887
rect 325559 698853 325651 698887
rect 340797 698887 340831 699125
rect 354597 698887 354631 699193
rect 354539 698853 354631 698887
rect 354689 698275 354723 699397
rect 6193 696643 6227 696745
rect 86969 696439 87003 696609
rect 22201 696371 22235 696405
rect 60841 696371 60875 696405
rect 22051 696337 22235 696371
rect 60691 696337 60875 696371
rect 6101 693379 6135 696337
rect 67649 696235 67683 696405
rect 80161 696371 80195 696405
rect 80011 696337 80195 696371
rect 96537 696371 96571 696609
rect 99389 696371 99423 696405
rect 99331 696337 99423 696371
rect 77217 696235 77251 696337
rect 108957 696303 108991 696405
rect 115857 696303 115891 696405
rect 143583 696337 143675 696371
rect 132509 696099 132543 696269
rect 138121 696099 138155 696337
rect 143641 696303 143675 696337
rect 154589 696303 154623 696473
rect 163881 696303 163915 696473
rect 164099 696405 164249 696439
rect 154715 696201 154773 696235
rect 154623 696133 154957 696167
rect 154715 696065 154865 696099
rect 17233 695555 17267 695657
rect 31769 695555 31803 695657
rect 46213 695555 46247 695997
rect 55873 695691 55907 695997
rect 62773 695691 62807 695997
rect 75193 695691 75227 695997
rect 82093 695691 82127 695997
rect 94513 695691 94547 695997
rect 123987 695997 124079 696031
rect 57805 695317 58023 695351
rect 57805 695147 57839 695317
rect 9689 694671 9723 694773
rect 19257 694671 19291 694841
rect 28825 694807 28859 694841
rect 28825 694773 28917 694807
rect 44189 694603 44223 694773
rect 53757 694603 53791 694705
rect 57897 694195 57931 695249
rect 57989 695215 58023 695317
rect 67465 694331 67499 695249
rect 75963 695181 76055 695215
rect 76021 695079 76055 695181
rect 75929 694671 75963 694773
rect 81357 694399 81391 695249
rect 95283 694909 95433 694943
rect 86969 694739 87003 694841
rect 86911 694705 87003 694739
rect 95801 694535 95835 695249
rect 98043 694841 98135 694875
rect 98101 694807 98135 694841
rect 100585 694603 100619 695249
rect 104909 694875 104943 695181
rect 106323 694773 106381 694807
rect 109969 694671 110003 695249
rect 114477 694875 114511 695113
rect 114569 694807 114603 695997
rect 114661 694875 114695 695113
rect 117237 694875 117271 695181
rect 110279 694773 110337 694807
rect 124045 694807 124079 695997
rect 124137 694875 124171 695997
rect 124355 695181 124447 695215
rect 124413 695147 124447 695181
rect 128311 695113 128369 695147
rect 138489 694875 138523 695997
rect 154715 695929 154865 695963
rect 154623 695793 155049 695827
rect 154715 695725 154957 695759
rect 154623 695657 154865 695691
rect 154623 695521 154865 695555
rect 125333 694807 125367 694841
rect 125609 694807 125643 694841
rect 124045 694773 124171 694807
rect 125333 694773 125517 694807
rect 125609 694773 125793 694807
rect 124137 694739 124171 694773
rect 125885 694739 125919 694841
rect 125735 694705 125919 694739
rect 137293 694739 137327 694841
rect 138247 694773 138397 694807
rect 147689 694739 147723 695113
rect 154589 695079 154623 695249
rect 156981 694739 157015 695113
rect 157441 695079 157475 695249
rect 167009 694739 167043 695249
rect 171609 695147 171643 696337
rect 173909 696303 173943 696473
rect 178693 696371 178727 696473
rect 186329 696371 186363 696473
rect 200715 696405 200865 696439
rect 205649 696371 205683 696609
rect 215217 696371 215251 696609
rect 224969 696371 225003 696881
rect 234537 696371 234571 696881
rect 244289 696371 244323 696881
rect 253857 696371 253891 696881
rect 263609 696371 263643 696881
rect 273177 696371 273211 696881
rect 282929 696371 282963 696881
rect 292497 696371 292531 696881
rect 174035 696201 174093 696235
rect 174035 696065 174185 696099
rect 174035 695929 174185 695963
rect 173943 695861 174277 695895
rect 297281 695691 297315 696881
rect 297373 696371 297407 696813
rect 174035 695657 174185 695691
rect 306941 695691 306975 696881
rect 307033 696371 307067 696813
rect 355241 695691 355275 696881
rect 355333 696371 355367 696813
rect 362141 695691 362175 696881
rect 364993 696371 365027 696813
rect 372261 696371 372295 696677
rect 374653 695691 374687 696813
rect 384313 695691 384347 696813
rect 393973 695691 394007 696337
rect 403633 695691 403667 696337
rect 567025 696167 567059 696269
rect 413293 695691 413327 696133
rect 422953 695691 422987 696133
rect 432337 695691 432371 696133
rect 442273 695691 442307 696133
rect 451289 695691 451323 695929
rect 461409 695691 461443 695929
rect 471253 695691 471287 695861
rect 483029 695827 483063 695929
rect 492597 695759 492631 695929
rect 492689 695691 492723 695929
rect 502257 695691 502291 695929
rect 173943 695589 174093 695623
rect 174035 695521 174185 695555
rect 125643 694501 125885 694535
rect 125735 694365 125793 694399
rect 125643 694297 125885 694331
rect 171517 694127 171551 695113
rect 176485 694127 176519 695181
rect 176577 694739 176611 695249
rect 186329 694739 186363 695249
rect 195897 694739 195931 695249
rect 355609 694739 355643 695453
rect 205649 694127 205683 694705
rect 215217 694127 215251 694705
rect 224969 694127 225003 694705
rect 234537 694127 234571 694705
rect 244289 694127 244323 694705
rect 253857 694127 253891 694705
rect 263609 694127 263643 694705
rect 273177 694127 273211 694705
rect 282929 694127 282963 694705
rect 292497 694127 292531 694705
rect 302157 694127 302191 694705
rect 364993 694739 365027 695453
rect 374653 694739 374687 695385
rect 384313 694739 384347 695385
rect 393973 694739 394007 695317
rect 403633 694739 403667 695317
rect 413293 694739 413327 695317
rect 422953 694739 422987 695317
rect 426541 695011 426575 695317
rect 432613 694739 432647 694977
rect 440709 694943 440743 695317
rect 441905 694739 441939 694977
rect 451289 694739 451323 694909
rect 461593 694739 461627 694909
rect 469229 694739 469263 695317
rect 302249 694127 302283 694705
rect 497565 694467 497599 695317
rect 511917 694263 511951 695317
<< viali >>
rect 241437 701641 241471 701675
rect 233249 699941 233283 699975
rect 200129 699737 200163 699771
rect 180993 699669 181027 699703
rect 180993 699193 181027 699227
rect 190193 699669 190227 699703
rect 190193 699193 190227 699227
rect 190745 699669 190779 699703
rect 190745 699193 190779 699227
rect 199853 699669 199887 699703
rect 199853 699193 199887 699227
rect 209697 699737 209731 699771
rect 200313 699669 200347 699703
rect 200313 699193 200347 699227
rect 209513 699669 209547 699703
rect 209513 699193 209547 699227
rect 200129 699125 200163 699159
rect 219449 699737 219483 699771
rect 210065 699669 210099 699703
rect 210065 699193 210099 699227
rect 219173 699669 219207 699703
rect 219173 699193 219207 699227
rect 209697 699125 209731 699159
rect 229017 699737 229051 699771
rect 219633 699669 219667 699703
rect 219633 699193 219667 699227
rect 228833 699669 228867 699703
rect 228833 699193 228867 699227
rect 219449 699125 219483 699159
rect 229385 699669 229419 699703
rect 229385 699193 229419 699227
rect 331229 700213 331263 700247
rect 241437 699737 241471 699771
rect 277961 699805 277995 699839
rect 278145 699737 278179 699771
rect 292221 699669 292255 699703
rect 292405 700009 292439 700043
rect 292497 700009 292531 700043
rect 302157 699873 302191 699907
rect 306389 699737 306423 699771
rect 306757 699873 306791 699907
rect 306849 699873 306883 699907
rect 318809 699873 318843 699907
rect 292497 699669 292531 699703
rect 292773 699669 292807 699703
rect 301973 699669 302007 699703
rect 302065 699669 302099 699703
rect 292589 699397 292623 699431
rect 302065 699397 302099 699431
rect 306481 699669 306515 699703
rect 233249 699193 233283 699227
rect 239505 699193 239539 699227
rect 264989 699193 265023 699227
rect 229017 699125 229051 699159
rect 239321 699125 239355 699159
rect 306389 699193 306423 699227
rect 306481 699193 306515 699227
rect 306665 699669 306699 699703
rect 265173 699125 265207 699159
rect 306665 699125 306699 699159
rect 325433 699873 325467 699907
rect 321477 699737 321511 699771
rect 321569 699737 321603 699771
rect 318809 699669 318843 699703
rect 325341 699669 325375 699703
rect 325341 699193 325375 699227
rect 306757 699125 306791 699159
rect 331229 699805 331263 699839
rect 336013 700213 336047 700247
rect 336013 699737 336047 699771
rect 338129 700213 338163 700247
rect 347697 700213 347731 700247
rect 347697 699805 347731 699839
rect 338129 699737 338163 699771
rect 354413 699737 354447 699771
rect 325985 699669 326019 699703
rect 325433 699125 325467 699159
rect 325617 699193 325651 699227
rect 325985 699193 326019 699227
rect 354321 699669 354355 699703
rect 354321 699193 354355 699227
rect 364257 699737 364291 699771
rect 354781 699669 354815 699703
rect 354689 699397 354723 699431
rect 354781 699397 354815 699431
rect 364165 699669 364199 699703
rect 364165 699397 364199 699431
rect 373733 699669 373767 699703
rect 373825 699669 373859 699703
rect 373825 699465 373859 699499
rect 373917 699465 373951 699499
rect 364257 699397 364291 699431
rect 340705 699125 340739 699159
rect 354413 699125 354447 699159
rect 354597 699193 354631 699227
rect 306481 698853 306515 698887
rect 325525 698853 325559 698887
rect 340797 698853 340831 698887
rect 354505 698853 354539 698887
rect 354689 698241 354723 698275
rect 224969 696881 225003 696915
rect 6193 696745 6227 696779
rect 6193 696609 6227 696643
rect 86969 696609 87003 696643
rect 22201 696405 22235 696439
rect 60841 696405 60875 696439
rect 6101 696337 6135 696371
rect 22017 696337 22051 696371
rect 60657 696337 60691 696371
rect 67649 696405 67683 696439
rect 80161 696405 80195 696439
rect 86969 696405 87003 696439
rect 96537 696609 96571 696643
rect 67649 696201 67683 696235
rect 77217 696337 77251 696371
rect 79977 696337 80011 696371
rect 205649 696609 205683 696643
rect 154589 696473 154623 696507
rect 99389 696405 99423 696439
rect 96537 696337 96571 696371
rect 99297 696337 99331 696371
rect 108957 696405 108991 696439
rect 108957 696269 108991 696303
rect 115857 696405 115891 696439
rect 138121 696337 138155 696371
rect 143549 696337 143583 696371
rect 115857 696269 115891 696303
rect 132509 696269 132543 696303
rect 77217 696201 77251 696235
rect 132509 696065 132543 696099
rect 143641 696269 143675 696303
rect 154589 696269 154623 696303
rect 163881 696473 163915 696507
rect 173909 696473 173943 696507
rect 164065 696405 164099 696439
rect 164249 696405 164283 696439
rect 163881 696269 163915 696303
rect 171609 696337 171643 696371
rect 154681 696201 154715 696235
rect 154773 696201 154807 696235
rect 154589 696133 154623 696167
rect 154957 696133 154991 696167
rect 138121 696065 138155 696099
rect 154681 696065 154715 696099
rect 154865 696065 154899 696099
rect 46213 695997 46247 696031
rect 17233 695657 17267 695691
rect 17233 695521 17267 695555
rect 31769 695657 31803 695691
rect 31769 695521 31803 695555
rect 55873 695997 55907 696031
rect 55873 695657 55907 695691
rect 62773 695997 62807 696031
rect 62773 695657 62807 695691
rect 75193 695997 75227 696031
rect 75193 695657 75227 695691
rect 82093 695997 82127 696031
rect 82093 695657 82127 695691
rect 94513 695997 94547 696031
rect 94513 695657 94547 695691
rect 114569 695997 114603 696031
rect 123953 695997 123987 696031
rect 46213 695521 46247 695555
rect 57805 695113 57839 695147
rect 57897 695249 57931 695283
rect 19257 694841 19291 694875
rect 9689 694773 9723 694807
rect 9689 694637 9723 694671
rect 28825 694841 28859 694875
rect 28917 694773 28951 694807
rect 44189 694773 44223 694807
rect 19257 694637 19291 694671
rect 44189 694569 44223 694603
rect 53757 694705 53791 694739
rect 53757 694569 53791 694603
rect 57989 695181 58023 695215
rect 67465 695249 67499 695283
rect 81357 695249 81391 695283
rect 75929 695181 75963 695215
rect 76021 695045 76055 695079
rect 75929 694773 75963 694807
rect 75929 694637 75963 694671
rect 95801 695249 95835 695283
rect 95249 694909 95283 694943
rect 95433 694909 95467 694943
rect 86969 694841 87003 694875
rect 86877 694705 86911 694739
rect 100585 695249 100619 695283
rect 98009 694841 98043 694875
rect 98101 694773 98135 694807
rect 109969 695249 110003 695283
rect 104909 695181 104943 695215
rect 104909 694841 104943 694875
rect 106289 694773 106323 694807
rect 106381 694773 106415 694807
rect 114477 695113 114511 695147
rect 114477 694841 114511 694875
rect 117237 695181 117271 695215
rect 114661 695113 114695 695147
rect 114661 694841 114695 694875
rect 117237 694841 117271 694875
rect 110245 694773 110279 694807
rect 110337 694773 110371 694807
rect 114569 694773 114603 694807
rect 124137 695997 124171 696031
rect 138489 695997 138523 696031
rect 124321 695181 124355 695215
rect 124413 695113 124447 695147
rect 128277 695113 128311 695147
rect 128369 695113 128403 695147
rect 154681 695929 154715 695963
rect 154865 695929 154899 695963
rect 154589 695793 154623 695827
rect 155049 695793 155083 695827
rect 154681 695725 154715 695759
rect 154957 695725 154991 695759
rect 154589 695657 154623 695691
rect 154865 695657 154899 695691
rect 154589 695521 154623 695555
rect 154865 695521 154899 695555
rect 154589 695249 154623 695283
rect 124137 694841 124171 694875
rect 125333 694841 125367 694875
rect 125609 694841 125643 694875
rect 125885 694841 125919 694875
rect 125517 694773 125551 694807
rect 125793 694773 125827 694807
rect 124137 694705 124171 694739
rect 125701 694705 125735 694739
rect 137293 694841 137327 694875
rect 138489 694841 138523 694875
rect 147689 695113 147723 695147
rect 138213 694773 138247 694807
rect 138397 694773 138431 694807
rect 137293 694705 137327 694739
rect 157441 695249 157475 695283
rect 154589 695045 154623 695079
rect 156981 695113 157015 695147
rect 147689 694705 147723 694739
rect 157441 695045 157475 695079
rect 167009 695249 167043 695283
rect 156981 694705 157015 694739
rect 178693 696473 178727 696507
rect 178693 696337 178727 696371
rect 186329 696473 186363 696507
rect 200681 696405 200715 696439
rect 200865 696405 200899 696439
rect 186329 696337 186363 696371
rect 205649 696337 205683 696371
rect 215217 696609 215251 696643
rect 215217 696337 215251 696371
rect 224969 696337 225003 696371
rect 234537 696881 234571 696915
rect 234537 696337 234571 696371
rect 244289 696881 244323 696915
rect 244289 696337 244323 696371
rect 253857 696881 253891 696915
rect 253857 696337 253891 696371
rect 263609 696881 263643 696915
rect 263609 696337 263643 696371
rect 273177 696881 273211 696915
rect 273177 696337 273211 696371
rect 282929 696881 282963 696915
rect 282929 696337 282963 696371
rect 292497 696881 292531 696915
rect 292497 696337 292531 696371
rect 297281 696881 297315 696915
rect 173909 696269 173943 696303
rect 174001 696201 174035 696235
rect 174093 696201 174127 696235
rect 174001 696065 174035 696099
rect 174185 696065 174219 696099
rect 174001 695929 174035 695963
rect 174185 695929 174219 695963
rect 173909 695861 173943 695895
rect 174277 695861 174311 695895
rect 306941 696881 306975 696915
rect 297373 696813 297407 696847
rect 297373 696337 297407 696371
rect 174001 695657 174035 695691
rect 174185 695657 174219 695691
rect 297281 695657 297315 695691
rect 355241 696881 355275 696915
rect 307033 696813 307067 696847
rect 307033 696337 307067 696371
rect 306941 695657 306975 695691
rect 362141 696881 362175 696915
rect 355333 696813 355367 696847
rect 355333 696337 355367 696371
rect 355241 695657 355275 695691
rect 364993 696813 365027 696847
rect 374653 696813 374687 696847
rect 364993 696337 365027 696371
rect 372261 696677 372295 696711
rect 372261 696337 372295 696371
rect 362141 695657 362175 695691
rect 374653 695657 374687 695691
rect 384313 696813 384347 696847
rect 384313 695657 384347 695691
rect 393973 696337 394007 696371
rect 393973 695657 394007 695691
rect 403633 696337 403667 696371
rect 567025 696269 567059 696303
rect 403633 695657 403667 695691
rect 413293 696133 413327 696167
rect 413293 695657 413327 695691
rect 422953 696133 422987 696167
rect 422953 695657 422987 695691
rect 432337 696133 432371 696167
rect 432337 695657 432371 695691
rect 442273 696133 442307 696167
rect 567025 696133 567059 696167
rect 442273 695657 442307 695691
rect 451289 695929 451323 695963
rect 451289 695657 451323 695691
rect 461409 695929 461443 695963
rect 483029 695929 483063 695963
rect 461409 695657 461443 695691
rect 471253 695861 471287 695895
rect 483029 695793 483063 695827
rect 492597 695929 492631 695963
rect 492597 695725 492631 695759
rect 492689 695929 492723 695963
rect 471253 695657 471287 695691
rect 492689 695657 492723 695691
rect 502257 695929 502291 695963
rect 502257 695657 502291 695691
rect 173909 695589 173943 695623
rect 174093 695589 174127 695623
rect 174001 695521 174035 695555
rect 174185 695521 174219 695555
rect 355609 695453 355643 695487
rect 176577 695249 176611 695283
rect 167009 694705 167043 694739
rect 171517 695113 171551 695147
rect 171609 695113 171643 695147
rect 176485 695181 176519 695215
rect 109969 694637 110003 694671
rect 100585 694569 100619 694603
rect 95801 694501 95835 694535
rect 125609 694501 125643 694535
rect 125885 694501 125919 694535
rect 81357 694365 81391 694399
rect 125701 694365 125735 694399
rect 125793 694365 125827 694399
rect 67465 694297 67499 694331
rect 125609 694297 125643 694331
rect 125885 694297 125919 694331
rect 57897 694161 57931 694195
rect 171517 694093 171551 694127
rect 176577 694705 176611 694739
rect 186329 695249 186363 695283
rect 186329 694705 186363 694739
rect 195897 695249 195931 695283
rect 195897 694705 195931 694739
rect 205649 694705 205683 694739
rect 176485 694093 176519 694127
rect 205649 694093 205683 694127
rect 215217 694705 215251 694739
rect 215217 694093 215251 694127
rect 224969 694705 225003 694739
rect 224969 694093 225003 694127
rect 234537 694705 234571 694739
rect 234537 694093 234571 694127
rect 244289 694705 244323 694739
rect 244289 694093 244323 694127
rect 253857 694705 253891 694739
rect 253857 694093 253891 694127
rect 263609 694705 263643 694739
rect 263609 694093 263643 694127
rect 273177 694705 273211 694739
rect 273177 694093 273211 694127
rect 282929 694705 282963 694739
rect 282929 694093 282963 694127
rect 292497 694705 292531 694739
rect 292497 694093 292531 694127
rect 302157 694705 302191 694739
rect 302157 694093 302191 694127
rect 302249 694705 302283 694739
rect 355609 694705 355643 694739
rect 364993 695453 365027 695487
rect 364993 694705 365027 694739
rect 374653 695385 374687 695419
rect 374653 694705 374687 694739
rect 384313 695385 384347 695419
rect 384313 694705 384347 694739
rect 393973 695317 394007 695351
rect 393973 694705 394007 694739
rect 403633 695317 403667 695351
rect 403633 694705 403667 694739
rect 413293 695317 413327 695351
rect 413293 694705 413327 694739
rect 422953 695317 422987 695351
rect 426541 695317 426575 695351
rect 440709 695317 440743 695351
rect 426541 694977 426575 695011
rect 432613 694977 432647 695011
rect 422953 694705 422987 694739
rect 469229 695317 469263 695351
rect 440709 694909 440743 694943
rect 441905 694977 441939 695011
rect 432613 694705 432647 694739
rect 441905 694705 441939 694739
rect 451289 694909 451323 694943
rect 451289 694705 451323 694739
rect 461593 694909 461627 694943
rect 461593 694705 461627 694739
rect 469229 694705 469263 694739
rect 497565 695317 497599 695351
rect 497565 694433 497599 694467
rect 511917 695317 511951 695351
rect 511917 694229 511951 694263
rect 302249 694093 302283 694127
rect 6101 693345 6135 693379
<< metal1 >>
rect 251634 701972 251640 702024
rect 251692 702012 251698 702024
rect 429838 702012 429844 702024
rect 251692 701984 429844 702012
rect 251692 701972 251698 701984
rect 429838 701972 429844 701984
rect 429896 701972 429902 702024
rect 237466 701904 237472 701956
rect 237524 701944 237530 701956
rect 494790 701944 494796 701956
rect 237524 701916 494796 701944
rect 237524 701904 237530 701916
rect 494790 701904 494796 701916
rect 494848 701904 494854 701956
rect 223298 701836 223304 701888
rect 223356 701876 223362 701888
rect 559650 701876 559656 701888
rect 223356 701848 559656 701876
rect 223356 701836 223362 701848
rect 559650 701836 559656 701848
rect 559708 701836 559714 701888
rect 1104 701786 582820 701808
rect 1104 701734 36822 701786
rect 36874 701734 36886 701786
rect 36938 701734 36950 701786
rect 37002 701734 37014 701786
rect 37066 701734 37078 701786
rect 37130 701734 37142 701786
rect 37194 701734 37206 701786
rect 37258 701734 37270 701786
rect 37322 701734 37334 701786
rect 37386 701734 72822 701786
rect 72874 701734 72886 701786
rect 72938 701734 72950 701786
rect 73002 701734 73014 701786
rect 73066 701734 73078 701786
rect 73130 701734 73142 701786
rect 73194 701734 73206 701786
rect 73258 701734 73270 701786
rect 73322 701734 73334 701786
rect 73386 701734 108822 701786
rect 108874 701734 108886 701786
rect 108938 701734 108950 701786
rect 109002 701734 109014 701786
rect 109066 701734 109078 701786
rect 109130 701734 109142 701786
rect 109194 701734 109206 701786
rect 109258 701734 109270 701786
rect 109322 701734 109334 701786
rect 109386 701734 144822 701786
rect 144874 701734 144886 701786
rect 144938 701734 144950 701786
rect 145002 701734 145014 701786
rect 145066 701734 145078 701786
rect 145130 701734 145142 701786
rect 145194 701734 145206 701786
rect 145258 701734 145270 701786
rect 145322 701734 145334 701786
rect 145386 701734 180822 701786
rect 180874 701734 180886 701786
rect 180938 701734 180950 701786
rect 181002 701734 181014 701786
rect 181066 701734 181078 701786
rect 181130 701734 181142 701786
rect 181194 701734 181206 701786
rect 181258 701734 181270 701786
rect 181322 701734 181334 701786
rect 181386 701734 216822 701786
rect 216874 701734 216886 701786
rect 216938 701734 216950 701786
rect 217002 701734 217014 701786
rect 217066 701734 217078 701786
rect 217130 701734 217142 701786
rect 217194 701734 217206 701786
rect 217258 701734 217270 701786
rect 217322 701734 217334 701786
rect 217386 701734 252822 701786
rect 252874 701734 252886 701786
rect 252938 701734 252950 701786
rect 253002 701734 253014 701786
rect 253066 701734 253078 701786
rect 253130 701734 253142 701786
rect 253194 701734 253206 701786
rect 253258 701734 253270 701786
rect 253322 701734 253334 701786
rect 253386 701734 288822 701786
rect 288874 701734 288886 701786
rect 288938 701734 288950 701786
rect 289002 701734 289014 701786
rect 289066 701734 289078 701786
rect 289130 701734 289142 701786
rect 289194 701734 289206 701786
rect 289258 701734 289270 701786
rect 289322 701734 289334 701786
rect 289386 701734 324822 701786
rect 324874 701734 324886 701786
rect 324938 701734 324950 701786
rect 325002 701734 325014 701786
rect 325066 701734 325078 701786
rect 325130 701734 325142 701786
rect 325194 701734 325206 701786
rect 325258 701734 325270 701786
rect 325322 701734 325334 701786
rect 325386 701734 360822 701786
rect 360874 701734 360886 701786
rect 360938 701734 360950 701786
rect 361002 701734 361014 701786
rect 361066 701734 361078 701786
rect 361130 701734 361142 701786
rect 361194 701734 361206 701786
rect 361258 701734 361270 701786
rect 361322 701734 361334 701786
rect 361386 701734 396822 701786
rect 396874 701734 396886 701786
rect 396938 701734 396950 701786
rect 397002 701734 397014 701786
rect 397066 701734 397078 701786
rect 397130 701734 397142 701786
rect 397194 701734 397206 701786
rect 397258 701734 397270 701786
rect 397322 701734 397334 701786
rect 397386 701734 432822 701786
rect 432874 701734 432886 701786
rect 432938 701734 432950 701786
rect 433002 701734 433014 701786
rect 433066 701734 433078 701786
rect 433130 701734 433142 701786
rect 433194 701734 433206 701786
rect 433258 701734 433270 701786
rect 433322 701734 433334 701786
rect 433386 701734 468822 701786
rect 468874 701734 468886 701786
rect 468938 701734 468950 701786
rect 469002 701734 469014 701786
rect 469066 701734 469078 701786
rect 469130 701734 469142 701786
rect 469194 701734 469206 701786
rect 469258 701734 469270 701786
rect 469322 701734 469334 701786
rect 469386 701734 504822 701786
rect 504874 701734 504886 701786
rect 504938 701734 504950 701786
rect 505002 701734 505014 701786
rect 505066 701734 505078 701786
rect 505130 701734 505142 701786
rect 505194 701734 505206 701786
rect 505258 701734 505270 701786
rect 505322 701734 505334 701786
rect 505386 701734 540822 701786
rect 540874 701734 540886 701786
rect 540938 701734 540950 701786
rect 541002 701734 541014 701786
rect 541066 701734 541078 701786
rect 541130 701734 541142 701786
rect 541194 701734 541206 701786
rect 541258 701734 541270 701786
rect 541322 701734 541334 701786
rect 541386 701734 576822 701786
rect 576874 701734 576886 701786
rect 576938 701734 576950 701786
rect 577002 701734 577014 701786
rect 577066 701734 577078 701786
rect 577130 701734 577142 701786
rect 577194 701734 577206 701786
rect 577258 701734 577270 701786
rect 577322 701734 577334 701786
rect 577386 701734 582820 701786
rect 1104 701712 582820 701734
rect 235166 701632 235172 701684
rect 235224 701672 235230 701684
rect 241425 701675 241483 701681
rect 241425 701672 241437 701675
rect 235224 701644 241437 701672
rect 235224 701632 235230 701644
rect 241425 701641 241437 701644
rect 241471 701641 241483 701675
rect 241425 701635 241483 701641
rect 1104 701242 582820 701264
rect 1104 701190 18822 701242
rect 18874 701190 18886 701242
rect 18938 701190 18950 701242
rect 19002 701190 19014 701242
rect 19066 701190 19078 701242
rect 19130 701190 19142 701242
rect 19194 701190 19206 701242
rect 19258 701190 19270 701242
rect 19322 701190 19334 701242
rect 19386 701190 54822 701242
rect 54874 701190 54886 701242
rect 54938 701190 54950 701242
rect 55002 701190 55014 701242
rect 55066 701190 55078 701242
rect 55130 701190 55142 701242
rect 55194 701190 55206 701242
rect 55258 701190 55270 701242
rect 55322 701190 55334 701242
rect 55386 701190 90822 701242
rect 90874 701190 90886 701242
rect 90938 701190 90950 701242
rect 91002 701190 91014 701242
rect 91066 701190 91078 701242
rect 91130 701190 91142 701242
rect 91194 701190 91206 701242
rect 91258 701190 91270 701242
rect 91322 701190 91334 701242
rect 91386 701190 126822 701242
rect 126874 701190 126886 701242
rect 126938 701190 126950 701242
rect 127002 701190 127014 701242
rect 127066 701190 127078 701242
rect 127130 701190 127142 701242
rect 127194 701190 127206 701242
rect 127258 701190 127270 701242
rect 127322 701190 127334 701242
rect 127386 701190 162822 701242
rect 162874 701190 162886 701242
rect 162938 701190 162950 701242
rect 163002 701190 163014 701242
rect 163066 701190 163078 701242
rect 163130 701190 163142 701242
rect 163194 701190 163206 701242
rect 163258 701190 163270 701242
rect 163322 701190 163334 701242
rect 163386 701190 198822 701242
rect 198874 701190 198886 701242
rect 198938 701190 198950 701242
rect 199002 701190 199014 701242
rect 199066 701190 199078 701242
rect 199130 701190 199142 701242
rect 199194 701190 199206 701242
rect 199258 701190 199270 701242
rect 199322 701190 199334 701242
rect 199386 701190 234822 701242
rect 234874 701190 234886 701242
rect 234938 701190 234950 701242
rect 235002 701190 235014 701242
rect 235066 701190 235078 701242
rect 235130 701190 235142 701242
rect 235194 701190 235206 701242
rect 235258 701190 235270 701242
rect 235322 701190 235334 701242
rect 235386 701190 270822 701242
rect 270874 701190 270886 701242
rect 270938 701190 270950 701242
rect 271002 701190 271014 701242
rect 271066 701190 271078 701242
rect 271130 701190 271142 701242
rect 271194 701190 271206 701242
rect 271258 701190 271270 701242
rect 271322 701190 271334 701242
rect 271386 701190 306822 701242
rect 306874 701190 306886 701242
rect 306938 701190 306950 701242
rect 307002 701190 307014 701242
rect 307066 701190 307078 701242
rect 307130 701190 307142 701242
rect 307194 701190 307206 701242
rect 307258 701190 307270 701242
rect 307322 701190 307334 701242
rect 307386 701190 342822 701242
rect 342874 701190 342886 701242
rect 342938 701190 342950 701242
rect 343002 701190 343014 701242
rect 343066 701190 343078 701242
rect 343130 701190 343142 701242
rect 343194 701190 343206 701242
rect 343258 701190 343270 701242
rect 343322 701190 343334 701242
rect 343386 701190 378822 701242
rect 378874 701190 378886 701242
rect 378938 701190 378950 701242
rect 379002 701190 379014 701242
rect 379066 701190 379078 701242
rect 379130 701190 379142 701242
rect 379194 701190 379206 701242
rect 379258 701190 379270 701242
rect 379322 701190 379334 701242
rect 379386 701190 414822 701242
rect 414874 701190 414886 701242
rect 414938 701190 414950 701242
rect 415002 701190 415014 701242
rect 415066 701190 415078 701242
rect 415130 701190 415142 701242
rect 415194 701190 415206 701242
rect 415258 701190 415270 701242
rect 415322 701190 415334 701242
rect 415386 701190 450822 701242
rect 450874 701190 450886 701242
rect 450938 701190 450950 701242
rect 451002 701190 451014 701242
rect 451066 701190 451078 701242
rect 451130 701190 451142 701242
rect 451194 701190 451206 701242
rect 451258 701190 451270 701242
rect 451322 701190 451334 701242
rect 451386 701190 486822 701242
rect 486874 701190 486886 701242
rect 486938 701190 486950 701242
rect 487002 701190 487014 701242
rect 487066 701190 487078 701242
rect 487130 701190 487142 701242
rect 487194 701190 487206 701242
rect 487258 701190 487270 701242
rect 487322 701190 487334 701242
rect 487386 701190 522822 701242
rect 522874 701190 522886 701242
rect 522938 701190 522950 701242
rect 523002 701190 523014 701242
rect 523066 701190 523078 701242
rect 523130 701190 523142 701242
rect 523194 701190 523206 701242
rect 523258 701190 523270 701242
rect 523322 701190 523334 701242
rect 523386 701190 558822 701242
rect 558874 701190 558886 701242
rect 558938 701190 558950 701242
rect 559002 701190 559014 701242
rect 559066 701190 559078 701242
rect 559130 701190 559142 701242
rect 559194 701190 559206 701242
rect 559258 701190 559270 701242
rect 559322 701190 559334 701242
rect 559386 701190 582820 701242
rect 1104 701168 582820 701190
rect 256418 700952 256424 701004
rect 256476 700992 256482 701004
rect 397454 700992 397460 701004
rect 256476 700964 397460 700992
rect 256476 700952 256482 700964
rect 397454 700952 397460 700964
rect 397512 700952 397518 701004
rect 154114 700884 154120 700936
rect 154172 700924 154178 700936
rect 317966 700924 317972 700936
rect 154172 700896 317972 700924
rect 154172 700884 154178 700896
rect 317966 700884 317972 700896
rect 318024 700884 318030 700936
rect 137830 700816 137836 700868
rect 137888 700856 137894 700868
rect 313182 700856 313188 700868
rect 137888 700828 313188 700856
rect 137888 700816 137894 700828
rect 313182 700816 313188 700828
rect 313240 700816 313246 700868
rect 105446 700748 105452 700800
rect 105504 700788 105510 700800
rect 322658 700788 322664 700800
rect 105504 700760 322664 700788
rect 105504 700748 105510 700760
rect 322658 700748 322664 700760
rect 322716 700748 322722 700800
rect 1104 700698 582820 700720
rect 1104 700646 36822 700698
rect 36874 700646 36886 700698
rect 36938 700646 36950 700698
rect 37002 700646 37014 700698
rect 37066 700646 37078 700698
rect 37130 700646 37142 700698
rect 37194 700646 37206 700698
rect 37258 700646 37270 700698
rect 37322 700646 37334 700698
rect 37386 700646 72822 700698
rect 72874 700646 72886 700698
rect 72938 700646 72950 700698
rect 73002 700646 73014 700698
rect 73066 700646 73078 700698
rect 73130 700646 73142 700698
rect 73194 700646 73206 700698
rect 73258 700646 73270 700698
rect 73322 700646 73334 700698
rect 73386 700646 108822 700698
rect 108874 700646 108886 700698
rect 108938 700646 108950 700698
rect 109002 700646 109014 700698
rect 109066 700646 109078 700698
rect 109130 700646 109142 700698
rect 109194 700646 109206 700698
rect 109258 700646 109270 700698
rect 109322 700646 109334 700698
rect 109386 700646 144822 700698
rect 144874 700646 144886 700698
rect 144938 700646 144950 700698
rect 145002 700646 145014 700698
rect 145066 700646 145078 700698
rect 145130 700646 145142 700698
rect 145194 700646 145206 700698
rect 145258 700646 145270 700698
rect 145322 700646 145334 700698
rect 145386 700646 180822 700698
rect 180874 700646 180886 700698
rect 180938 700646 180950 700698
rect 181002 700646 181014 700698
rect 181066 700646 181078 700698
rect 181130 700646 181142 700698
rect 181194 700646 181206 700698
rect 181258 700646 181270 700698
rect 181322 700646 181334 700698
rect 181386 700646 216822 700698
rect 216874 700646 216886 700698
rect 216938 700646 216950 700698
rect 217002 700646 217014 700698
rect 217066 700646 217078 700698
rect 217130 700646 217142 700698
rect 217194 700646 217206 700698
rect 217258 700646 217270 700698
rect 217322 700646 217334 700698
rect 217386 700646 252822 700698
rect 252874 700646 252886 700698
rect 252938 700646 252950 700698
rect 253002 700646 253014 700698
rect 253066 700646 253078 700698
rect 253130 700646 253142 700698
rect 253194 700646 253206 700698
rect 253258 700646 253270 700698
rect 253322 700646 253334 700698
rect 253386 700646 288822 700698
rect 288874 700646 288886 700698
rect 288938 700646 288950 700698
rect 289002 700646 289014 700698
rect 289066 700646 289078 700698
rect 289130 700646 289142 700698
rect 289194 700646 289206 700698
rect 289258 700646 289270 700698
rect 289322 700646 289334 700698
rect 289386 700646 324822 700698
rect 324874 700646 324886 700698
rect 324938 700646 324950 700698
rect 325002 700646 325014 700698
rect 325066 700646 325078 700698
rect 325130 700646 325142 700698
rect 325194 700646 325206 700698
rect 325258 700646 325270 700698
rect 325322 700646 325334 700698
rect 325386 700646 360822 700698
rect 360874 700646 360886 700698
rect 360938 700646 360950 700698
rect 361002 700646 361014 700698
rect 361066 700646 361078 700698
rect 361130 700646 361142 700698
rect 361194 700646 361206 700698
rect 361258 700646 361270 700698
rect 361322 700646 361334 700698
rect 361386 700646 396822 700698
rect 396874 700646 396886 700698
rect 396938 700646 396950 700698
rect 397002 700646 397014 700698
rect 397066 700646 397078 700698
rect 397130 700646 397142 700698
rect 397194 700646 397206 700698
rect 397258 700646 397270 700698
rect 397322 700646 397334 700698
rect 397386 700646 432822 700698
rect 432874 700646 432886 700698
rect 432938 700646 432950 700698
rect 433002 700646 433014 700698
rect 433066 700646 433078 700698
rect 433130 700646 433142 700698
rect 433194 700646 433206 700698
rect 433258 700646 433270 700698
rect 433322 700646 433334 700698
rect 433386 700646 468822 700698
rect 468874 700646 468886 700698
rect 468938 700646 468950 700698
rect 469002 700646 469014 700698
rect 469066 700646 469078 700698
rect 469130 700646 469142 700698
rect 469194 700646 469206 700698
rect 469258 700646 469270 700698
rect 469322 700646 469334 700698
rect 469386 700646 504822 700698
rect 504874 700646 504886 700698
rect 504938 700646 504950 700698
rect 505002 700646 505014 700698
rect 505066 700646 505078 700698
rect 505130 700646 505142 700698
rect 505194 700646 505206 700698
rect 505258 700646 505270 700698
rect 505322 700646 505334 700698
rect 505386 700646 540822 700698
rect 540874 700646 540886 700698
rect 540938 700646 540950 700698
rect 541002 700646 541014 700698
rect 541066 700646 541078 700698
rect 541130 700646 541142 700698
rect 541194 700646 541206 700698
rect 541258 700646 541270 700698
rect 541322 700646 541334 700698
rect 541386 700646 576822 700698
rect 576874 700646 576886 700698
rect 576938 700646 576950 700698
rect 577002 700646 577014 700698
rect 577066 700646 577078 700698
rect 577130 700646 577142 700698
rect 577194 700646 577206 700698
rect 577258 700646 577270 700698
rect 577322 700646 577334 700698
rect 577386 700646 582820 700698
rect 1104 700624 582820 700646
rect 242250 700544 242256 700596
rect 242308 700584 242314 700596
rect 462314 700584 462320 700596
rect 242308 700556 462320 700584
rect 242308 700544 242314 700556
rect 462314 700544 462320 700556
rect 462372 700544 462378 700596
rect 246942 700476 246948 700528
rect 247000 700516 247006 700528
rect 478506 700516 478512 700528
rect 247000 700488 478512 700516
rect 247000 700476 247006 700488
rect 478506 700476 478512 700488
rect 478564 700476 478570 700528
rect 89162 700408 89168 700460
rect 89220 700448 89226 700460
rect 332134 700448 332140 700460
rect 89220 700420 332140 700448
rect 89220 700408 89226 700420
rect 332134 700408 332140 700420
rect 332192 700408 332198 700460
rect 202782 700340 202788 700392
rect 202840 700380 202846 700392
rect 292574 700380 292580 700392
rect 202840 700352 292580 700380
rect 202840 700340 202846 700352
rect 292574 700340 292580 700352
rect 292632 700340 292638 700392
rect 292666 700340 292672 700392
rect 292724 700380 292730 700392
rect 300118 700380 300124 700392
rect 292724 700352 300124 700380
rect 292724 700340 292730 700352
rect 300118 700340 300124 700352
rect 300176 700340 300182 700392
rect 300210 700340 300216 700392
rect 300268 700380 300274 700392
rect 543458 700380 543464 700392
rect 300268 700352 543464 700380
rect 300268 700340 300274 700352
rect 543458 700340 543464 700352
rect 543516 700340 543522 700392
rect 72694 700272 72700 700324
rect 72752 700312 72758 700324
rect 327442 700312 327448 700324
rect 72752 700284 327448 700312
rect 72752 700272 72758 700284
rect 327442 700272 327448 700284
rect 327500 700272 327506 700324
rect 170306 700204 170312 700256
rect 170364 700244 170370 700256
rect 308490 700244 308496 700256
rect 170364 700216 308496 700244
rect 170364 700204 170370 700216
rect 308490 700204 308496 700216
rect 308548 700204 308554 700256
rect 331217 700247 331275 700253
rect 331217 700213 331229 700247
rect 331263 700244 331275 700247
rect 336001 700247 336059 700253
rect 336001 700244 336013 700247
rect 331263 700216 336013 700244
rect 331263 700213 331275 700216
rect 331217 700207 331275 700213
rect 336001 700213 336013 700216
rect 336047 700213 336059 700247
rect 336001 700207 336059 700213
rect 338117 700247 338175 700253
rect 338117 700213 338129 700247
rect 338163 700244 338175 700247
rect 347685 700247 347743 700253
rect 347685 700244 347697 700247
rect 338163 700216 347697 700244
rect 338163 700213 338175 700216
rect 338117 700207 338175 700213
rect 347685 700213 347697 700216
rect 347731 700213 347743 700247
rect 347685 700207 347743 700213
rect 1104 700154 582820 700176
rect 1104 700102 18822 700154
rect 18874 700102 18886 700154
rect 18938 700102 18950 700154
rect 19002 700102 19014 700154
rect 19066 700102 19078 700154
rect 19130 700102 19142 700154
rect 19194 700102 19206 700154
rect 19258 700102 19270 700154
rect 19322 700102 19334 700154
rect 19386 700102 54822 700154
rect 54874 700102 54886 700154
rect 54938 700102 54950 700154
rect 55002 700102 55014 700154
rect 55066 700102 55078 700154
rect 55130 700102 55142 700154
rect 55194 700102 55206 700154
rect 55258 700102 55270 700154
rect 55322 700102 55334 700154
rect 55386 700102 90822 700154
rect 90874 700102 90886 700154
rect 90938 700102 90950 700154
rect 91002 700102 91014 700154
rect 91066 700102 91078 700154
rect 91130 700102 91142 700154
rect 91194 700102 91206 700154
rect 91258 700102 91270 700154
rect 91322 700102 91334 700154
rect 91386 700102 126822 700154
rect 126874 700102 126886 700154
rect 126938 700102 126950 700154
rect 127002 700102 127014 700154
rect 127066 700102 127078 700154
rect 127130 700102 127142 700154
rect 127194 700102 127206 700154
rect 127258 700102 127270 700154
rect 127322 700102 127334 700154
rect 127386 700102 162822 700154
rect 162874 700102 162886 700154
rect 162938 700102 162950 700154
rect 163002 700102 163014 700154
rect 163066 700102 163078 700154
rect 163130 700102 163142 700154
rect 163194 700102 163206 700154
rect 163258 700102 163270 700154
rect 163322 700102 163334 700154
rect 163386 700102 198822 700154
rect 198874 700102 198886 700154
rect 198938 700102 198950 700154
rect 199002 700102 199014 700154
rect 199066 700102 199078 700154
rect 199130 700102 199142 700154
rect 199194 700102 199206 700154
rect 199258 700102 199270 700154
rect 199322 700102 199334 700154
rect 199386 700102 234822 700154
rect 234874 700102 234886 700154
rect 234938 700102 234950 700154
rect 235002 700102 235014 700154
rect 235066 700102 235078 700154
rect 235130 700102 235142 700154
rect 235194 700102 235206 700154
rect 235258 700102 235270 700154
rect 235322 700102 235334 700154
rect 235386 700102 270822 700154
rect 270874 700102 270886 700154
rect 270938 700102 270950 700154
rect 271002 700102 271014 700154
rect 271066 700102 271078 700154
rect 271130 700102 271142 700154
rect 271194 700102 271206 700154
rect 271258 700102 271270 700154
rect 271322 700102 271334 700154
rect 271386 700102 306822 700154
rect 306874 700102 306886 700154
rect 306938 700102 306950 700154
rect 307002 700102 307014 700154
rect 307066 700102 307078 700154
rect 307130 700102 307142 700154
rect 307194 700102 307206 700154
rect 307258 700102 307270 700154
rect 307322 700102 307334 700154
rect 307386 700102 342822 700154
rect 342874 700102 342886 700154
rect 342938 700102 342950 700154
rect 343002 700102 343014 700154
rect 343066 700102 343078 700154
rect 343130 700102 343142 700154
rect 343194 700102 343206 700154
rect 343258 700102 343270 700154
rect 343322 700102 343334 700154
rect 343386 700102 378822 700154
rect 378874 700102 378886 700154
rect 378938 700102 378950 700154
rect 379002 700102 379014 700154
rect 379066 700102 379078 700154
rect 379130 700102 379142 700154
rect 379194 700102 379206 700154
rect 379258 700102 379270 700154
rect 379322 700102 379334 700154
rect 379386 700102 414822 700154
rect 414874 700102 414886 700154
rect 414938 700102 414950 700154
rect 415002 700102 415014 700154
rect 415066 700102 415078 700154
rect 415130 700102 415142 700154
rect 415194 700102 415206 700154
rect 415258 700102 415270 700154
rect 415322 700102 415334 700154
rect 415386 700102 450822 700154
rect 450874 700102 450886 700154
rect 450938 700102 450950 700154
rect 451002 700102 451014 700154
rect 451066 700102 451078 700154
rect 451130 700102 451142 700154
rect 451194 700102 451206 700154
rect 451258 700102 451270 700154
rect 451322 700102 451334 700154
rect 451386 700102 486822 700154
rect 486874 700102 486886 700154
rect 486938 700102 486950 700154
rect 487002 700102 487014 700154
rect 487066 700102 487078 700154
rect 487130 700102 487142 700154
rect 487194 700102 487206 700154
rect 487258 700102 487270 700154
rect 487322 700102 487334 700154
rect 487386 700102 522822 700154
rect 522874 700102 522886 700154
rect 522938 700102 522950 700154
rect 523002 700102 523014 700154
rect 523066 700102 523078 700154
rect 523130 700102 523142 700154
rect 523194 700102 523206 700154
rect 523258 700102 523270 700154
rect 523322 700102 523334 700154
rect 523386 700102 558822 700154
rect 558874 700102 558886 700154
rect 558938 700102 558950 700154
rect 559002 700102 559014 700154
rect 559066 700102 559078 700154
rect 559130 700102 559142 700154
rect 559194 700102 559206 700154
rect 559258 700102 559270 700154
rect 559322 700102 559334 700154
rect 559386 700102 582820 700154
rect 1104 700080 582820 700102
rect 267642 700000 267648 700052
rect 267700 700040 267706 700052
rect 283742 700040 283748 700052
rect 267700 700012 283748 700040
rect 267700 700000 267706 700012
rect 283742 700000 283748 700012
rect 283800 700000 283806 700052
rect 283834 700000 283840 700052
rect 283892 700040 283898 700052
rect 289446 700040 289452 700052
rect 283892 700012 289452 700040
rect 283892 700000 283898 700012
rect 289446 700000 289452 700012
rect 289504 700000 289510 700052
rect 289538 700000 289544 700052
rect 289596 700040 289602 700052
rect 292393 700043 292451 700049
rect 292393 700040 292405 700043
rect 289596 700012 292405 700040
rect 289596 700000 289602 700012
rect 292393 700009 292405 700012
rect 292439 700009 292451 700043
rect 292393 700003 292451 700009
rect 292485 700043 292543 700049
rect 292485 700009 292497 700043
rect 292531 700040 292543 700043
rect 413646 700040 413652 700052
rect 292531 700012 413652 700040
rect 292531 700009 292543 700012
rect 292485 700003 292543 700009
rect 413646 700000 413652 700012
rect 413704 700000 413710 700052
rect 233237 699975 233295 699981
rect 233237 699941 233249 699975
rect 233283 699972 233295 699975
rect 244182 699972 244188 699984
rect 233283 699944 244188 699972
rect 233283 699941 233295 699944
rect 233237 699935 233295 699941
rect 244182 699932 244188 699944
rect 244240 699932 244246 699984
rect 251082 699932 251088 699984
rect 251140 699972 251146 699984
rect 253842 699972 253848 699984
rect 251140 699944 253848 699972
rect 251140 699932 251146 699944
rect 253842 699932 253848 699944
rect 253900 699932 253906 699984
rect 265894 699932 265900 699984
rect 265952 699972 265958 699984
rect 364978 699972 364984 699984
rect 265952 699944 364984 699972
rect 265952 699932 265958 699944
rect 364978 699932 364984 699944
rect 365036 699932 365042 699984
rect 218974 699864 218980 699916
rect 219032 699904 219038 699916
rect 302050 699904 302056 699916
rect 219032 699876 302056 699904
rect 219032 699864 219038 699876
rect 302050 699864 302056 699876
rect 302108 699864 302114 699916
rect 302145 699907 302203 699913
rect 302145 699873 302157 699907
rect 302191 699904 302203 699907
rect 306745 699907 306803 699913
rect 306745 699904 306757 699907
rect 302191 699876 306757 699904
rect 302191 699873 302203 699876
rect 302145 699867 302203 699873
rect 306745 699873 306757 699876
rect 306791 699873 306803 699907
rect 306745 699867 306803 699873
rect 306837 699907 306895 699913
rect 306837 699873 306849 699907
rect 306883 699904 306895 699907
rect 318797 699907 318855 699913
rect 306883 699876 316724 699904
rect 306883 699873 306895 699876
rect 306837 699867 306895 699873
rect 270494 699836 270500 699848
rect 241440 699808 241560 699836
rect 241440 699777 241468 699808
rect 241532 699780 241560 699808
rect 253952 699808 270500 699836
rect 200117 699771 200175 699777
rect 200117 699737 200129 699771
rect 200163 699768 200175 699771
rect 209685 699771 209743 699777
rect 209685 699768 209697 699771
rect 200163 699740 209697 699768
rect 200163 699737 200175 699740
rect 200117 699731 200175 699737
rect 209685 699737 209697 699740
rect 209731 699737 209743 699771
rect 209685 699731 209743 699737
rect 219437 699771 219495 699777
rect 219437 699737 219449 699771
rect 219483 699768 219495 699771
rect 229005 699771 229063 699777
rect 229005 699768 229017 699771
rect 219483 699740 229017 699768
rect 219483 699737 219495 699740
rect 219437 699731 219495 699737
rect 229005 699737 229017 699740
rect 229051 699737 229063 699771
rect 229005 699731 229063 699737
rect 241425 699771 241483 699777
rect 241425 699737 241437 699771
rect 241471 699737 241483 699771
rect 241425 699731 241483 699737
rect 241514 699728 241520 699780
rect 241572 699728 241578 699780
rect 251082 699728 251088 699780
rect 251140 699768 251146 699780
rect 253952 699768 253980 699808
rect 270494 699796 270500 699808
rect 270552 699796 270558 699848
rect 270586 699796 270592 699848
rect 270644 699836 270650 699848
rect 277949 699839 278007 699845
rect 277949 699836 277961 699839
rect 270644 699808 277961 699836
rect 270644 699796 270650 699808
rect 277949 699805 277961 699808
rect 277995 699805 278007 699839
rect 292482 699836 292488 699848
rect 277949 699799 278007 699805
rect 278056 699808 292488 699836
rect 251140 699740 253980 699768
rect 251140 699728 251146 699740
rect 263870 699728 263876 699780
rect 263928 699768 263934 699780
rect 273530 699768 273536 699780
rect 263928 699740 273536 699768
rect 263928 699728 263934 699740
rect 273530 699728 273536 699740
rect 273588 699728 273594 699780
rect 275738 699728 275744 699780
rect 275796 699768 275802 699780
rect 278056 699768 278084 699808
rect 292482 699796 292488 699808
rect 292540 699796 292546 699848
rect 301958 699796 301964 699848
rect 302016 699836 302022 699848
rect 302016 699808 311940 699836
rect 302016 699796 302022 699808
rect 275796 699740 278084 699768
rect 278133 699771 278191 699777
rect 275796 699728 275802 699740
rect 278133 699737 278145 699771
rect 278179 699768 278191 699771
rect 292298 699768 292304 699780
rect 278179 699740 292304 699768
rect 278179 699737 278191 699740
rect 278133 699731 278191 699737
rect 292298 699728 292304 699740
rect 292356 699728 292362 699780
rect 292666 699728 292672 699780
rect 292724 699768 292730 699780
rect 306377 699771 306435 699777
rect 306377 699768 306389 699771
rect 292724 699740 306389 699768
rect 292724 699728 292730 699740
rect 306377 699737 306389 699740
rect 306423 699737 306435 699771
rect 311912 699768 311940 699808
rect 316696 699768 316724 699876
rect 318797 699873 318809 699907
rect 318843 699904 318855 699907
rect 325421 699907 325479 699913
rect 318843 699876 321600 699904
rect 318843 699873 318855 699876
rect 318797 699867 318855 699873
rect 321572 699836 321600 699876
rect 325421 699873 325433 699907
rect 325467 699904 325479 699907
rect 340782 699904 340788 699916
rect 325467 699876 340788 699904
rect 325467 699873 325479 699876
rect 325421 699867 325479 699873
rect 340782 699864 340788 699876
rect 340840 699864 340846 699916
rect 331217 699839 331275 699845
rect 331217 699836 331229 699839
rect 321572 699808 331229 699836
rect 331217 699805 331229 699808
rect 331263 699805 331275 699839
rect 331217 699799 331275 699805
rect 347685 699839 347743 699845
rect 347685 699805 347697 699839
rect 347731 699836 347743 699839
rect 348786 699836 348792 699848
rect 347731 699808 348792 699836
rect 347731 699805 347743 699808
rect 347685 699799 347743 699805
rect 348786 699796 348792 699808
rect 348844 699796 348850 699848
rect 321465 699771 321523 699777
rect 321465 699768 321477 699771
rect 311912 699740 312032 699768
rect 316696 699740 321477 699768
rect 306377 699731 306435 699737
rect 179322 699660 179328 699712
rect 179380 699700 179386 699712
rect 180981 699703 181039 699709
rect 180981 699700 180993 699703
rect 179380 699672 180993 699700
rect 179380 699660 179386 699672
rect 180981 699669 180993 699672
rect 181027 699669 181039 699703
rect 180981 699663 181039 699669
rect 190181 699703 190239 699709
rect 190181 699669 190193 699703
rect 190227 699700 190239 699703
rect 190733 699703 190791 699709
rect 190733 699700 190745 699703
rect 190227 699672 190745 699700
rect 190227 699669 190239 699672
rect 190181 699663 190239 699669
rect 190733 699669 190745 699672
rect 190779 699669 190791 699703
rect 190733 699663 190791 699669
rect 199841 699703 199899 699709
rect 199841 699669 199853 699703
rect 199887 699700 199899 699703
rect 200301 699703 200359 699709
rect 200301 699700 200313 699703
rect 199887 699672 200313 699700
rect 199887 699669 199899 699672
rect 199841 699663 199899 699669
rect 200301 699669 200313 699672
rect 200347 699669 200359 699703
rect 200301 699663 200359 699669
rect 209501 699703 209559 699709
rect 209501 699669 209513 699703
rect 209547 699700 209559 699703
rect 210053 699703 210111 699709
rect 210053 699700 210065 699703
rect 209547 699672 210065 699700
rect 209547 699669 209559 699672
rect 209501 699663 209559 699669
rect 210053 699669 210065 699672
rect 210099 699669 210111 699703
rect 210053 699663 210111 699669
rect 219161 699703 219219 699709
rect 219161 699669 219173 699703
rect 219207 699700 219219 699703
rect 219621 699703 219679 699709
rect 219621 699700 219633 699703
rect 219207 699672 219633 699700
rect 219207 699669 219219 699672
rect 219161 699663 219219 699669
rect 219621 699669 219633 699672
rect 219667 699669 219679 699703
rect 219621 699663 219679 699669
rect 228821 699703 228879 699709
rect 228821 699669 228833 699703
rect 228867 699700 228879 699703
rect 229373 699703 229431 699709
rect 229373 699700 229385 699703
rect 228867 699672 229385 699700
rect 228867 699669 228879 699672
rect 228821 699663 228879 699669
rect 229373 699669 229385 699672
rect 229419 699669 229431 699703
rect 229373 699663 229431 699669
rect 273162 699660 273168 699712
rect 273220 699700 273226 699712
rect 282914 699700 282920 699712
rect 273220 699672 282920 699700
rect 273220 699660 273226 699672
rect 282914 699660 282920 699672
rect 282972 699660 282978 699712
rect 288434 699660 288440 699712
rect 288492 699700 288498 699712
rect 292209 699703 292267 699709
rect 292209 699700 292221 699703
rect 288492 699672 292221 699700
rect 288492 699660 288498 699672
rect 292209 699669 292221 699672
rect 292255 699669 292267 699703
rect 292209 699663 292267 699669
rect 292485 699703 292543 699709
rect 292485 699669 292497 699703
rect 292531 699700 292543 699703
rect 292574 699700 292580 699712
rect 292531 699672 292580 699700
rect 292531 699669 292543 699672
rect 292485 699663 292543 699669
rect 292574 699660 292580 699672
rect 292632 699660 292638 699712
rect 292761 699703 292819 699709
rect 292761 699669 292773 699703
rect 292807 699700 292819 699703
rect 301961 699703 302019 699709
rect 301961 699700 301973 699703
rect 292807 699672 301973 699700
rect 292807 699669 292819 699672
rect 292761 699663 292819 699669
rect 301961 699669 301973 699672
rect 302007 699669 302019 699703
rect 301961 699663 302019 699669
rect 302053 699703 302111 699709
rect 302053 699669 302065 699703
rect 302099 699700 302111 699703
rect 306469 699703 306527 699709
rect 306469 699700 306481 699703
rect 302099 699672 306481 699700
rect 302099 699669 302111 699672
rect 302053 699663 302111 699669
rect 306469 699669 306481 699672
rect 306515 699669 306527 699703
rect 306469 699663 306527 699669
rect 306653 699703 306711 699709
rect 306653 699669 306665 699703
rect 306699 699700 306711 699703
rect 311894 699700 311900 699712
rect 306699 699672 311900 699700
rect 306699 699669 306711 699672
rect 306653 699663 306711 699669
rect 311894 699660 311900 699672
rect 311952 699660 311958 699712
rect 312004 699700 312032 699740
rect 321465 699737 321477 699740
rect 321511 699737 321523 699771
rect 321465 699731 321523 699737
rect 321557 699771 321615 699777
rect 321557 699737 321569 699771
rect 321603 699768 321615 699771
rect 332502 699768 332508 699780
rect 321603 699740 332508 699768
rect 321603 699737 321615 699740
rect 321557 699731 321615 699737
rect 332502 699728 332508 699740
rect 332560 699728 332566 699780
rect 336001 699771 336059 699777
rect 336001 699737 336013 699771
rect 336047 699768 336059 699771
rect 338117 699771 338175 699777
rect 338117 699768 338129 699771
rect 336047 699740 338129 699768
rect 336047 699737 336059 699740
rect 336001 699731 336059 699737
rect 338117 699737 338129 699740
rect 338163 699737 338175 699771
rect 338117 699731 338175 699737
rect 354401 699771 354459 699777
rect 354401 699737 354413 699771
rect 354447 699768 354459 699771
rect 364245 699771 364303 699777
rect 364245 699768 364257 699771
rect 354447 699740 364257 699768
rect 354447 699737 354459 699740
rect 354401 699731 354459 699737
rect 364245 699737 364257 699740
rect 364291 699737 364303 699771
rect 364245 699731 364303 699737
rect 318797 699703 318855 699709
rect 318797 699700 318809 699703
rect 312004 699672 318809 699700
rect 318797 699669 318809 699672
rect 318843 699669 318855 699703
rect 318797 699663 318855 699669
rect 325329 699703 325387 699709
rect 325329 699669 325341 699703
rect 325375 699700 325387 699703
rect 325973 699703 326031 699709
rect 325973 699700 325985 699703
rect 325375 699672 325985 699700
rect 325375 699669 325387 699672
rect 325329 699663 325387 699669
rect 325973 699669 325985 699672
rect 326019 699669 326031 699703
rect 325973 699663 326031 699669
rect 331214 699660 331220 699712
rect 331272 699700 331278 699712
rect 343542 699700 343548 699712
rect 331272 699672 343548 699700
rect 331272 699660 331278 699672
rect 343542 699660 343548 699672
rect 343600 699660 343606 699712
rect 354309 699703 354367 699709
rect 354309 699669 354321 699703
rect 354355 699700 354367 699703
rect 354769 699703 354827 699709
rect 354769 699700 354781 699703
rect 354355 699672 354781 699700
rect 354355 699669 354367 699672
rect 354309 699663 354367 699669
rect 354769 699669 354781 699672
rect 354815 699669 354827 699703
rect 354769 699663 354827 699669
rect 364153 699703 364211 699709
rect 364153 699669 364165 699703
rect 364199 699700 364211 699703
rect 373721 699703 373779 699709
rect 373721 699700 373733 699703
rect 364199 699672 373733 699700
rect 364199 699669 364211 699672
rect 364153 699663 364211 699669
rect 373721 699669 373733 699672
rect 373767 699669 373779 699703
rect 373721 699663 373779 699669
rect 373813 699703 373871 699709
rect 373813 699669 373825 699703
rect 373859 699700 373871 699703
rect 373994 699700 374000 699712
rect 373859 699672 374000 699700
rect 373859 699669 373871 699672
rect 373813 699663 373871 699669
rect 373994 699660 374000 699672
rect 374052 699660 374058 699712
rect 1104 699610 582820 699632
rect 1104 699558 36822 699610
rect 36874 699558 36886 699610
rect 36938 699558 36950 699610
rect 37002 699558 37014 699610
rect 37066 699558 37078 699610
rect 37130 699558 37142 699610
rect 37194 699558 37206 699610
rect 37258 699558 37270 699610
rect 37322 699558 37334 699610
rect 37386 699558 72822 699610
rect 72874 699558 72886 699610
rect 72938 699558 72950 699610
rect 73002 699558 73014 699610
rect 73066 699558 73078 699610
rect 73130 699558 73142 699610
rect 73194 699558 73206 699610
rect 73258 699558 73270 699610
rect 73322 699558 73334 699610
rect 73386 699558 108822 699610
rect 108874 699558 108886 699610
rect 108938 699558 108950 699610
rect 109002 699558 109014 699610
rect 109066 699558 109078 699610
rect 109130 699558 109142 699610
rect 109194 699558 109206 699610
rect 109258 699558 109270 699610
rect 109322 699558 109334 699610
rect 109386 699558 144822 699610
rect 144874 699558 144886 699610
rect 144938 699558 144950 699610
rect 145002 699558 145014 699610
rect 145066 699558 145078 699610
rect 145130 699558 145142 699610
rect 145194 699558 145206 699610
rect 145258 699558 145270 699610
rect 145322 699558 145334 699610
rect 145386 699558 180822 699610
rect 180874 699558 180886 699610
rect 180938 699558 180950 699610
rect 181002 699558 181014 699610
rect 181066 699558 181078 699610
rect 181130 699558 181142 699610
rect 181194 699558 181206 699610
rect 181258 699558 181270 699610
rect 181322 699558 181334 699610
rect 181386 699558 216822 699610
rect 216874 699558 216886 699610
rect 216938 699558 216950 699610
rect 217002 699558 217014 699610
rect 217066 699558 217078 699610
rect 217130 699558 217142 699610
rect 217194 699558 217206 699610
rect 217258 699558 217270 699610
rect 217322 699558 217334 699610
rect 217386 699558 252822 699610
rect 252874 699558 252886 699610
rect 252938 699558 252950 699610
rect 253002 699558 253014 699610
rect 253066 699558 253078 699610
rect 253130 699558 253142 699610
rect 253194 699558 253206 699610
rect 253258 699558 253270 699610
rect 253322 699558 253334 699610
rect 253386 699558 288822 699610
rect 288874 699558 288886 699610
rect 288938 699558 288950 699610
rect 289002 699558 289014 699610
rect 289066 699558 289078 699610
rect 289130 699558 289142 699610
rect 289194 699558 289206 699610
rect 289258 699558 289270 699610
rect 289322 699558 289334 699610
rect 289386 699558 324822 699610
rect 324874 699558 324886 699610
rect 324938 699558 324950 699610
rect 325002 699558 325014 699610
rect 325066 699558 325078 699610
rect 325130 699558 325142 699610
rect 325194 699558 325206 699610
rect 325258 699558 325270 699610
rect 325322 699558 325334 699610
rect 325386 699558 360822 699610
rect 360874 699558 360886 699610
rect 360938 699558 360950 699610
rect 361002 699558 361014 699610
rect 361066 699558 361078 699610
rect 361130 699558 361142 699610
rect 361194 699558 361206 699610
rect 361258 699558 361270 699610
rect 361322 699558 361334 699610
rect 361386 699558 396822 699610
rect 396874 699558 396886 699610
rect 396938 699558 396950 699610
rect 397002 699558 397014 699610
rect 397066 699558 397078 699610
rect 397130 699558 397142 699610
rect 397194 699558 397206 699610
rect 397258 699558 397270 699610
rect 397322 699558 397334 699610
rect 397386 699558 432822 699610
rect 432874 699558 432886 699610
rect 432938 699558 432950 699610
rect 433002 699558 433014 699610
rect 433066 699558 433078 699610
rect 433130 699558 433142 699610
rect 433194 699558 433206 699610
rect 433258 699558 433270 699610
rect 433322 699558 433334 699610
rect 433386 699558 468822 699610
rect 468874 699558 468886 699610
rect 468938 699558 468950 699610
rect 469002 699558 469014 699610
rect 469066 699558 469078 699610
rect 469130 699558 469142 699610
rect 469194 699558 469206 699610
rect 469258 699558 469270 699610
rect 469322 699558 469334 699610
rect 469386 699558 504822 699610
rect 504874 699558 504886 699610
rect 504938 699558 504950 699610
rect 505002 699558 505014 699610
rect 505066 699558 505078 699610
rect 505130 699558 505142 699610
rect 505194 699558 505206 699610
rect 505258 699558 505270 699610
rect 505322 699558 505334 699610
rect 505386 699558 540822 699610
rect 540874 699558 540886 699610
rect 540938 699558 540950 699610
rect 541002 699558 541014 699610
rect 541066 699558 541078 699610
rect 541130 699558 541142 699610
rect 541194 699558 541206 699610
rect 541258 699558 541270 699610
rect 541322 699558 541334 699610
rect 541386 699558 576822 699610
rect 576874 699558 576886 699610
rect 576938 699558 576950 699610
rect 577002 699558 577014 699610
rect 577066 699558 577078 699610
rect 577130 699558 577142 699610
rect 577194 699558 577206 699610
rect 577258 699558 577270 699610
rect 577322 699558 577334 699610
rect 577386 699558 582820 699610
rect 1104 699536 582820 699558
rect 86034 699456 86040 699508
rect 86092 699496 86098 699508
rect 373813 699499 373871 699505
rect 373813 699496 373825 699499
rect 86092 699468 373825 699496
rect 86092 699456 86098 699468
rect 373813 699465 373825 699468
rect 373859 699465 373871 699499
rect 373813 699459 373871 699465
rect 373905 699499 373963 699505
rect 373905 699465 373917 699499
rect 373951 699496 373963 699499
rect 403158 699496 403164 699508
rect 373951 699468 403164 699496
rect 373951 699465 373963 699468
rect 373905 699459 373963 699465
rect 403158 699456 403164 699468
rect 403216 699456 403222 699508
rect 404262 699456 404268 699508
rect 404320 699496 404326 699508
rect 417326 699496 417332 699508
rect 404320 699468 417332 699496
rect 404320 699456 404326 699468
rect 417326 699456 417332 699468
rect 417384 699456 417390 699508
rect 71774 699388 71780 699440
rect 71832 699428 71838 699440
rect 273254 699428 273260 699440
rect 71832 699400 273260 699428
rect 71832 699388 71838 699400
rect 273254 699388 273260 699400
rect 273312 699388 273318 699440
rect 273346 699388 273352 699440
rect 273404 699428 273410 699440
rect 282914 699428 282920 699440
rect 273404 699400 282920 699428
rect 273404 699388 273410 699400
rect 282914 699388 282920 699400
rect 282972 699388 282978 699440
rect 283006 699388 283012 699440
rect 283064 699428 283070 699440
rect 292577 699431 292635 699437
rect 292577 699428 292589 699431
rect 283064 699400 292589 699428
rect 283064 699388 283070 699400
rect 292577 699397 292589 699400
rect 292623 699397 292635 699431
rect 292577 699391 292635 699397
rect 292666 699388 292672 699440
rect 292724 699428 292730 699440
rect 302053 699431 302111 699437
rect 302053 699428 302065 699431
rect 292724 699400 302065 699428
rect 292724 699388 292730 699400
rect 302053 699397 302065 699400
rect 302099 699397 302111 699431
rect 302053 699391 302111 699397
rect 302142 699388 302148 699440
rect 302200 699428 302206 699440
rect 354677 699431 354735 699437
rect 354677 699428 354689 699431
rect 302200 699400 354689 699428
rect 302200 699388 302206 699400
rect 354677 699397 354689 699400
rect 354723 699397 354735 699431
rect 354677 699391 354735 699397
rect 354769 699431 354827 699437
rect 354769 699397 354781 699431
rect 354815 699428 354827 699431
rect 364153 699431 364211 699437
rect 364153 699428 364165 699431
rect 354815 699400 364165 699428
rect 354815 699397 354827 699400
rect 354769 699391 354827 699397
rect 364153 699397 364165 699400
rect 364199 699397 364211 699431
rect 364153 699391 364211 699397
rect 364245 699431 364303 699437
rect 364245 699397 364257 699431
rect 364291 699428 364303 699431
rect 431586 699428 431592 699440
rect 364291 699400 431592 699428
rect 364291 699397 364303 699400
rect 364245 699391 364303 699397
rect 431586 699388 431592 699400
rect 431644 699388 431650 699440
rect 114370 699320 114376 699372
rect 114428 699360 114434 699372
rect 407942 699360 407948 699372
rect 114428 699332 407948 699360
rect 114428 699320 114434 699332
rect 407942 699320 407948 699332
rect 408000 699320 408006 699372
rect 161750 699252 161756 699304
rect 161808 699292 161814 699304
rect 577866 699292 577872 699304
rect 161808 699264 577872 699292
rect 161808 699252 161814 699264
rect 577866 699252 577872 699264
rect 577924 699252 577930 699304
rect 5166 699184 5172 699236
rect 5224 699224 5230 699236
rect 180981 699227 181039 699233
rect 5224 699196 180932 699224
rect 5224 699184 5230 699196
rect 133322 699116 133328 699168
rect 133380 699156 133386 699168
rect 180794 699156 180800 699168
rect 133380 699128 180800 699156
rect 133380 699116 133386 699128
rect 180794 699116 180800 699128
rect 180852 699116 180858 699168
rect 180904 699156 180932 699196
rect 180981 699193 180993 699227
rect 181027 699224 181039 699227
rect 190181 699227 190239 699233
rect 190181 699224 190193 699227
rect 181027 699196 190193 699224
rect 181027 699193 181039 699196
rect 180981 699187 181039 699193
rect 190181 699193 190193 699196
rect 190227 699193 190239 699227
rect 190733 699227 190791 699233
rect 190181 699187 190239 699193
rect 190288 699196 190592 699224
rect 190288 699156 190316 699196
rect 180904 699128 190316 699156
rect 190362 699116 190368 699168
rect 190420 699156 190426 699168
rect 190454 699156 190460 699168
rect 190420 699128 190460 699156
rect 190420 699116 190426 699128
rect 190454 699116 190460 699128
rect 190512 699116 190518 699168
rect 190564 699156 190592 699196
rect 190733 699193 190745 699227
rect 190779 699224 190791 699227
rect 199841 699227 199899 699233
rect 199841 699224 199853 699227
rect 190779 699196 199853 699224
rect 190779 699193 190791 699196
rect 190733 699187 190791 699193
rect 199841 699193 199853 699196
rect 199887 699193 199899 699227
rect 200301 699227 200359 699233
rect 199841 699187 199899 699193
rect 199948 699196 200252 699224
rect 199948 699156 199976 699196
rect 190564 699128 199976 699156
rect 200022 699116 200028 699168
rect 200080 699156 200086 699168
rect 200117 699159 200175 699165
rect 200117 699156 200129 699159
rect 200080 699128 200129 699156
rect 200080 699116 200086 699128
rect 200117 699125 200129 699128
rect 200163 699125 200175 699159
rect 200224 699156 200252 699196
rect 200301 699193 200313 699227
rect 200347 699224 200359 699227
rect 209501 699227 209559 699233
rect 209501 699224 209513 699227
rect 200347 699196 209513 699224
rect 200347 699193 200359 699196
rect 200301 699187 200359 699193
rect 209501 699193 209513 699196
rect 209547 699193 209559 699227
rect 210053 699227 210111 699233
rect 209501 699187 209559 699193
rect 209608 699196 209912 699224
rect 209608 699156 209636 699196
rect 200224 699128 209636 699156
rect 209685 699159 209743 699165
rect 200117 699119 200175 699125
rect 209685 699125 209697 699159
rect 209731 699156 209743 699159
rect 209774 699156 209780 699168
rect 209731 699128 209780 699156
rect 209731 699125 209743 699128
rect 209685 699119 209743 699125
rect 209774 699116 209780 699128
rect 209832 699116 209838 699168
rect 209884 699156 209912 699196
rect 210053 699193 210065 699227
rect 210099 699224 210111 699227
rect 219161 699227 219219 699233
rect 219161 699224 219173 699227
rect 210099 699196 219173 699224
rect 210099 699193 210111 699196
rect 210053 699187 210111 699193
rect 219161 699193 219173 699196
rect 219207 699193 219219 699227
rect 219621 699227 219679 699233
rect 219161 699187 219219 699193
rect 219268 699196 219572 699224
rect 219268 699156 219296 699196
rect 209884 699128 219296 699156
rect 219342 699116 219348 699168
rect 219400 699156 219406 699168
rect 219437 699159 219495 699165
rect 219437 699156 219449 699159
rect 219400 699128 219449 699156
rect 219400 699116 219406 699128
rect 219437 699125 219449 699128
rect 219483 699125 219495 699159
rect 219544 699156 219572 699196
rect 219621 699193 219633 699227
rect 219667 699224 219679 699227
rect 228821 699227 228879 699233
rect 228821 699224 228833 699227
rect 219667 699196 228833 699224
rect 219667 699193 219679 699196
rect 219621 699187 219679 699193
rect 228821 699193 228833 699196
rect 228867 699193 228879 699227
rect 229373 699227 229431 699233
rect 228821 699187 228879 699193
rect 228928 699196 229232 699224
rect 228928 699156 228956 699196
rect 219544 699128 228956 699156
rect 229005 699159 229063 699165
rect 219437 699119 219495 699125
rect 229005 699125 229017 699159
rect 229051 699156 229063 699159
rect 229094 699156 229100 699168
rect 229051 699128 229100 699156
rect 229051 699125 229063 699128
rect 229005 699119 229063 699125
rect 229094 699116 229100 699128
rect 229152 699116 229158 699168
rect 229204 699156 229232 699196
rect 229373 699193 229385 699227
rect 229419 699224 229431 699227
rect 233237 699227 233295 699233
rect 233237 699224 233249 699227
rect 229419 699196 233249 699224
rect 229419 699193 229431 699196
rect 229373 699187 229431 699193
rect 233237 699193 233249 699196
rect 233283 699193 233295 699227
rect 233237 699187 233295 699193
rect 234706 699184 234712 699236
rect 234764 699224 234770 699236
rect 239493 699227 239551 699233
rect 234764 699196 239444 699224
rect 234764 699184 234770 699196
rect 239309 699159 239367 699165
rect 239309 699156 239321 699159
rect 229204 699128 239321 699156
rect 239309 699125 239321 699128
rect 239355 699125 239367 699159
rect 239416 699156 239444 699196
rect 239493 699193 239505 699227
rect 239539 699224 239551 699227
rect 239539 699196 253796 699224
rect 239539 699193 239551 699196
rect 239493 699187 239551 699193
rect 244090 699156 244096 699168
rect 239416 699128 244096 699156
rect 239309 699119 239367 699125
rect 244090 699116 244096 699128
rect 244148 699116 244154 699168
rect 244182 699116 244188 699168
rect 244240 699156 244246 699168
rect 253658 699156 253664 699168
rect 244240 699128 253664 699156
rect 244240 699116 244246 699128
rect 253658 699116 253664 699128
rect 253716 699116 253722 699168
rect 253768 699156 253796 699196
rect 253842 699184 253848 699236
rect 253900 699224 253906 699236
rect 264977 699227 265035 699233
rect 264977 699224 264989 699227
rect 253900 699196 264989 699224
rect 253900 699184 253906 699196
rect 264977 699193 264989 699196
rect 265023 699193 265035 699227
rect 306377 699227 306435 699233
rect 306377 699224 306389 699227
rect 264977 699187 265035 699193
rect 265084 699196 306389 699224
rect 265084 699156 265112 699196
rect 306377 699193 306389 699196
rect 306423 699193 306435 699227
rect 306377 699187 306435 699193
rect 306469 699227 306527 699233
rect 306469 699193 306481 699227
rect 306515 699224 306527 699227
rect 325329 699227 325387 699233
rect 325329 699224 325341 699227
rect 306515 699196 325341 699224
rect 306515 699193 306527 699196
rect 306469 699187 306527 699193
rect 325329 699193 325341 699196
rect 325375 699193 325387 699227
rect 325329 699187 325387 699193
rect 325605 699227 325663 699233
rect 325605 699193 325617 699227
rect 325651 699224 325663 699227
rect 325973 699227 326031 699233
rect 325651 699196 325832 699224
rect 325651 699193 325663 699196
rect 325605 699187 325663 699193
rect 253768 699128 265112 699156
rect 265161 699159 265219 699165
rect 265161 699125 265173 699159
rect 265207 699156 265219 699159
rect 282730 699156 282736 699168
rect 265207 699128 282736 699156
rect 265207 699125 265219 699128
rect 265161 699119 265219 699125
rect 282730 699116 282736 699128
rect 282788 699116 282794 699168
rect 282822 699116 282828 699168
rect 282880 699156 282886 699168
rect 282914 699156 282920 699168
rect 282880 699128 282920 699156
rect 282880 699116 282886 699128
rect 282914 699116 282920 699128
rect 282972 699116 282978 699168
rect 283006 699116 283012 699168
rect 283064 699156 283070 699168
rect 292390 699156 292396 699168
rect 283064 699128 292396 699156
rect 283064 699116 283070 699128
rect 292390 699116 292396 699128
rect 292448 699116 292454 699168
rect 292482 699116 292488 699168
rect 292540 699156 292546 699168
rect 306653 699159 306711 699165
rect 306653 699156 306665 699159
rect 292540 699128 306665 699156
rect 292540 699116 292546 699128
rect 306653 699125 306665 699128
rect 306699 699125 306711 699159
rect 306653 699119 306711 699125
rect 306745 699159 306803 699165
rect 306745 699125 306757 699159
rect 306791 699156 306803 699159
rect 325421 699159 325479 699165
rect 325421 699156 325433 699159
rect 306791 699128 325433 699156
rect 306791 699125 306803 699128
rect 306745 699119 306803 699125
rect 325421 699125 325433 699128
rect 325467 699125 325479 699159
rect 325421 699119 325479 699125
rect 325510 699116 325516 699168
rect 325568 699156 325574 699168
rect 325694 699156 325700 699168
rect 325568 699128 325700 699156
rect 325568 699116 325574 699128
rect 325694 699116 325700 699128
rect 325752 699116 325758 699168
rect 325804 699156 325832 699196
rect 325973 699193 325985 699227
rect 326019 699224 326031 699227
rect 354309 699227 354367 699233
rect 354309 699224 354321 699227
rect 326019 699196 354321 699224
rect 326019 699193 326031 699196
rect 325973 699187 326031 699193
rect 354309 699193 354321 699196
rect 354355 699193 354367 699227
rect 354309 699187 354367 699193
rect 354585 699227 354643 699233
rect 354585 699193 354597 699227
rect 354631 699224 354643 699227
rect 445754 699224 445760 699236
rect 354631 699196 445760 699224
rect 354631 699193 354643 699196
rect 354585 699187 354643 699193
rect 445754 699184 445760 699196
rect 445812 699184 445818 699236
rect 340693 699159 340751 699165
rect 340693 699156 340705 699159
rect 325804 699128 340705 699156
rect 340693 699125 340705 699128
rect 340739 699125 340751 699159
rect 340693 699119 340751 699125
rect 340782 699116 340788 699168
rect 340840 699156 340846 699168
rect 354401 699159 354459 699165
rect 354401 699156 354413 699159
rect 340840 699128 354413 699156
rect 340840 699116 340846 699128
rect 354401 699125 354413 699128
rect 354447 699125 354459 699159
rect 354401 699119 354459 699125
rect 354490 699116 354496 699168
rect 354548 699156 354554 699168
rect 579154 699156 579160 699168
rect 354548 699128 579160 699156
rect 354548 699116 354554 699128
rect 579154 699116 579160 699128
rect 579212 699116 579218 699168
rect 1104 699066 582820 699088
rect 1104 699014 18822 699066
rect 18874 699014 18886 699066
rect 18938 699014 18950 699066
rect 19002 699014 19014 699066
rect 19066 699014 19078 699066
rect 19130 699014 19142 699066
rect 19194 699014 19206 699066
rect 19258 699014 19270 699066
rect 19322 699014 19334 699066
rect 19386 699014 54822 699066
rect 54874 699014 54886 699066
rect 54938 699014 54950 699066
rect 55002 699014 55014 699066
rect 55066 699014 55078 699066
rect 55130 699014 55142 699066
rect 55194 699014 55206 699066
rect 55258 699014 55270 699066
rect 55322 699014 55334 699066
rect 55386 699014 90822 699066
rect 90874 699014 90886 699066
rect 90938 699014 90950 699066
rect 91002 699014 91014 699066
rect 91066 699014 91078 699066
rect 91130 699014 91142 699066
rect 91194 699014 91206 699066
rect 91258 699014 91270 699066
rect 91322 699014 91334 699066
rect 91386 699014 126822 699066
rect 126874 699014 126886 699066
rect 126938 699014 126950 699066
rect 127002 699014 127014 699066
rect 127066 699014 127078 699066
rect 127130 699014 127142 699066
rect 127194 699014 127206 699066
rect 127258 699014 127270 699066
rect 127322 699014 127334 699066
rect 127386 699014 162822 699066
rect 162874 699014 162886 699066
rect 162938 699014 162950 699066
rect 163002 699014 163014 699066
rect 163066 699014 163078 699066
rect 163130 699014 163142 699066
rect 163194 699014 163206 699066
rect 163258 699014 163270 699066
rect 163322 699014 163334 699066
rect 163386 699014 198822 699066
rect 198874 699014 198886 699066
rect 198938 699014 198950 699066
rect 199002 699014 199014 699066
rect 199066 699014 199078 699066
rect 199130 699014 199142 699066
rect 199194 699014 199206 699066
rect 199258 699014 199270 699066
rect 199322 699014 199334 699066
rect 199386 699014 234822 699066
rect 234874 699014 234886 699066
rect 234938 699014 234950 699066
rect 235002 699014 235014 699066
rect 235066 699014 235078 699066
rect 235130 699014 235142 699066
rect 235194 699014 235206 699066
rect 235258 699014 235270 699066
rect 235322 699014 235334 699066
rect 235386 699014 270822 699066
rect 270874 699014 270886 699066
rect 270938 699014 270950 699066
rect 271002 699014 271014 699066
rect 271066 699014 271078 699066
rect 271130 699014 271142 699066
rect 271194 699014 271206 699066
rect 271258 699014 271270 699066
rect 271322 699014 271334 699066
rect 271386 699014 306822 699066
rect 306874 699014 306886 699066
rect 306938 699014 306950 699066
rect 307002 699014 307014 699066
rect 307066 699014 307078 699066
rect 307130 699014 307142 699066
rect 307194 699014 307206 699066
rect 307258 699014 307270 699066
rect 307322 699014 307334 699066
rect 307386 699014 342822 699066
rect 342874 699014 342886 699066
rect 342938 699014 342950 699066
rect 343002 699014 343014 699066
rect 343066 699014 343078 699066
rect 343130 699014 343142 699066
rect 343194 699014 343206 699066
rect 343258 699014 343270 699066
rect 343322 699014 343334 699066
rect 343386 699014 378822 699066
rect 378874 699014 378886 699066
rect 378938 699014 378950 699066
rect 379002 699014 379014 699066
rect 379066 699014 379078 699066
rect 379130 699014 379142 699066
rect 379194 699014 379206 699066
rect 379258 699014 379270 699066
rect 379322 699014 379334 699066
rect 379386 699014 414822 699066
rect 414874 699014 414886 699066
rect 414938 699014 414950 699066
rect 415002 699014 415014 699066
rect 415066 699014 415078 699066
rect 415130 699014 415142 699066
rect 415194 699014 415206 699066
rect 415258 699014 415270 699066
rect 415322 699014 415334 699066
rect 415386 699014 450822 699066
rect 450874 699014 450886 699066
rect 450938 699014 450950 699066
rect 451002 699014 451014 699066
rect 451066 699014 451078 699066
rect 451130 699014 451142 699066
rect 451194 699014 451206 699066
rect 451258 699014 451270 699066
rect 451322 699014 451334 699066
rect 451386 699014 486822 699066
rect 486874 699014 486886 699066
rect 486938 699014 486950 699066
rect 487002 699014 487014 699066
rect 487066 699014 487078 699066
rect 487130 699014 487142 699066
rect 487194 699014 487206 699066
rect 487258 699014 487270 699066
rect 487322 699014 487334 699066
rect 487386 699014 522822 699066
rect 522874 699014 522886 699066
rect 522938 699014 522950 699066
rect 523002 699014 523014 699066
rect 523066 699014 523078 699066
rect 523130 699014 523142 699066
rect 523194 699014 523206 699066
rect 523258 699014 523270 699066
rect 523322 699014 523334 699066
rect 523386 699014 558822 699066
rect 558874 699014 558886 699066
rect 558938 699014 558950 699066
rect 559002 699014 559014 699066
rect 559066 699014 559078 699066
rect 559130 699014 559142 699066
rect 559194 699014 559206 699066
rect 559258 699014 559270 699066
rect 559322 699014 559334 699066
rect 559386 699014 582820 699066
rect 1104 698992 582820 699014
rect 48130 698912 48136 698964
rect 48188 698952 48194 698964
rect 119706 698952 119712 698964
rect 48188 698924 119712 698952
rect 48188 698912 48194 698924
rect 119706 698912 119712 698924
rect 119764 698912 119770 698964
rect 128630 698912 128636 698964
rect 128688 698952 128694 698964
rect 576578 698952 576584 698964
rect 128688 698924 576584 698952
rect 128688 698912 128694 698924
rect 576578 698912 576584 698924
rect 576636 698912 576642 698964
rect 119154 698844 119160 698896
rect 119212 698884 119218 698896
rect 253750 698884 253756 698896
rect 119212 698856 253756 698884
rect 119212 698844 119218 698856
rect 253750 698844 253756 698856
rect 253808 698844 253814 698896
rect 253842 698844 253848 698896
rect 253900 698884 253906 698896
rect 263594 698884 263600 698896
rect 253900 698856 263600 698884
rect 253900 698844 253906 698856
rect 263594 698844 263600 698856
rect 263652 698844 263658 698896
rect 263686 698844 263692 698896
rect 263744 698884 263750 698896
rect 306374 698884 306380 698896
rect 263744 698856 306380 698884
rect 263744 698844 263750 698856
rect 306374 698844 306380 698856
rect 306432 698844 306438 698896
rect 306469 698887 306527 698893
rect 306469 698853 306481 698887
rect 306515 698884 306527 698887
rect 325513 698887 325571 698893
rect 325513 698884 325525 698887
rect 306515 698856 325525 698884
rect 306515 698853 306527 698856
rect 306469 698847 306527 698853
rect 325513 698853 325525 698856
rect 325559 698853 325571 698887
rect 325513 698847 325571 698853
rect 325602 698844 325608 698896
rect 325660 698884 325666 698896
rect 340690 698884 340696 698896
rect 325660 698856 340696 698884
rect 325660 698844 325666 698856
rect 340690 698844 340696 698856
rect 340748 698844 340754 698896
rect 340785 698887 340843 698893
rect 340785 698853 340797 698887
rect 340831 698884 340843 698887
rect 354493 698887 354551 698893
rect 354493 698884 354505 698887
rect 340831 698856 354505 698884
rect 340831 698853 340843 698856
rect 340785 698847 340843 698853
rect 354493 698853 354505 698856
rect 354539 698853 354551 698887
rect 354493 698847 354551 698853
rect 354582 698844 354588 698896
rect 354640 698884 354646 698896
rect 577682 698884 577688 698896
rect 354640 698856 577688 698884
rect 354640 698844 354646 698856
rect 577682 698844 577688 698856
rect 577740 698844 577746 698896
rect 5258 698776 5264 698828
rect 5316 698816 5322 698828
rect 474182 698816 474188 698828
rect 5316 698788 474188 698816
rect 5316 698776 5322 698788
rect 474182 698776 474188 698788
rect 474240 698776 474246 698828
rect 33962 698708 33968 698760
rect 34020 698748 34026 698760
rect 89714 698748 89720 698760
rect 34020 698720 89720 698748
rect 34020 698708 34026 698720
rect 89714 698708 89720 698720
rect 89772 698708 89778 698760
rect 104986 698708 104992 698760
rect 105044 698748 105050 698760
rect 577590 698748 577596 698760
rect 105044 698720 577596 698748
rect 105044 698708 105050 698720
rect 577590 698708 577596 698720
rect 577648 698708 577654 698760
rect 4982 698640 4988 698692
rect 5040 698680 5046 698692
rect 488350 698680 488356 698692
rect 5040 698652 488356 698680
rect 5040 698640 5046 698652
rect 488350 698640 488356 698652
rect 488408 698640 488414 698692
rect 90726 698572 90732 698624
rect 90784 698612 90790 698624
rect 576394 698612 576400 698624
rect 90784 698584 576400 698612
rect 90784 698572 90790 698584
rect 576394 698572 576400 698584
rect 576452 698572 576458 698624
rect 1104 698522 582820 698544
rect 1104 698470 36822 698522
rect 36874 698470 36886 698522
rect 36938 698470 36950 698522
rect 37002 698470 37014 698522
rect 37066 698470 37078 698522
rect 37130 698470 37142 698522
rect 37194 698470 37206 698522
rect 37258 698470 37270 698522
rect 37322 698470 37334 698522
rect 37386 698470 72822 698522
rect 72874 698470 72886 698522
rect 72938 698470 72950 698522
rect 73002 698470 73014 698522
rect 73066 698470 73078 698522
rect 73130 698470 73142 698522
rect 73194 698470 73206 698522
rect 73258 698470 73270 698522
rect 73322 698470 73334 698522
rect 73386 698470 108822 698522
rect 108874 698470 108886 698522
rect 108938 698470 108950 698522
rect 109002 698470 109014 698522
rect 109066 698470 109078 698522
rect 109130 698470 109142 698522
rect 109194 698470 109206 698522
rect 109258 698470 109270 698522
rect 109322 698470 109334 698522
rect 109386 698470 144822 698522
rect 144874 698470 144886 698522
rect 144938 698470 144950 698522
rect 145002 698470 145014 698522
rect 145066 698470 145078 698522
rect 145130 698470 145142 698522
rect 145194 698470 145206 698522
rect 145258 698470 145270 698522
rect 145322 698470 145334 698522
rect 145386 698470 180822 698522
rect 180874 698470 180886 698522
rect 180938 698470 180950 698522
rect 181002 698470 181014 698522
rect 181066 698470 181078 698522
rect 181130 698470 181142 698522
rect 181194 698470 181206 698522
rect 181258 698470 181270 698522
rect 181322 698470 181334 698522
rect 181386 698470 216822 698522
rect 216874 698470 216886 698522
rect 216938 698470 216950 698522
rect 217002 698470 217014 698522
rect 217066 698470 217078 698522
rect 217130 698470 217142 698522
rect 217194 698470 217206 698522
rect 217258 698470 217270 698522
rect 217322 698470 217334 698522
rect 217386 698470 252822 698522
rect 252874 698470 252886 698522
rect 252938 698470 252950 698522
rect 253002 698470 253014 698522
rect 253066 698470 253078 698522
rect 253130 698470 253142 698522
rect 253194 698470 253206 698522
rect 253258 698470 253270 698522
rect 253322 698470 253334 698522
rect 253386 698470 288822 698522
rect 288874 698470 288886 698522
rect 288938 698470 288950 698522
rect 289002 698470 289014 698522
rect 289066 698470 289078 698522
rect 289130 698470 289142 698522
rect 289194 698470 289206 698522
rect 289258 698470 289270 698522
rect 289322 698470 289334 698522
rect 289386 698470 324822 698522
rect 324874 698470 324886 698522
rect 324938 698470 324950 698522
rect 325002 698470 325014 698522
rect 325066 698470 325078 698522
rect 325130 698470 325142 698522
rect 325194 698470 325206 698522
rect 325258 698470 325270 698522
rect 325322 698470 325334 698522
rect 325386 698470 360822 698522
rect 360874 698470 360886 698522
rect 360938 698470 360950 698522
rect 361002 698470 361014 698522
rect 361066 698470 361078 698522
rect 361130 698470 361142 698522
rect 361194 698470 361206 698522
rect 361258 698470 361270 698522
rect 361322 698470 361334 698522
rect 361386 698470 396822 698522
rect 396874 698470 396886 698522
rect 396938 698470 396950 698522
rect 397002 698470 397014 698522
rect 397066 698470 397078 698522
rect 397130 698470 397142 698522
rect 397194 698470 397206 698522
rect 397258 698470 397270 698522
rect 397322 698470 397334 698522
rect 397386 698470 432822 698522
rect 432874 698470 432886 698522
rect 432938 698470 432950 698522
rect 433002 698470 433014 698522
rect 433066 698470 433078 698522
rect 433130 698470 433142 698522
rect 433194 698470 433206 698522
rect 433258 698470 433270 698522
rect 433322 698470 433334 698522
rect 433386 698470 468822 698522
rect 468874 698470 468886 698522
rect 468938 698470 468950 698522
rect 469002 698470 469014 698522
rect 469066 698470 469078 698522
rect 469130 698470 469142 698522
rect 469194 698470 469206 698522
rect 469258 698470 469270 698522
rect 469322 698470 469334 698522
rect 469386 698470 504822 698522
rect 504874 698470 504886 698522
rect 504938 698470 504950 698522
rect 505002 698470 505014 698522
rect 505066 698470 505078 698522
rect 505130 698470 505142 698522
rect 505194 698470 505206 698522
rect 505258 698470 505270 698522
rect 505322 698470 505334 698522
rect 505386 698470 540822 698522
rect 540874 698470 540886 698522
rect 540938 698470 540950 698522
rect 541002 698470 541014 698522
rect 541066 698470 541078 698522
rect 541130 698470 541142 698522
rect 541194 698470 541206 698522
rect 541258 698470 541270 698522
rect 541322 698470 541334 698522
rect 541386 698470 576822 698522
rect 576874 698470 576886 698522
rect 576938 698470 576950 698522
rect 577002 698470 577014 698522
rect 577066 698470 577078 698522
rect 577130 698470 577142 698522
rect 577194 698470 577206 698522
rect 577258 698470 577270 698522
rect 577322 698470 577334 698522
rect 577386 698470 582820 698522
rect 1104 698448 582820 698470
rect 76558 698368 76564 698420
rect 76616 698408 76622 698420
rect 578878 698408 578884 698420
rect 76616 698380 578884 698408
rect 76616 698368 76622 698380
rect 578878 698368 578884 698380
rect 578936 698368 578942 698420
rect 62298 698300 62304 698352
rect 62356 698340 62362 698352
rect 576302 698340 576308 698352
rect 62356 698312 576308 698340
rect 62356 698300 62362 698312
rect 576302 698300 576308 698312
rect 576360 698300 576366 698352
rect 5718 698232 5724 698284
rect 5776 698272 5782 698284
rect 351086 698272 351092 698284
rect 5776 698244 351092 698272
rect 5776 698232 5782 698244
rect 351086 698232 351092 698244
rect 351144 698232 351150 698284
rect 354677 698275 354735 698281
rect 354677 698241 354689 698275
rect 354723 698272 354735 698275
rect 354723 698244 365392 698272
rect 354723 698241 354735 698244
rect 354677 698235 354735 698241
rect 5810 698164 5816 698216
rect 5868 698204 5874 698216
rect 365254 698204 365260 698216
rect 5868 698176 365260 698204
rect 5868 698164 5874 698176
rect 365254 698164 365260 698176
rect 365312 698164 365318 698216
rect 365364 698204 365392 698244
rect 580626 698204 580632 698216
rect 365364 698176 580632 698204
rect 580626 698164 580632 698176
rect 580684 698164 580690 698216
rect 209038 698096 209044 698148
rect 209096 698136 209102 698148
rect 574554 698136 574560 698148
rect 209096 698108 574560 698136
rect 209096 698096 209102 698108
rect 574554 698096 574560 698108
rect 574612 698096 574618 698148
rect 5902 698028 5908 698080
rect 5960 698068 5966 698080
rect 5960 698040 6132 698068
rect 5960 698028 5966 698040
rect 6104 698000 6132 698040
rect 213822 698028 213828 698080
rect 213880 698068 213886 698080
rect 579614 698068 579620 698080
rect 213880 698040 579620 698068
rect 213880 698028 213886 698040
rect 579614 698028 579620 698040
rect 579672 698028 579678 698080
rect 379514 698000 379520 698012
rect 1104 697904 6000 698000
rect 6104 697972 379520 698000
rect 379514 697960 379520 697972
rect 379572 697960 379578 698012
rect 194870 697892 194876 697944
rect 194928 697932 194934 697944
rect 574646 697932 574652 697944
rect 194928 697904 574652 697932
rect 194928 697892 194934 697904
rect 574646 697892 574652 697904
rect 574704 697892 574710 697944
rect 578000 697904 582820 698000
rect 5994 697824 6000 697876
rect 6052 697864 6058 697876
rect 393682 697864 393688 697876
rect 6052 697836 393688 697864
rect 6052 697824 6058 697836
rect 393682 697824 393688 697836
rect 393740 697824 393746 697876
rect 7374 697756 7380 697808
rect 7432 697796 7438 697808
rect 398374 697796 398380 697808
rect 7432 697768 398380 697796
rect 7432 697756 7438 697768
rect 398374 697756 398380 697768
rect 398432 697756 398438 697808
rect 180702 697688 180708 697740
rect 180760 697728 180766 697740
rect 575382 697728 575388 697740
rect 180760 697700 575388 697728
rect 180760 697688 180766 697700
rect 575382 697688 575388 697700
rect 575440 697688 575446 697740
rect 6086 697620 6092 697672
rect 6144 697660 6150 697672
rect 407850 697660 407856 697672
rect 6144 697632 407856 697660
rect 6144 697620 6150 697632
rect 407850 697620 407856 697632
rect 407908 697620 407914 697672
rect 407942 697620 407948 697672
rect 408000 697660 408006 697672
rect 580810 697660 580816 697672
rect 408000 697632 580816 697660
rect 408000 697620 408006 697632
rect 580810 697620 580816 697632
rect 580868 697620 580874 697672
rect 166442 697552 166448 697604
rect 166500 697592 166506 697604
rect 577958 697592 577964 697604
rect 166500 697564 577964 697592
rect 166500 697552 166506 697564
rect 577958 697552 577964 697564
rect 578016 697552 578022 697604
rect 6730 697484 6736 697536
rect 6788 697524 6794 697536
rect 422110 697524 422116 697536
rect 6788 697496 422116 697524
rect 6788 697484 6794 697496
rect 422110 697484 422116 697496
rect 422168 697484 422174 697536
rect 1104 697360 6000 697456
rect 152274 697416 152280 697468
rect 152332 697456 152338 697468
rect 576762 697456 576768 697468
rect 152332 697428 576768 697456
rect 152332 697416 152338 697428
rect 576762 697416 576768 697428
rect 576820 697416 576826 697468
rect 6638 697348 6644 697400
rect 6696 697388 6702 697400
rect 436278 697388 436284 697400
rect 6696 697360 436284 697388
rect 6696 697348 6702 697360
rect 436278 697348 436284 697360
rect 436336 697348 436342 697400
rect 578000 697360 582820 697456
rect 6454 697280 6460 697332
rect 6512 697320 6518 697332
rect 455230 697320 455236 697332
rect 6512 697292 455236 697320
rect 6512 697280 6518 697292
rect 455230 697280 455236 697292
rect 455288 697280 455294 697332
rect 6362 697212 6368 697264
rect 6420 697252 6426 697264
rect 464706 697252 464712 697264
rect 6420 697224 464712 697252
rect 6420 697212 6426 697224
rect 464706 697212 464712 697224
rect 464764 697212 464770 697264
rect 7926 697144 7932 697196
rect 7984 697184 7990 697196
rect 493042 697184 493048 697196
rect 7984 697156 493048 697184
rect 7984 697144 7990 697156
rect 493042 697144 493048 697156
rect 493100 697144 493106 697196
rect 7558 697076 7564 697128
rect 7616 697116 7622 697128
rect 535638 697116 535644 697128
rect 7616 697088 535644 697116
rect 7616 697076 7622 697088
rect 535638 697076 535644 697088
rect 535696 697076 535702 697128
rect 38654 697008 38660 697060
rect 38712 697048 38718 697060
rect 574922 697048 574928 697060
rect 38712 697020 574928 697048
rect 38712 697008 38718 697020
rect 574922 697008 574928 697020
rect 574980 697008 574986 697060
rect 24486 696940 24492 696992
rect 24544 696980 24550 696992
rect 576210 696980 576216 696992
rect 24544 696952 576216 696980
rect 24544 696940 24550 696952
rect 576210 696940 576216 696952
rect 576268 696940 576274 696992
rect 224957 696915 225015 696921
rect 1104 696816 6000 696912
rect 224957 696881 224969 696915
rect 225003 696912 225015 696915
rect 234525 696915 234583 696921
rect 234525 696912 234537 696915
rect 225003 696884 234537 696912
rect 225003 696881 225015 696884
rect 224957 696875 225015 696881
rect 234525 696881 234537 696884
rect 234571 696881 234583 696915
rect 234525 696875 234583 696881
rect 244277 696915 244335 696921
rect 244277 696881 244289 696915
rect 244323 696912 244335 696915
rect 253845 696915 253903 696921
rect 253845 696912 253857 696915
rect 244323 696884 253857 696912
rect 244323 696881 244335 696884
rect 244277 696875 244335 696881
rect 253845 696881 253857 696884
rect 253891 696881 253903 696915
rect 253845 696875 253903 696881
rect 263597 696915 263655 696921
rect 263597 696881 263609 696915
rect 263643 696912 263655 696915
rect 273165 696915 273223 696921
rect 273165 696912 273177 696915
rect 263643 696884 273177 696912
rect 263643 696881 263655 696884
rect 263597 696875 263655 696881
rect 273165 696881 273177 696884
rect 273211 696881 273223 696915
rect 273165 696875 273223 696881
rect 282917 696915 282975 696921
rect 282917 696881 282929 696915
rect 282963 696912 282975 696915
rect 292485 696915 292543 696921
rect 292485 696912 292497 696915
rect 282963 696884 292497 696912
rect 282963 696881 282975 696884
rect 282917 696875 282975 696881
rect 292485 696881 292497 696884
rect 292531 696881 292543 696915
rect 292485 696875 292543 696881
rect 297269 696915 297327 696921
rect 297269 696881 297281 696915
rect 297315 696912 297327 696915
rect 306929 696915 306987 696921
rect 306929 696912 306941 696915
rect 297315 696884 306941 696912
rect 297315 696881 297327 696884
rect 297269 696875 297327 696881
rect 306929 696881 306941 696884
rect 306975 696881 306987 696915
rect 306929 696875 306987 696881
rect 355229 696915 355287 696921
rect 355229 696881 355241 696915
rect 355275 696912 355287 696915
rect 362129 696915 362187 696921
rect 362129 696912 362141 696915
rect 355275 696884 362141 696912
rect 355275 696881 355287 696884
rect 355229 696875 355287 696881
rect 362129 696881 362141 696884
rect 362175 696881 362187 696915
rect 362129 696875 362187 696881
rect 373994 696872 374000 696924
rect 374052 696912 374058 696924
rect 374822 696912 374828 696924
rect 374052 696884 374828 696912
rect 374052 696872 374058 696884
rect 374822 696872 374828 696884
rect 374880 696872 374886 696924
rect 289722 696844 289728 696856
rect 6104 696816 289728 696844
rect 3970 696736 3976 696788
rect 4028 696776 4034 696788
rect 6104 696776 6132 696816
rect 289722 696804 289728 696816
rect 289780 696804 289786 696856
rect 297361 696847 297419 696853
rect 297361 696813 297373 696847
rect 297407 696844 297419 696847
rect 307021 696847 307079 696853
rect 307021 696844 307033 696847
rect 297407 696816 307033 696844
rect 297407 696813 297419 696816
rect 297361 696807 297419 696813
rect 307021 696813 307033 696816
rect 307067 696813 307079 696847
rect 307021 696807 307079 696813
rect 355321 696847 355379 696853
rect 355321 696813 355333 696847
rect 355367 696844 355379 696847
rect 364981 696847 365039 696853
rect 364981 696844 364993 696847
rect 355367 696816 364993 696844
rect 355367 696813 355379 696816
rect 355321 696807 355379 696813
rect 364981 696813 364993 696816
rect 365027 696813 365039 696847
rect 364981 696807 365039 696813
rect 374641 696847 374699 696853
rect 374641 696813 374653 696847
rect 374687 696844 374699 696847
rect 384301 696847 384359 696853
rect 384301 696844 384313 696847
rect 374687 696816 384313 696844
rect 374687 696813 374699 696816
rect 374641 696807 374699 696813
rect 384301 696813 384313 696816
rect 384347 696813 384359 696847
rect 578000 696816 582820 696912
rect 384301 696807 384359 696813
rect 4028 696748 6132 696776
rect 6181 696779 6239 696785
rect 4028 696736 4034 696748
rect 6181 696745 6193 696779
rect 6227 696776 6239 696779
rect 404262 696776 404268 696788
rect 6227 696748 404268 696776
rect 6227 696745 6239 696748
rect 6181 696739 6239 696745
rect 404262 696736 404268 696748
rect 404320 696736 404326 696788
rect 4706 696668 4712 696720
rect 4764 696708 4770 696720
rect 360562 696708 360568 696720
rect 4764 696680 360568 696708
rect 4764 696668 4770 696680
rect 360562 696668 360568 696680
rect 360620 696668 360626 696720
rect 372249 696711 372307 696717
rect 372249 696677 372261 696711
rect 372295 696708 372307 696711
rect 388990 696708 388996 696720
rect 372295 696680 388996 696708
rect 372295 696677 372307 696680
rect 372249 696671 372307 696677
rect 388990 696668 388996 696680
rect 389048 696668 389054 696720
rect 3326 696600 3332 696652
rect 3384 696640 3390 696652
rect 6181 696643 6239 696649
rect 6181 696640 6193 696643
rect 3384 696612 6193 696640
rect 3384 696600 3390 696612
rect 6181 696609 6193 696612
rect 6227 696609 6239 696643
rect 6181 696603 6239 696609
rect 86957 696643 87015 696649
rect 86957 696609 86969 696643
rect 87003 696640 87015 696643
rect 96525 696643 96583 696649
rect 96525 696640 96537 696643
rect 87003 696612 96537 696640
rect 87003 696609 87015 696612
rect 86957 696603 87015 696609
rect 96525 696609 96537 696612
rect 96571 696609 96583 696643
rect 96525 696603 96583 696609
rect 205637 696643 205695 696649
rect 205637 696609 205649 696643
rect 205683 696640 205695 696643
rect 215205 696643 215263 696649
rect 215205 696640 215217 696643
rect 205683 696612 215217 696640
rect 205683 696609 205695 696612
rect 205637 696603 205695 696609
rect 215205 696609 215217 696612
rect 215251 696609 215263 696643
rect 215205 696603 215263 696609
rect 218514 696600 218520 696652
rect 218572 696640 218578 696652
rect 578786 696640 578792 696652
rect 218572 696612 578792 696640
rect 218572 696600 218578 696612
rect 578786 696600 578792 696612
rect 578844 696600 578850 696652
rect 5442 696532 5448 696584
rect 5500 696572 5506 696584
rect 374730 696572 374736 696584
rect 5500 696544 374736 696572
rect 5500 696532 5506 696544
rect 374730 696532 374736 696544
rect 374788 696532 374794 696584
rect 374822 696532 374828 696584
rect 374880 696572 374886 696584
rect 580718 696572 580724 696584
rect 374880 696544 580724 696572
rect 374880 696532 374886 696544
rect 580718 696532 580724 696544
rect 580776 696532 580782 696584
rect 154577 696507 154635 696513
rect 154577 696473 154589 696507
rect 154623 696504 154635 696507
rect 163869 696507 163927 696513
rect 163869 696504 163881 696507
rect 154623 696476 163881 696504
rect 154623 696473 154635 696476
rect 154577 696467 154635 696473
rect 163869 696473 163881 696476
rect 163915 696473 163927 696507
rect 163869 696467 163927 696473
rect 173897 696507 173955 696513
rect 173897 696473 173909 696507
rect 173943 696504 173955 696507
rect 178681 696507 178739 696513
rect 178681 696504 178693 696507
rect 173943 696476 178693 696504
rect 173943 696473 173955 696476
rect 173897 696467 173955 696473
rect 178681 696473 178693 696476
rect 178727 696473 178739 696507
rect 178681 696467 178739 696473
rect 186317 696507 186375 696513
rect 186317 696473 186329 696507
rect 186363 696504 186375 696507
rect 186363 696476 200804 696504
rect 186363 696473 186375 696476
rect 186317 696467 186375 696473
rect 22189 696439 22247 696445
rect 22189 696405 22201 696439
rect 22235 696436 22247 696439
rect 60829 696439 60887 696445
rect 22235 696408 46888 696436
rect 22235 696405 22247 696408
rect 22189 696399 22247 696405
rect 6089 696371 6147 696377
rect 1104 696272 6000 696368
rect 6089 696337 6101 696371
rect 6135 696368 6147 696371
rect 22005 696371 22063 696377
rect 22005 696368 22017 696371
rect 6135 696340 22017 696368
rect 6135 696337 6147 696340
rect 6089 696331 6147 696337
rect 22005 696337 22017 696340
rect 22051 696337 22063 696371
rect 22005 696331 22063 696337
rect 46860 696300 46888 696408
rect 60829 696405 60841 696439
rect 60875 696436 60887 696439
rect 67637 696439 67695 696445
rect 67637 696436 67649 696439
rect 60875 696408 67649 696436
rect 60875 696405 60887 696408
rect 60829 696399 60887 696405
rect 67637 696405 67649 696408
rect 67683 696405 67695 696439
rect 67637 696399 67695 696405
rect 80149 696439 80207 696445
rect 80149 696405 80161 696439
rect 80195 696436 80207 696439
rect 86957 696439 87015 696445
rect 86957 696436 86969 696439
rect 80195 696408 86969 696436
rect 80195 696405 80207 696408
rect 80149 696399 80207 696405
rect 86957 696405 86969 696408
rect 87003 696405 87015 696439
rect 86957 696399 87015 696405
rect 99377 696439 99435 696445
rect 99377 696405 99389 696439
rect 99423 696436 99435 696439
rect 108945 696439 109003 696445
rect 108945 696436 108957 696439
rect 99423 696408 108957 696436
rect 99423 696405 99435 696408
rect 99377 696399 99435 696405
rect 108945 696405 108957 696408
rect 108991 696405 109003 696439
rect 108945 696399 109003 696405
rect 115845 696439 115903 696445
rect 115845 696405 115857 696439
rect 115891 696436 115903 696439
rect 115891 696408 118740 696436
rect 115891 696405 115903 696408
rect 115845 696399 115903 696405
rect 60645 696371 60703 696377
rect 60645 696368 60657 696371
rect 46952 696340 60657 696368
rect 46952 696300 46980 696340
rect 60645 696337 60657 696340
rect 60691 696337 60703 696371
rect 60645 696331 60703 696337
rect 77205 696371 77263 696377
rect 77205 696337 77217 696371
rect 77251 696368 77263 696371
rect 79965 696371 80023 696377
rect 79965 696368 79977 696371
rect 77251 696340 79977 696368
rect 77251 696337 77263 696340
rect 77205 696331 77263 696337
rect 79965 696337 79977 696340
rect 80011 696337 80023 696371
rect 79965 696331 80023 696337
rect 96525 696371 96583 696377
rect 96525 696337 96537 696371
rect 96571 696368 96583 696371
rect 99285 696371 99343 696377
rect 99285 696368 99297 696371
rect 96571 696340 99297 696368
rect 96571 696337 96583 696340
rect 96525 696331 96583 696337
rect 99285 696337 99297 696340
rect 99331 696337 99343 696371
rect 99285 696331 99343 696337
rect 46860 696272 46980 696300
rect 108945 696303 109003 696309
rect 108945 696269 108957 696303
rect 108991 696300 109003 696303
rect 115845 696303 115903 696309
rect 115845 696300 115857 696303
rect 108991 696272 115857 696300
rect 108991 696269 109003 696272
rect 108945 696263 109003 696269
rect 115845 696269 115857 696272
rect 115891 696269 115903 696303
rect 118712 696300 118740 696408
rect 119706 696396 119712 696448
rect 119764 696436 119770 696448
rect 164053 696439 164111 696445
rect 164053 696436 164065 696439
rect 119764 696408 164065 696436
rect 119764 696396 119770 696408
rect 164053 696405 164065 696408
rect 164099 696405 164111 696439
rect 164053 696399 164111 696405
rect 164237 696439 164295 696445
rect 164237 696405 164249 696439
rect 164283 696436 164295 696439
rect 200669 696439 200727 696445
rect 200669 696436 200681 696439
rect 164283 696408 200681 696436
rect 164283 696405 164295 696408
rect 164237 696399 164295 696405
rect 200669 696405 200681 696408
rect 200715 696405 200727 696439
rect 200669 696399 200727 696405
rect 138109 696371 138167 696377
rect 138109 696337 138121 696371
rect 138155 696368 138167 696371
rect 143537 696371 143595 696377
rect 143537 696368 143549 696371
rect 138155 696340 143549 696368
rect 138155 696337 138167 696340
rect 138109 696331 138167 696337
rect 143537 696337 143549 696340
rect 143583 696337 143595 696371
rect 143537 696331 143595 696337
rect 171594 696328 171600 696380
rect 171652 696368 171658 696380
rect 178681 696371 178739 696377
rect 171652 696340 171697 696368
rect 171652 696328 171658 696340
rect 178681 696337 178693 696371
rect 178727 696368 178739 696371
rect 186317 696371 186375 696377
rect 186317 696368 186329 696371
rect 178727 696340 186329 696368
rect 178727 696337 178739 696340
rect 178681 696331 178739 696337
rect 186317 696337 186329 696340
rect 186363 696337 186375 696371
rect 200776 696368 200804 696476
rect 204346 696464 204352 696516
rect 204404 696504 204410 696516
rect 579522 696504 579528 696516
rect 204404 696476 579528 696504
rect 204404 696464 204410 696476
rect 579522 696464 579528 696476
rect 579580 696464 579586 696516
rect 200853 696439 200911 696445
rect 200853 696405 200865 696439
rect 200899 696436 200911 696439
rect 580442 696436 580448 696448
rect 200899 696408 580448 696436
rect 200899 696405 200911 696408
rect 200853 696399 200911 696405
rect 580442 696396 580448 696408
rect 580500 696396 580506 696448
rect 205637 696371 205695 696377
rect 205637 696368 205649 696371
rect 200776 696340 205649 696368
rect 186317 696331 186375 696337
rect 205637 696337 205649 696340
rect 205683 696337 205695 696371
rect 205637 696331 205695 696337
rect 215205 696371 215263 696377
rect 215205 696337 215217 696371
rect 215251 696368 215263 696371
rect 224957 696371 225015 696377
rect 224957 696368 224969 696371
rect 215251 696340 224969 696368
rect 215251 696337 215263 696340
rect 215205 696331 215263 696337
rect 224957 696337 224969 696340
rect 225003 696337 225015 696371
rect 224957 696331 225015 696337
rect 234525 696371 234583 696377
rect 234525 696337 234537 696371
rect 234571 696368 234583 696371
rect 244277 696371 244335 696377
rect 244277 696368 244289 696371
rect 234571 696340 244289 696368
rect 234571 696337 234583 696340
rect 234525 696331 234583 696337
rect 244277 696337 244289 696340
rect 244323 696337 244335 696371
rect 244277 696331 244335 696337
rect 253845 696371 253903 696377
rect 253845 696337 253857 696371
rect 253891 696368 253903 696371
rect 263597 696371 263655 696377
rect 263597 696368 263609 696371
rect 253891 696340 263609 696368
rect 253891 696337 253903 696340
rect 253845 696331 253903 696337
rect 263597 696337 263609 696340
rect 263643 696337 263655 696371
rect 263597 696331 263655 696337
rect 273165 696371 273223 696377
rect 273165 696337 273177 696371
rect 273211 696368 273223 696371
rect 282917 696371 282975 696377
rect 282917 696368 282929 696371
rect 273211 696340 282929 696368
rect 273211 696337 273223 696340
rect 273165 696331 273223 696337
rect 282917 696337 282929 696340
rect 282963 696337 282975 696371
rect 282917 696331 282975 696337
rect 292485 696371 292543 696377
rect 292485 696337 292497 696371
rect 292531 696368 292543 696371
rect 297361 696371 297419 696377
rect 297361 696368 297373 696371
rect 292531 696340 297373 696368
rect 292531 696337 292543 696340
rect 292485 696331 292543 696337
rect 297361 696337 297373 696340
rect 297407 696337 297419 696371
rect 297361 696331 297419 696337
rect 307021 696371 307079 696377
rect 307021 696337 307033 696371
rect 307067 696368 307079 696371
rect 355321 696371 355379 696377
rect 355321 696368 355333 696371
rect 307067 696340 355333 696368
rect 307067 696337 307079 696340
rect 307021 696331 307079 696337
rect 355321 696337 355333 696340
rect 355367 696337 355379 696371
rect 355321 696331 355379 696337
rect 364981 696371 365039 696377
rect 364981 696337 364993 696371
rect 365027 696368 365039 696371
rect 372249 696371 372307 696377
rect 372249 696368 372261 696371
rect 365027 696340 372261 696368
rect 365027 696337 365039 696340
rect 364981 696331 365039 696337
rect 372249 696337 372261 696340
rect 372295 696337 372307 696371
rect 372249 696331 372307 696337
rect 393961 696371 394019 696377
rect 393961 696337 393973 696371
rect 394007 696368 394019 696371
rect 403621 696371 403679 696377
rect 403621 696368 403633 696371
rect 394007 696340 403633 696368
rect 394007 696337 394019 696340
rect 393961 696331 394019 696337
rect 403621 696337 403633 696340
rect 403667 696337 403679 696371
rect 403621 696331 403679 696337
rect 132497 696303 132555 696309
rect 132497 696300 132509 696303
rect 118712 696272 132509 696300
rect 115845 696263 115903 696269
rect 132497 696269 132509 696272
rect 132543 696269 132555 696303
rect 132497 696263 132555 696269
rect 143629 696303 143687 696309
rect 143629 696269 143641 696303
rect 143675 696300 143687 696303
rect 154577 696303 154635 696309
rect 154577 696300 154589 696303
rect 143675 696272 154589 696300
rect 143675 696269 143687 696272
rect 143629 696263 143687 696269
rect 154577 696269 154589 696272
rect 154623 696269 154635 696303
rect 154577 696263 154635 696269
rect 163869 696303 163927 696309
rect 163869 696269 163881 696303
rect 163915 696300 163927 696303
rect 173897 696303 173955 696309
rect 173897 696300 173909 696303
rect 163915 696272 173909 696300
rect 163915 696269 163927 696272
rect 163869 696263 163927 696269
rect 173897 696269 173909 696272
rect 173943 696269 173955 696303
rect 173897 696263 173955 696269
rect 190178 696260 190184 696312
rect 190236 696300 190242 696312
rect 567013 696303 567071 696309
rect 567013 696300 567025 696303
rect 190236 696272 567025 696300
rect 190236 696260 190242 696272
rect 567013 696269 567025 696272
rect 567059 696269 567071 696303
rect 578000 696272 582820 696368
rect 567013 696263 567071 696269
rect 67637 696235 67695 696241
rect 67637 696201 67649 696235
rect 67683 696232 67695 696235
rect 77205 696235 77263 696241
rect 77205 696232 77217 696235
rect 67683 696204 77217 696232
rect 67683 696201 67695 696204
rect 67637 696195 67695 696201
rect 77205 696201 77217 696204
rect 77251 696201 77263 696235
rect 77205 696195 77263 696201
rect 89714 696192 89720 696244
rect 89772 696232 89778 696244
rect 154669 696235 154727 696241
rect 154669 696232 154681 696235
rect 89772 696204 154681 696232
rect 89772 696192 89778 696204
rect 154669 696201 154681 696204
rect 154715 696201 154727 696235
rect 154669 696195 154727 696201
rect 154761 696235 154819 696241
rect 154761 696201 154773 696235
rect 154807 696232 154819 696235
rect 173989 696235 174047 696241
rect 173989 696232 174001 696235
rect 154807 696204 174001 696232
rect 154807 696201 154819 696204
rect 154761 696195 154819 696201
rect 173989 696201 174001 696204
rect 174035 696201 174047 696235
rect 173989 696195 174047 696201
rect 174081 696235 174139 696241
rect 174081 696201 174093 696235
rect 174127 696232 174139 696235
rect 580258 696232 580264 696244
rect 174127 696204 580264 696232
rect 174127 696201 174139 696204
rect 174081 696195 174139 696201
rect 580258 696192 580264 696204
rect 580316 696192 580322 696244
rect 6822 696124 6828 696176
rect 6880 696164 6886 696176
rect 154577 696167 154635 696173
rect 154577 696164 154589 696167
rect 6880 696136 154589 696164
rect 6880 696124 6886 696136
rect 154577 696133 154589 696136
rect 154623 696133 154635 696167
rect 154577 696127 154635 696133
rect 154945 696167 155003 696173
rect 154945 696133 154957 696167
rect 154991 696164 155003 696167
rect 173894 696164 173900 696176
rect 154991 696136 173900 696164
rect 154991 696133 155003 696136
rect 154945 696127 155003 696133
rect 173894 696124 173900 696136
rect 173952 696124 173958 696176
rect 174354 696124 174360 696176
rect 174412 696164 174418 696176
rect 412634 696164 412640 696176
rect 174412 696136 412640 696164
rect 174412 696124 174418 696136
rect 412634 696124 412640 696136
rect 412692 696124 412698 696176
rect 413281 696167 413339 696173
rect 413281 696133 413293 696167
rect 413327 696164 413339 696167
rect 422941 696167 422999 696173
rect 422941 696164 422953 696167
rect 413327 696136 422953 696164
rect 413327 696133 413339 696136
rect 413281 696127 413339 696133
rect 422941 696133 422953 696136
rect 422987 696133 422999 696167
rect 422941 696127 422999 696133
rect 432325 696167 432383 696173
rect 432325 696133 432337 696167
rect 432371 696164 432383 696167
rect 442261 696167 442319 696173
rect 442261 696164 442273 696167
rect 432371 696136 442273 696164
rect 432371 696133 432383 696136
rect 432325 696127 432383 696133
rect 442261 696133 442273 696136
rect 442307 696133 442319 696167
rect 442261 696127 442319 696133
rect 567013 696167 567071 696173
rect 567013 696133 567025 696167
rect 567059 696164 567071 696167
rect 579430 696164 579436 696176
rect 567059 696136 579436 696164
rect 567059 696133 567071 696136
rect 567013 696127 567071 696133
rect 579430 696124 579436 696136
rect 579488 696124 579494 696176
rect 132497 696099 132555 696105
rect 132497 696065 132509 696099
rect 132543 696096 132555 696099
rect 138109 696099 138167 696105
rect 138109 696096 138121 696099
rect 132543 696068 138121 696096
rect 132543 696065 132555 696068
rect 132497 696059 132555 696065
rect 138109 696065 138121 696068
rect 138155 696065 138167 696099
rect 138109 696059 138167 696065
rect 147582 696056 147588 696108
rect 147640 696096 147646 696108
rect 154669 696099 154727 696105
rect 154669 696096 154681 696099
rect 147640 696068 154681 696096
rect 147640 696056 147646 696068
rect 154669 696065 154681 696068
rect 154715 696065 154727 696099
rect 154669 696059 154727 696065
rect 154853 696099 154911 696105
rect 154853 696065 154865 696099
rect 154899 696096 154911 696099
rect 173989 696099 174047 696105
rect 173989 696096 174001 696099
rect 154899 696068 174001 696096
rect 154899 696065 154911 696068
rect 154853 696059 154911 696065
rect 173989 696065 174001 696068
rect 174035 696065 174047 696099
rect 173989 696059 174047 696065
rect 174173 696099 174231 696105
rect 174173 696065 174185 696099
rect 174219 696096 174231 696099
rect 579246 696096 579252 696108
rect 174219 696068 579252 696096
rect 174219 696065 174231 696068
rect 174173 696059 174231 696065
rect 579246 696056 579252 696068
rect 579304 696056 579310 696108
rect 46201 696031 46259 696037
rect 46201 695997 46213 696031
rect 46247 696028 46259 696031
rect 55861 696031 55919 696037
rect 55861 696028 55873 696031
rect 46247 696000 55873 696028
rect 46247 695997 46259 696000
rect 46201 695991 46259 695997
rect 55861 695997 55873 696000
rect 55907 695997 55919 696031
rect 55861 695991 55919 695997
rect 62761 696031 62819 696037
rect 62761 695997 62773 696031
rect 62807 696028 62819 696031
rect 75181 696031 75239 696037
rect 75181 696028 75193 696031
rect 62807 696000 75193 696028
rect 62807 695997 62819 696000
rect 62761 695991 62819 695997
rect 75181 695997 75193 696000
rect 75227 695997 75239 696031
rect 75181 695991 75239 695997
rect 82081 696031 82139 696037
rect 82081 695997 82093 696031
rect 82127 696028 82139 696031
rect 94501 696031 94559 696037
rect 94501 696028 94513 696031
rect 82127 696000 94513 696028
rect 82127 695997 82139 696000
rect 82081 695991 82139 695997
rect 94501 695997 94513 696000
rect 94547 695997 94559 696031
rect 94501 695991 94559 695997
rect 114557 696031 114615 696037
rect 114557 695997 114569 696031
rect 114603 696028 114615 696031
rect 123941 696031 123999 696037
rect 123941 696028 123953 696031
rect 114603 696000 123953 696028
rect 114603 695997 114615 696000
rect 114557 695991 114615 695997
rect 123941 695997 123953 696000
rect 123987 695997 123999 696031
rect 123941 695991 123999 695997
rect 124030 695988 124036 696040
rect 124088 696028 124094 696040
rect 124125 696031 124183 696037
rect 124125 696028 124137 696031
rect 124088 696000 124137 696028
rect 124088 695988 124094 696000
rect 124125 695997 124137 696000
rect 124171 695997 124183 696031
rect 138474 696028 138480 696040
rect 138435 696000 138480 696028
rect 124125 695991 124183 695997
rect 138474 695988 138480 696000
rect 138532 695988 138538 696040
rect 143074 695988 143080 696040
rect 143132 696028 143138 696040
rect 173894 696028 173900 696040
rect 143132 696000 173900 696028
rect 143132 695988 143138 696000
rect 173894 695988 173900 696000
rect 173952 695988 173958 696040
rect 174262 695988 174268 696040
rect 174320 696028 174326 696040
rect 577774 696028 577780 696040
rect 174320 696000 577780 696028
rect 174320 695988 174326 696000
rect 577774 695988 577780 696000
rect 577832 695988 577838 696040
rect 6546 695920 6552 695972
rect 6604 695960 6610 695972
rect 154669 695963 154727 695969
rect 154669 695960 154681 695963
rect 6604 695932 154681 695960
rect 6604 695920 6610 695932
rect 154669 695929 154681 695932
rect 154715 695929 154727 695963
rect 154669 695923 154727 695929
rect 154853 695963 154911 695969
rect 154853 695929 154865 695963
rect 154899 695960 154911 695963
rect 173989 695963 174047 695969
rect 173989 695960 174001 695963
rect 154899 695932 174001 695960
rect 154899 695929 154911 695932
rect 154853 695923 154911 695929
rect 173989 695929 174001 695932
rect 174035 695929 174047 695963
rect 173989 695923 174047 695929
rect 174173 695963 174231 695969
rect 174173 695929 174185 695963
rect 174219 695960 174231 695963
rect 450078 695960 450084 695972
rect 174219 695932 450084 695960
rect 174219 695929 174231 695932
rect 174173 695923 174231 695929
rect 450078 695920 450084 695932
rect 450136 695920 450142 695972
rect 451277 695963 451335 695969
rect 451277 695929 451289 695963
rect 451323 695960 451335 695963
rect 461397 695963 461455 695969
rect 461397 695960 461409 695963
rect 451323 695932 461409 695960
rect 451323 695929 451335 695932
rect 451277 695923 451335 695929
rect 461397 695929 461409 695932
rect 461443 695929 461455 695963
rect 461397 695923 461455 695929
rect 483017 695963 483075 695969
rect 483017 695929 483029 695963
rect 483063 695960 483075 695963
rect 492585 695963 492643 695969
rect 492585 695960 492597 695963
rect 483063 695932 492597 695960
rect 483063 695929 483075 695932
rect 483017 695923 483075 695929
rect 492585 695929 492597 695932
rect 492631 695929 492643 695963
rect 492585 695923 492643 695929
rect 492677 695963 492735 695969
rect 492677 695929 492689 695963
rect 492723 695960 492735 695963
rect 502245 695963 502303 695969
rect 502245 695960 502257 695963
rect 492723 695932 502257 695960
rect 492723 695929 492735 695932
rect 492677 695923 492735 695929
rect 502245 695929 502257 695932
rect 502291 695929 502303 695963
rect 502245 695923 502303 695929
rect 5074 695852 5080 695904
rect 5132 695892 5138 695904
rect 173897 695895 173955 695901
rect 173897 695892 173909 695895
rect 5132 695864 173909 695892
rect 5132 695852 5138 695864
rect 173897 695861 173909 695864
rect 173943 695861 173955 695895
rect 173897 695855 173955 695861
rect 174265 695895 174323 695901
rect 174265 695861 174277 695895
rect 174311 695892 174323 695895
rect 459646 695892 459652 695904
rect 174311 695864 459652 695892
rect 174311 695861 174323 695864
rect 174265 695855 174323 695861
rect 459646 695852 459652 695864
rect 459704 695852 459710 695904
rect 471241 695895 471299 695901
rect 471241 695861 471253 695895
rect 471287 695892 471299 695895
rect 471287 695864 479656 695892
rect 471287 695861 471299 695864
rect 471241 695855 471299 695861
rect 1104 695728 6000 695824
rect 6270 695784 6276 695836
rect 6328 695824 6334 695836
rect 154577 695827 154635 695833
rect 154577 695824 154589 695827
rect 6328 695796 154589 695824
rect 6328 695784 6334 695796
rect 154577 695793 154589 695796
rect 154623 695793 154635 695827
rect 154577 695787 154635 695793
rect 155037 695827 155095 695833
rect 155037 695793 155049 695827
rect 155083 695824 155095 695827
rect 478782 695824 478788 695836
rect 155083 695796 478788 695824
rect 155083 695793 155095 695796
rect 155037 695787 155095 695793
rect 478782 695784 478788 695796
rect 478840 695784 478846 695836
rect 479628 695824 479656 695864
rect 483017 695827 483075 695833
rect 483017 695824 483029 695827
rect 479628 695796 483029 695824
rect 483017 695793 483029 695796
rect 483063 695793 483075 695827
rect 483017 695787 483075 695793
rect 154669 695759 154727 695765
rect 154669 695756 154681 695759
rect 6104 695728 154681 695756
rect 3694 695648 3700 695700
rect 3752 695688 3758 695700
rect 6104 695688 6132 695728
rect 154669 695725 154681 695728
rect 154715 695725 154727 695759
rect 154669 695719 154727 695725
rect 154945 695759 155003 695765
rect 154945 695725 154957 695759
rect 154991 695756 155003 695759
rect 483382 695756 483388 695768
rect 154991 695728 483388 695756
rect 154991 695725 155003 695728
rect 154945 695719 155003 695725
rect 483382 695716 483388 695728
rect 483440 695716 483446 695768
rect 492585 695759 492643 695765
rect 492585 695725 492597 695759
rect 492631 695756 492643 695759
rect 502334 695756 502340 695768
rect 492631 695728 492720 695756
rect 492631 695725 492643 695728
rect 492585 695719 492643 695725
rect 492692 695697 492720 695728
rect 502260 695728 502340 695756
rect 502260 695697 502288 695728
rect 502334 695716 502340 695728
rect 502392 695716 502398 695768
rect 578000 695728 582820 695824
rect 3752 695660 6132 695688
rect 17221 695691 17279 695697
rect 3752 695648 3758 695660
rect 17221 695657 17233 695691
rect 17267 695688 17279 695691
rect 31757 695691 31815 695697
rect 31757 695688 31769 695691
rect 17267 695660 31769 695688
rect 17267 695657 17279 695660
rect 17221 695651 17279 695657
rect 31757 695657 31769 695660
rect 31803 695657 31815 695691
rect 31757 695651 31815 695657
rect 55861 695691 55919 695697
rect 55861 695657 55873 695691
rect 55907 695688 55919 695691
rect 62761 695691 62819 695697
rect 62761 695688 62773 695691
rect 55907 695660 62773 695688
rect 55907 695657 55919 695660
rect 55861 695651 55919 695657
rect 62761 695657 62773 695660
rect 62807 695657 62819 695691
rect 62761 695651 62819 695657
rect 75181 695691 75239 695697
rect 75181 695657 75193 695691
rect 75227 695688 75239 695691
rect 82081 695691 82139 695697
rect 82081 695688 82093 695691
rect 75227 695660 82093 695688
rect 75227 695657 75239 695660
rect 75181 695651 75239 695657
rect 82081 695657 82093 695660
rect 82127 695657 82139 695691
rect 82081 695651 82139 695657
rect 94501 695691 94559 695697
rect 94501 695657 94513 695691
rect 94547 695688 94559 695691
rect 154577 695691 154635 695697
rect 154577 695688 154589 695691
rect 94547 695660 154589 695688
rect 94547 695657 94559 695660
rect 94501 695651 94559 695657
rect 154577 695657 154589 695660
rect 154623 695657 154635 695691
rect 154577 695651 154635 695657
rect 154853 695691 154911 695697
rect 154853 695657 154865 695691
rect 154899 695688 154911 695691
rect 173989 695691 174047 695697
rect 173989 695688 174001 695691
rect 154899 695660 174001 695688
rect 154899 695657 154911 695660
rect 154853 695651 154911 695657
rect 173989 695657 174001 695660
rect 174035 695657 174047 695691
rect 173989 695651 174047 695657
rect 174173 695691 174231 695697
rect 174173 695657 174185 695691
rect 174219 695688 174231 695691
rect 297269 695691 297327 695697
rect 297269 695688 297281 695691
rect 174219 695660 297281 695688
rect 174219 695657 174231 695660
rect 174173 695651 174231 695657
rect 297269 695657 297281 695660
rect 297315 695657 297327 695691
rect 297269 695651 297327 695657
rect 306929 695691 306987 695697
rect 306929 695657 306941 695691
rect 306975 695688 306987 695691
rect 355229 695691 355287 695697
rect 355229 695688 355241 695691
rect 306975 695660 355241 695688
rect 306975 695657 306987 695660
rect 306929 695651 306987 695657
rect 355229 695657 355241 695660
rect 355275 695657 355287 695691
rect 355229 695651 355287 695657
rect 362129 695691 362187 695697
rect 362129 695657 362141 695691
rect 362175 695688 362187 695691
rect 374641 695691 374699 695697
rect 374641 695688 374653 695691
rect 362175 695660 374653 695688
rect 362175 695657 362187 695660
rect 362129 695651 362187 695657
rect 374641 695657 374653 695660
rect 374687 695657 374699 695691
rect 374641 695651 374699 695657
rect 384301 695691 384359 695697
rect 384301 695657 384313 695691
rect 384347 695688 384359 695691
rect 393961 695691 394019 695697
rect 393961 695688 393973 695691
rect 384347 695660 393973 695688
rect 384347 695657 384359 695660
rect 384301 695651 384359 695657
rect 393961 695657 393973 695660
rect 394007 695657 394019 695691
rect 393961 695651 394019 695657
rect 403621 695691 403679 695697
rect 403621 695657 403633 695691
rect 403667 695688 403679 695691
rect 413281 695691 413339 695697
rect 413281 695688 413293 695691
rect 403667 695660 413293 695688
rect 403667 695657 403679 695660
rect 403621 695651 403679 695657
rect 413281 695657 413293 695660
rect 413327 695657 413339 695691
rect 413281 695651 413339 695657
rect 422941 695691 422999 695697
rect 422941 695657 422953 695691
rect 422987 695688 422999 695691
rect 432325 695691 432383 695697
rect 432325 695688 432337 695691
rect 422987 695660 432337 695688
rect 422987 695657 422999 695660
rect 422941 695651 422999 695657
rect 432325 695657 432337 695660
rect 432371 695657 432383 695691
rect 432325 695651 432383 695657
rect 442261 695691 442319 695697
rect 442261 695657 442273 695691
rect 442307 695688 442319 695691
rect 451277 695691 451335 695697
rect 451277 695688 451289 695691
rect 442307 695660 451289 695688
rect 442307 695657 442319 695660
rect 442261 695651 442319 695657
rect 451277 695657 451289 695660
rect 451323 695657 451335 695691
rect 451277 695651 451335 695657
rect 461397 695691 461455 695697
rect 461397 695657 461409 695691
rect 461443 695688 461455 695691
rect 471241 695691 471299 695697
rect 471241 695688 471253 695691
rect 461443 695660 471253 695688
rect 461443 695657 461455 695660
rect 461397 695651 461455 695657
rect 471241 695657 471253 695660
rect 471287 695657 471299 695691
rect 471241 695651 471299 695657
rect 492677 695691 492735 695697
rect 492677 695657 492689 695691
rect 492723 695657 492735 695691
rect 492677 695651 492735 695657
rect 502245 695691 502303 695697
rect 502245 695657 502257 695691
rect 502291 695657 502303 695691
rect 502245 695651 502303 695657
rect 7742 695580 7748 695632
rect 7800 695620 7806 695632
rect 173897 695623 173955 695629
rect 173897 695620 173909 695623
rect 7800 695592 154712 695620
rect 7800 695580 7806 695592
rect 4890 695512 4896 695564
rect 4948 695552 4954 695564
rect 17221 695555 17279 695561
rect 17221 695552 17233 695555
rect 4948 695524 17233 695552
rect 4948 695512 4954 695524
rect 17221 695521 17233 695524
rect 17267 695521 17279 695555
rect 17221 695515 17279 695521
rect 31757 695555 31815 695561
rect 31757 695521 31769 695555
rect 31803 695552 31815 695555
rect 46201 695555 46259 695561
rect 46201 695552 46213 695555
rect 31803 695524 46213 695552
rect 31803 695521 31815 695524
rect 31757 695515 31815 695521
rect 46201 695521 46213 695524
rect 46247 695521 46259 695555
rect 46201 695515 46259 695521
rect 53282 695512 53288 695564
rect 53340 695552 53346 695564
rect 154577 695555 154635 695561
rect 154577 695552 154589 695555
rect 53340 695524 154589 695552
rect 53340 695512 53346 695524
rect 154577 695521 154589 695524
rect 154623 695521 154635 695555
rect 154684 695552 154712 695592
rect 154776 695592 173909 695620
rect 154776 695552 154804 695592
rect 173897 695589 173909 695592
rect 173943 695589 173955 695623
rect 173897 695583 173955 695589
rect 174081 695623 174139 695629
rect 174081 695589 174093 695623
rect 174127 695620 174139 695623
rect 506934 695620 506940 695632
rect 174127 695592 506940 695620
rect 174127 695589 174139 695592
rect 174081 695583 174139 695589
rect 506934 695580 506940 695592
rect 506992 695580 506998 695632
rect 154684 695524 154804 695552
rect 154853 695555 154911 695561
rect 154577 695515 154635 695521
rect 154853 695521 154865 695555
rect 154899 695552 154911 695555
rect 173989 695555 174047 695561
rect 173989 695552 174001 695555
rect 154899 695524 174001 695552
rect 154899 695521 154911 695524
rect 154853 695515 154911 695521
rect 173989 695521 174001 695524
rect 174035 695521 174047 695555
rect 173989 695515 174047 695521
rect 174173 695555 174231 695561
rect 174173 695521 174185 695555
rect 174219 695552 174231 695555
rect 577498 695552 577504 695564
rect 174219 695524 577504 695552
rect 174219 695521 174231 695524
rect 174173 695515 174231 695521
rect 577498 695512 577504 695524
rect 577556 695512 577562 695564
rect 7190 695444 7196 695496
rect 7248 695484 7254 695496
rect 355502 695484 355508 695496
rect 7248 695456 355508 695484
rect 7248 695444 7254 695456
rect 355502 695444 355508 695456
rect 355560 695444 355566 695496
rect 355597 695487 355655 695493
rect 355597 695453 355609 695487
rect 355643 695484 355655 695487
rect 364981 695487 365039 695493
rect 364981 695484 364993 695487
rect 355643 695456 364993 695484
rect 355643 695453 355655 695456
rect 355597 695447 355655 695453
rect 364981 695453 364993 695456
rect 365027 695453 365039 695487
rect 364981 695447 365039 695453
rect 7282 695376 7288 695428
rect 7340 695416 7346 695428
rect 369946 695416 369952 695428
rect 7340 695388 369952 695416
rect 7340 695376 7346 695388
rect 369946 695376 369952 695388
rect 370004 695376 370010 695428
rect 374641 695419 374699 695425
rect 374641 695385 374653 695419
rect 374687 695416 374699 695419
rect 384301 695419 384359 695425
rect 384301 695416 384313 695419
rect 374687 695388 384313 695416
rect 374687 695385 374699 695388
rect 374641 695379 374699 695385
rect 384301 695385 384313 695388
rect 384347 695385 384359 695419
rect 384301 695379 384359 695385
rect 3234 695308 3240 695360
rect 3292 695348 3298 695360
rect 383838 695348 383844 695360
rect 3292 695320 383844 695348
rect 3292 695308 3298 695320
rect 383838 695308 383844 695320
rect 383896 695308 383902 695360
rect 393961 695351 394019 695357
rect 393961 695317 393973 695351
rect 394007 695348 394019 695351
rect 403621 695351 403679 695357
rect 403621 695348 403633 695351
rect 394007 695320 403633 695348
rect 394007 695317 394019 695320
rect 393961 695311 394019 695317
rect 403621 695317 403633 695320
rect 403667 695317 403679 695351
rect 403621 695311 403679 695317
rect 413281 695351 413339 695357
rect 413281 695317 413293 695351
rect 413327 695348 413339 695351
rect 422941 695351 422999 695357
rect 422941 695348 422953 695351
rect 413327 695320 422953 695348
rect 413327 695317 413339 695320
rect 413281 695311 413339 695317
rect 422941 695317 422953 695320
rect 422987 695317 422999 695351
rect 426526 695348 426532 695360
rect 426487 695320 426532 695348
rect 422941 695311 422999 695317
rect 426526 695308 426532 695320
rect 426584 695308 426590 695360
rect 440694 695348 440700 695360
rect 440655 695320 440700 695348
rect 440694 695308 440700 695320
rect 440752 695308 440758 695360
rect 469214 695348 469220 695360
rect 469175 695320 469220 695348
rect 469214 695308 469220 695320
rect 469272 695308 469278 695360
rect 497550 695348 497556 695360
rect 497511 695320 497556 695348
rect 497550 695308 497556 695320
rect 497608 695308 497614 695360
rect 511902 695348 511908 695360
rect 511863 695320 511908 695348
rect 511902 695308 511908 695320
rect 511960 695308 511966 695360
rect 578142 695348 578148 695360
rect 577516 695320 578148 695348
rect 57882 695280 57888 695292
rect 1104 695184 6000 695280
rect 57843 695252 57888 695280
rect 57882 695240 57888 695252
rect 57940 695240 57946 695292
rect 67450 695280 67456 695292
rect 67411 695252 67456 695280
rect 67450 695240 67456 695252
rect 67508 695240 67514 695292
rect 81342 695280 81348 695292
rect 81303 695252 81348 695280
rect 81342 695240 81348 695252
rect 81400 695240 81406 695292
rect 95786 695280 95792 695292
rect 95747 695252 95792 695280
rect 95786 695240 95792 695252
rect 95844 695240 95850 695292
rect 100570 695280 100576 695292
rect 100531 695252 100576 695280
rect 100570 695240 100576 695252
rect 100628 695240 100634 695292
rect 109954 695280 109960 695292
rect 109915 695252 109960 695280
rect 109954 695240 109960 695252
rect 110012 695240 110018 695292
rect 154577 695283 154635 695289
rect 154577 695280 154589 695283
rect 138032 695252 154589 695280
rect 57977 695215 58035 695221
rect 6104 695184 28948 695212
rect 4062 695036 4068 695088
rect 4120 695076 4126 695088
rect 6104 695076 6132 695184
rect 28920 695144 28948 695184
rect 33796 695184 45600 695212
rect 33796 695144 33824 695184
rect 28920 695116 33824 695144
rect 45572 695144 45600 695184
rect 57977 695181 57989 695215
rect 58023 695212 58035 695215
rect 75917 695215 75975 695221
rect 75917 695212 75929 695215
rect 58023 695184 75929 695212
rect 58023 695181 58035 695184
rect 57977 695175 58035 695181
rect 75917 695181 75929 695184
rect 75963 695181 75975 695215
rect 104897 695215 104955 695221
rect 104897 695212 104909 695215
rect 75917 695175 75975 695181
rect 104820 695184 104909 695212
rect 57793 695147 57851 695153
rect 57793 695144 57805 695147
rect 45572 695116 57805 695144
rect 57793 695113 57805 695116
rect 57839 695113 57851 695147
rect 104820 695144 104848 695184
rect 104897 695181 104909 695184
rect 104943 695181 104955 695215
rect 104897 695175 104955 695181
rect 117225 695215 117283 695221
rect 117225 695181 117237 695215
rect 117271 695212 117283 695215
rect 124309 695215 124367 695221
rect 124309 695212 124321 695215
rect 117271 695184 124321 695212
rect 117271 695181 117283 695184
rect 117225 695175 117283 695181
rect 124309 695181 124321 695184
rect 124355 695181 124367 695215
rect 124309 695175 124367 695181
rect 57793 695107 57851 695113
rect 79520 695116 104848 695144
rect 114465 695147 114523 695153
rect 4120 695048 6132 695076
rect 76009 695079 76067 695085
rect 4120 695036 4126 695048
rect 76009 695045 76021 695079
rect 76055 695076 76067 695079
rect 79520 695076 79548 695116
rect 114465 695113 114477 695147
rect 114511 695144 114523 695147
rect 114649 695147 114707 695153
rect 114649 695144 114661 695147
rect 114511 695116 114661 695144
rect 114511 695113 114523 695116
rect 114465 695107 114523 695113
rect 114649 695113 114661 695116
rect 114695 695113 114707 695147
rect 114649 695107 114707 695113
rect 124401 695147 124459 695153
rect 124401 695113 124413 695147
rect 124447 695144 124459 695147
rect 128265 695147 128323 695153
rect 128265 695144 128277 695147
rect 124447 695116 128277 695144
rect 124447 695113 124459 695116
rect 124401 695107 124459 695113
rect 128265 695113 128277 695116
rect 128311 695113 128323 695147
rect 128265 695107 128323 695113
rect 128357 695147 128415 695153
rect 128357 695113 128369 695147
rect 128403 695144 128415 695147
rect 138032 695144 138060 695252
rect 154577 695249 154589 695252
rect 154623 695249 154635 695283
rect 157426 695280 157432 695292
rect 157387 695252 157432 695280
rect 154577 695243 154635 695249
rect 157426 695240 157432 695252
rect 157484 695240 157490 695292
rect 166997 695283 167055 695289
rect 166997 695249 167009 695283
rect 167043 695280 167055 695283
rect 176565 695283 176623 695289
rect 176565 695280 176577 695283
rect 167043 695252 176577 695280
rect 167043 695249 167055 695252
rect 166997 695243 167055 695249
rect 176565 695249 176577 695252
rect 176611 695249 176623 695283
rect 176565 695243 176623 695249
rect 179322 695240 179328 695292
rect 179380 695240 179386 695292
rect 185762 695240 185768 695292
rect 185820 695240 185826 695292
rect 186317 695283 186375 695289
rect 186317 695249 186329 695283
rect 186363 695280 186375 695283
rect 195885 695283 195943 695289
rect 195885 695280 195897 695283
rect 186363 695252 195897 695280
rect 186363 695249 186375 695252
rect 186317 695243 186375 695249
rect 195885 695249 195897 695252
rect 195931 695249 195943 695283
rect 195885 695243 195943 695249
rect 199930 695240 199936 695292
rect 199988 695280 199994 695292
rect 577406 695280 577412 695292
rect 199988 695252 577412 695280
rect 199988 695240 199994 695252
rect 577406 695240 577412 695252
rect 577464 695240 577470 695292
rect 176473 695215 176531 695221
rect 176473 695181 176485 695215
rect 176519 695212 176531 695215
rect 179340 695212 179368 695240
rect 176519 695184 179368 695212
rect 185780 695212 185808 695240
rect 577516 695212 577544 695320
rect 578142 695308 578148 695320
rect 578200 695308 578206 695360
rect 185780 695184 577544 695212
rect 578000 695184 582820 695280
rect 176519 695181 176531 695184
rect 176473 695175 176531 695181
rect 128403 695116 138060 695144
rect 147677 695147 147735 695153
rect 128403 695113 128415 695116
rect 128357 695107 128415 695113
rect 147677 695113 147689 695147
rect 147723 695144 147735 695147
rect 156969 695147 157027 695153
rect 156969 695144 156981 695147
rect 147723 695116 156981 695144
rect 147723 695113 147735 695116
rect 147677 695107 147735 695113
rect 156969 695113 156981 695116
rect 157015 695113 157027 695147
rect 171505 695147 171563 695153
rect 171505 695144 171517 695147
rect 156969 695107 157027 695113
rect 157352 695116 171517 695144
rect 76055 695048 79548 695076
rect 154577 695079 154635 695085
rect 76055 695045 76067 695048
rect 76009 695039 76067 695045
rect 154577 695045 154589 695079
rect 154623 695076 154635 695079
rect 157352 695076 157380 695116
rect 171505 695113 171517 695116
rect 171551 695113 171563 695147
rect 171505 695107 171563 695113
rect 171597 695147 171655 695153
rect 171597 695113 171609 695147
rect 171643 695144 171655 695147
rect 578050 695144 578056 695156
rect 171643 695116 578056 695144
rect 171643 695113 171655 695116
rect 171597 695107 171655 695113
rect 578050 695104 578056 695116
rect 578108 695104 578114 695156
rect 154623 695048 157380 695076
rect 157429 695079 157487 695085
rect 154623 695045 154635 695048
rect 154577 695039 154635 695045
rect 157429 695045 157441 695079
rect 157475 695076 157487 695079
rect 576026 695076 576032 695088
rect 157475 695048 576032 695076
rect 157475 695045 157487 695048
rect 157429 695039 157487 695045
rect 576026 695036 576032 695048
rect 576084 695036 576090 695088
rect 7466 694968 7472 695020
rect 7524 695008 7530 695020
rect 426529 695011 426587 695017
rect 426529 695008 426541 695011
rect 7524 694980 426541 695008
rect 7524 694968 7530 694980
rect 426529 694977 426541 694980
rect 426575 694977 426587 695011
rect 426529 694971 426587 694977
rect 432601 695011 432659 695017
rect 432601 694977 432613 695011
rect 432647 695008 432659 695011
rect 441893 695011 441951 695017
rect 441893 695008 441905 695011
rect 432647 694980 441905 695008
rect 432647 694977 432659 694980
rect 432601 694971 432659 694977
rect 441893 694977 441905 694980
rect 441939 694977 441951 695011
rect 441893 694971 441951 694977
rect 3878 694900 3884 694952
rect 3936 694940 3942 694952
rect 95237 694943 95295 694949
rect 95237 694940 95249 694943
rect 3936 694912 95249 694940
rect 3936 694900 3942 694912
rect 95237 694909 95249 694912
rect 95283 694909 95295 694943
rect 95237 694903 95295 694909
rect 95421 694943 95479 694949
rect 95421 694909 95433 694943
rect 95467 694940 95479 694943
rect 440697 694943 440755 694949
rect 440697 694940 440709 694943
rect 95467 694912 440709 694940
rect 95467 694909 95479 694912
rect 95421 694903 95479 694909
rect 440697 694909 440709 694912
rect 440743 694909 440755 694943
rect 440697 694903 440755 694909
rect 451277 694943 451335 694949
rect 451277 694909 451289 694943
rect 451323 694940 451335 694943
rect 461581 694943 461639 694949
rect 461581 694940 461593 694943
rect 451323 694912 461593 694940
rect 451323 694909 451335 694912
rect 451277 694903 451335 694909
rect 461581 694909 461593 694912
rect 461627 694909 461639 694943
rect 461581 694903 461639 694909
rect 19245 694875 19303 694881
rect 19245 694841 19257 694875
rect 19291 694872 19303 694875
rect 28813 694875 28871 694881
rect 28813 694872 28825 694875
rect 19291 694844 28825 694872
rect 19291 694841 19303 694844
rect 19245 694835 19303 694841
rect 28813 694841 28825 694844
rect 28859 694841 28871 694875
rect 28813 694835 28871 694841
rect 86957 694875 87015 694881
rect 86957 694841 86969 694875
rect 87003 694872 87015 694875
rect 97997 694875 98055 694881
rect 97997 694872 98009 694875
rect 87003 694844 98009 694872
rect 87003 694841 87015 694844
rect 86957 694835 87015 694841
rect 97997 694841 98009 694844
rect 98043 694841 98055 694875
rect 97997 694835 98055 694841
rect 104897 694875 104955 694881
rect 104897 694841 104909 694875
rect 104943 694872 104955 694875
rect 114465 694875 114523 694881
rect 114465 694872 114477 694875
rect 104943 694844 114477 694872
rect 104943 694841 104955 694844
rect 104897 694835 104955 694841
rect 114465 694841 114477 694844
rect 114511 694841 114523 694875
rect 114465 694835 114523 694841
rect 114649 694875 114707 694881
rect 114649 694841 114661 694875
rect 114695 694872 114707 694875
rect 117225 694875 117283 694881
rect 117225 694872 117237 694875
rect 114695 694844 117237 694872
rect 114695 694841 114707 694844
rect 114649 694835 114707 694841
rect 117225 694841 117237 694844
rect 117271 694841 117283 694875
rect 117225 694835 117283 694841
rect 124125 694875 124183 694881
rect 124125 694841 124137 694875
rect 124171 694872 124183 694875
rect 125321 694875 125379 694881
rect 125321 694872 125333 694875
rect 124171 694844 125333 694872
rect 124171 694841 124183 694844
rect 124125 694835 124183 694841
rect 125321 694841 125333 694844
rect 125367 694841 125379 694875
rect 125321 694835 125379 694841
rect 125597 694875 125655 694881
rect 125597 694841 125609 694875
rect 125643 694841 125655 694875
rect 125597 694835 125655 694841
rect 125873 694875 125931 694881
rect 125873 694841 125885 694875
rect 125919 694872 125931 694875
rect 137281 694875 137339 694881
rect 137281 694872 137293 694875
rect 125919 694844 137293 694872
rect 125919 694841 125931 694844
rect 125873 694835 125931 694841
rect 137281 694841 137293 694844
rect 137327 694841 137339 694875
rect 137281 694835 137339 694841
rect 138477 694875 138535 694881
rect 138477 694841 138489 694875
rect 138523 694872 138535 694875
rect 576670 694872 576676 694884
rect 138523 694844 576676 694872
rect 138523 694841 138535 694844
rect 138477 694835 138535 694841
rect 3786 694764 3792 694816
rect 3844 694804 3850 694816
rect 9677 694807 9735 694813
rect 9677 694804 9689 694807
rect 3844 694776 9689 694804
rect 3844 694764 3850 694776
rect 9677 694773 9689 694776
rect 9723 694773 9735 694807
rect 9677 694767 9735 694773
rect 28905 694807 28963 694813
rect 28905 694773 28917 694807
rect 28951 694804 28963 694807
rect 44177 694807 44235 694813
rect 44177 694804 44189 694807
rect 28951 694776 33824 694804
rect 28951 694773 28963 694776
rect 28905 694767 28963 694773
rect 33796 694736 33824 694776
rect 41156 694776 44189 694804
rect 41156 694736 41184 694776
rect 44177 694773 44189 694776
rect 44223 694773 44235 694807
rect 75917 694807 75975 694813
rect 75917 694804 75929 694807
rect 44177 694767 44235 694773
rect 67560 694776 75929 694804
rect 1104 694640 6000 694736
rect 33796 694708 41184 694736
rect 53745 694739 53803 694745
rect 53745 694705 53757 694739
rect 53791 694736 53803 694739
rect 67560 694736 67588 694776
rect 75917 694773 75929 694776
rect 75963 694773 75975 694807
rect 75917 694767 75975 694773
rect 98089 694807 98147 694813
rect 98089 694773 98101 694807
rect 98135 694804 98147 694807
rect 106277 694807 106335 694813
rect 106277 694804 106289 694807
rect 98135 694776 106289 694804
rect 98135 694773 98147 694776
rect 98089 694767 98147 694773
rect 106277 694773 106289 694776
rect 106323 694773 106335 694807
rect 106277 694767 106335 694773
rect 106369 694807 106427 694813
rect 106369 694773 106381 694807
rect 106415 694804 106427 694807
rect 110233 694807 110291 694813
rect 110233 694804 110245 694807
rect 106415 694776 110245 694804
rect 106415 694773 106427 694776
rect 106369 694767 106427 694773
rect 110233 694773 110245 694776
rect 110279 694773 110291 694807
rect 110233 694767 110291 694773
rect 110325 694807 110383 694813
rect 110325 694773 110337 694807
rect 110371 694804 110383 694807
rect 114557 694807 114615 694813
rect 114557 694804 114569 694807
rect 110371 694776 114569 694804
rect 110371 694773 110383 694776
rect 110325 694767 110383 694773
rect 114557 694773 114569 694776
rect 114603 694773 114615 694807
rect 114557 694767 114615 694773
rect 125505 694807 125563 694813
rect 125505 694773 125517 694807
rect 125551 694804 125563 694807
rect 125612 694804 125640 694835
rect 576670 694832 576676 694844
rect 576728 694832 576734 694884
rect 125551 694776 125640 694804
rect 125781 694807 125839 694813
rect 125551 694773 125563 694776
rect 125505 694767 125563 694773
rect 125781 694773 125793 694807
rect 125827 694804 125839 694807
rect 138201 694807 138259 694813
rect 138201 694804 138213 694807
rect 125827 694776 138213 694804
rect 125827 694773 125839 694776
rect 125781 694767 125839 694773
rect 138201 694773 138213 694776
rect 138247 694773 138259 694807
rect 138201 694767 138259 694773
rect 138385 694807 138443 694813
rect 138385 694773 138397 694807
rect 138431 694804 138443 694807
rect 579062 694804 579068 694816
rect 138431 694776 579068 694804
rect 138431 694773 138443 694776
rect 138385 694767 138443 694773
rect 579062 694764 579068 694776
rect 579120 694764 579126 694816
rect 86865 694739 86923 694745
rect 86865 694736 86877 694739
rect 53791 694708 57836 694736
rect 53791 694705 53803 694708
rect 53745 694699 53803 694705
rect 9677 694671 9735 694677
rect 9677 694637 9689 694671
rect 9723 694668 9735 694671
rect 19245 694671 19303 694677
rect 19245 694668 19257 694671
rect 9723 694640 19257 694668
rect 9723 694637 9735 694640
rect 9677 694631 9735 694637
rect 19245 694637 19257 694640
rect 19291 694637 19303 694671
rect 57808 694668 57836 694708
rect 57992 694708 67588 694736
rect 85500 694708 86877 694736
rect 57992 694668 58020 694708
rect 57808 694640 58020 694668
rect 75917 694671 75975 694677
rect 19245 694631 19303 694637
rect 75917 694637 75929 694671
rect 75963 694668 75975 694671
rect 85500 694668 85528 694708
rect 86865 694705 86877 694708
rect 86911 694705 86923 694739
rect 86865 694699 86923 694705
rect 124125 694739 124183 694745
rect 124125 694705 124137 694739
rect 124171 694736 124183 694739
rect 125689 694739 125747 694745
rect 125689 694736 125701 694739
rect 124171 694708 125701 694736
rect 124171 694705 124183 694708
rect 124125 694699 124183 694705
rect 125689 694705 125701 694708
rect 125735 694705 125747 694739
rect 125689 694699 125747 694705
rect 137281 694739 137339 694745
rect 137281 694705 137293 694739
rect 137327 694736 137339 694739
rect 147677 694739 147735 694745
rect 147677 694736 147689 694739
rect 137327 694708 147689 694736
rect 137327 694705 137339 694708
rect 137281 694699 137339 694705
rect 147677 694705 147689 694708
rect 147723 694705 147735 694739
rect 147677 694699 147735 694705
rect 156969 694739 157027 694745
rect 156969 694705 156981 694739
rect 157015 694736 157027 694739
rect 166997 694739 167055 694745
rect 166997 694736 167009 694739
rect 157015 694708 167009 694736
rect 157015 694705 157027 694708
rect 156969 694699 157027 694705
rect 166997 694705 167009 694708
rect 167043 694705 167055 694739
rect 166997 694699 167055 694705
rect 176565 694739 176623 694745
rect 176565 694705 176577 694739
rect 176611 694736 176623 694739
rect 186317 694739 186375 694745
rect 186317 694736 186329 694739
rect 176611 694708 186329 694736
rect 176611 694705 176623 694708
rect 176565 694699 176623 694705
rect 186317 694705 186329 694708
rect 186363 694705 186375 694739
rect 186317 694699 186375 694705
rect 195885 694739 195943 694745
rect 195885 694705 195897 694739
rect 195931 694736 195943 694739
rect 205637 694739 205695 694745
rect 205637 694736 205649 694739
rect 195931 694708 205649 694736
rect 195931 694705 195943 694708
rect 195885 694699 195943 694705
rect 205637 694705 205649 694708
rect 205683 694705 205695 694739
rect 205637 694699 205695 694705
rect 215205 694739 215263 694745
rect 215205 694705 215217 694739
rect 215251 694736 215263 694739
rect 224957 694739 225015 694745
rect 224957 694736 224969 694739
rect 215251 694708 224969 694736
rect 215251 694705 215263 694708
rect 215205 694699 215263 694705
rect 224957 694705 224969 694708
rect 225003 694705 225015 694739
rect 224957 694699 225015 694705
rect 234525 694739 234583 694745
rect 234525 694705 234537 694739
rect 234571 694736 234583 694739
rect 244277 694739 244335 694745
rect 244277 694736 244289 694739
rect 234571 694708 244289 694736
rect 234571 694705 234583 694708
rect 234525 694699 234583 694705
rect 244277 694705 244289 694708
rect 244323 694705 244335 694739
rect 244277 694699 244335 694705
rect 253845 694739 253903 694745
rect 253845 694705 253857 694739
rect 253891 694736 253903 694739
rect 263597 694739 263655 694745
rect 263597 694736 263609 694739
rect 253891 694708 263609 694736
rect 253891 694705 253903 694708
rect 253845 694699 253903 694705
rect 263597 694705 263609 694708
rect 263643 694705 263655 694739
rect 263597 694699 263655 694705
rect 273165 694739 273223 694745
rect 273165 694705 273177 694739
rect 273211 694736 273223 694739
rect 282917 694739 282975 694745
rect 282917 694736 282929 694739
rect 273211 694708 282929 694736
rect 273211 694705 273223 694708
rect 273165 694699 273223 694705
rect 282917 694705 282929 694708
rect 282963 694705 282975 694739
rect 282917 694699 282975 694705
rect 292485 694739 292543 694745
rect 292485 694705 292497 694739
rect 292531 694736 292543 694739
rect 302145 694739 302203 694745
rect 302145 694736 302157 694739
rect 292531 694708 302157 694736
rect 292531 694705 292543 694708
rect 292485 694699 292543 694705
rect 302145 694705 302157 694708
rect 302191 694705 302203 694739
rect 302145 694699 302203 694705
rect 302237 694739 302295 694745
rect 302237 694705 302249 694739
rect 302283 694736 302295 694739
rect 355597 694739 355655 694745
rect 355597 694736 355609 694739
rect 302283 694708 355609 694736
rect 302283 694705 302295 694708
rect 302237 694699 302295 694705
rect 355597 694705 355609 694708
rect 355643 694705 355655 694739
rect 355597 694699 355655 694705
rect 364981 694739 365039 694745
rect 364981 694705 364993 694739
rect 365027 694736 365039 694739
rect 374641 694739 374699 694745
rect 374641 694736 374653 694739
rect 365027 694708 374653 694736
rect 365027 694705 365039 694708
rect 364981 694699 365039 694705
rect 374641 694705 374653 694708
rect 374687 694705 374699 694739
rect 374641 694699 374699 694705
rect 384301 694739 384359 694745
rect 384301 694705 384313 694739
rect 384347 694736 384359 694739
rect 393961 694739 394019 694745
rect 393961 694736 393973 694739
rect 384347 694708 393973 694736
rect 384347 694705 384359 694708
rect 384301 694699 384359 694705
rect 393961 694705 393973 694708
rect 394007 694705 394019 694739
rect 393961 694699 394019 694705
rect 403621 694739 403679 694745
rect 403621 694705 403633 694739
rect 403667 694736 403679 694739
rect 413281 694739 413339 694745
rect 413281 694736 413293 694739
rect 403667 694708 413293 694736
rect 403667 694705 403679 694708
rect 403621 694699 403679 694705
rect 413281 694705 413293 694708
rect 413327 694705 413339 694739
rect 413281 694699 413339 694705
rect 422941 694739 422999 694745
rect 422941 694705 422953 694739
rect 422987 694736 422999 694739
rect 432601 694739 432659 694745
rect 432601 694736 432613 694739
rect 422987 694708 432613 694736
rect 422987 694705 422999 694708
rect 422941 694699 422999 694705
rect 432601 694705 432613 694708
rect 432647 694705 432659 694739
rect 432601 694699 432659 694705
rect 441893 694739 441951 694745
rect 441893 694705 441905 694739
rect 441939 694736 441951 694739
rect 451277 694739 451335 694745
rect 451277 694736 451289 694739
rect 441939 694708 451289 694736
rect 441939 694705 441951 694708
rect 441893 694699 441951 694705
rect 451277 694705 451289 694708
rect 451323 694705 451335 694739
rect 451277 694699 451335 694705
rect 461581 694739 461639 694745
rect 461581 694705 461593 694739
rect 461627 694736 461639 694739
rect 469217 694739 469275 694745
rect 469217 694736 469229 694739
rect 461627 694708 469229 694736
rect 461627 694705 461639 694708
rect 461581 694699 461639 694705
rect 469217 694705 469229 694708
rect 469263 694705 469275 694739
rect 469217 694699 469275 694705
rect 75963 694640 85528 694668
rect 109957 694671 110015 694677
rect 75963 694637 75975 694640
rect 75917 694631 75975 694637
rect 109957 694637 109969 694671
rect 110003 694668 110015 694671
rect 576486 694668 576492 694680
rect 110003 694640 576492 694668
rect 110003 694637 110015 694640
rect 109957 694631 110015 694637
rect 576486 694628 576492 694640
rect 576544 694628 576550 694680
rect 578000 694640 582820 694736
rect 44177 694603 44235 694609
rect 44177 694569 44189 694603
rect 44223 694600 44235 694603
rect 53745 694603 53803 694609
rect 53745 694600 53757 694603
rect 44223 694572 53757 694600
rect 44223 694569 44235 694572
rect 44177 694563 44235 694569
rect 53745 694569 53757 694572
rect 53791 694569 53803 694603
rect 53745 694563 53803 694569
rect 100573 694603 100631 694609
rect 100573 694569 100585 694603
rect 100619 694600 100631 694603
rect 578970 694600 578976 694612
rect 100619 694572 578976 694600
rect 100619 694569 100631 694572
rect 100573 694563 100631 694569
rect 578970 694560 578976 694572
rect 579028 694560 579034 694612
rect 95789 694535 95847 694541
rect 95789 694501 95801 694535
rect 95835 694532 95847 694535
rect 125597 694535 125655 694541
rect 125597 694532 125609 694535
rect 95835 694504 125609 694532
rect 95835 694501 95847 694504
rect 95789 694495 95847 694501
rect 125597 694501 125609 694504
rect 125643 694501 125655 694535
rect 125597 694495 125655 694501
rect 125873 694535 125931 694541
rect 125873 694501 125885 694535
rect 125919 694532 125931 694535
rect 575290 694532 575296 694544
rect 125919 694504 575296 694532
rect 125919 694501 125931 694504
rect 125873 694495 125931 694501
rect 575290 694492 575296 694504
rect 575348 694492 575354 694544
rect 7834 694424 7840 694476
rect 7892 694464 7898 694476
rect 497553 694467 497611 694473
rect 497553 694464 497565 694467
rect 7892 694436 497565 694464
rect 7892 694424 7898 694436
rect 497553 694433 497565 694436
rect 497599 694433 497611 694467
rect 497553 694427 497611 694433
rect 81345 694399 81403 694405
rect 81345 694365 81357 694399
rect 81391 694396 81403 694399
rect 125689 694399 125747 694405
rect 125689 694396 125701 694399
rect 81391 694368 125701 694396
rect 81391 694365 81403 694368
rect 81345 694359 81403 694365
rect 125689 694365 125701 694368
rect 125735 694365 125747 694399
rect 125689 694359 125747 694365
rect 125781 694399 125839 694405
rect 125781 694365 125793 694399
rect 125827 694396 125839 694399
rect 575198 694396 575204 694408
rect 125827 694368 575204 694396
rect 125827 694365 125839 694368
rect 125781 694359 125839 694365
rect 575198 694356 575204 694368
rect 575256 694356 575262 694408
rect 67453 694331 67511 694337
rect 67453 694297 67465 694331
rect 67499 694328 67511 694331
rect 125597 694331 125655 694337
rect 125597 694328 125609 694331
rect 67499 694300 125609 694328
rect 67499 694297 67511 694300
rect 67453 694291 67511 694297
rect 125597 694297 125609 694300
rect 125643 694297 125655 694331
rect 125597 694291 125655 694297
rect 125873 694331 125931 694337
rect 125873 694297 125885 694331
rect 125919 694328 125931 694331
rect 575106 694328 575112 694340
rect 125919 694300 575112 694328
rect 125919 694297 125931 694300
rect 125873 694291 125931 694297
rect 575106 694288 575112 694300
rect 575164 694288 575170 694340
rect 3602 694220 3608 694272
rect 3660 694260 3666 694272
rect 511905 694263 511963 694269
rect 511905 694260 511917 694263
rect 3660 694232 511917 694260
rect 3660 694220 3666 694232
rect 511905 694229 511917 694232
rect 511951 694229 511963 694263
rect 511905 694223 511963 694229
rect 57885 694195 57943 694201
rect 1104 694096 6000 694192
rect 57885 694161 57897 694195
rect 57931 694192 57943 694195
rect 575014 694192 575020 694204
rect 57931 694164 575020 694192
rect 57931 694161 57943 694164
rect 57885 694155 57943 694161
rect 575014 694152 575020 694164
rect 575072 694152 575078 694204
rect 171505 694127 171563 694133
rect 171505 694093 171517 694127
rect 171551 694124 171563 694127
rect 176473 694127 176531 694133
rect 176473 694124 176485 694127
rect 171551 694096 176485 694124
rect 171551 694093 171563 694096
rect 171505 694087 171563 694093
rect 176473 694093 176485 694096
rect 176519 694093 176531 694127
rect 176473 694087 176531 694093
rect 205637 694127 205695 694133
rect 205637 694093 205649 694127
rect 205683 694124 205695 694127
rect 215205 694127 215263 694133
rect 215205 694124 215217 694127
rect 205683 694096 215217 694124
rect 205683 694093 205695 694096
rect 205637 694087 205695 694093
rect 215205 694093 215217 694096
rect 215251 694093 215263 694127
rect 215205 694087 215263 694093
rect 224957 694127 225015 694133
rect 224957 694093 224969 694127
rect 225003 694124 225015 694127
rect 234525 694127 234583 694133
rect 234525 694124 234537 694127
rect 225003 694096 234537 694124
rect 225003 694093 225015 694096
rect 224957 694087 225015 694093
rect 234525 694093 234537 694096
rect 234571 694093 234583 694127
rect 234525 694087 234583 694093
rect 244277 694127 244335 694133
rect 244277 694093 244289 694127
rect 244323 694124 244335 694127
rect 253845 694127 253903 694133
rect 253845 694124 253857 694127
rect 244323 694096 253857 694124
rect 244323 694093 244335 694096
rect 244277 694087 244335 694093
rect 253845 694093 253857 694096
rect 253891 694093 253903 694127
rect 253845 694087 253903 694093
rect 263597 694127 263655 694133
rect 263597 694093 263609 694127
rect 263643 694124 263655 694127
rect 273165 694127 273223 694133
rect 273165 694124 273177 694127
rect 263643 694096 273177 694124
rect 263643 694093 263655 694096
rect 263597 694087 263655 694093
rect 273165 694093 273177 694096
rect 273211 694093 273223 694127
rect 273165 694087 273223 694093
rect 282917 694127 282975 694133
rect 282917 694093 282929 694127
rect 282963 694124 282975 694127
rect 292485 694127 292543 694133
rect 292485 694124 292497 694127
rect 282963 694096 292497 694124
rect 282963 694093 282975 694096
rect 282917 694087 282975 694093
rect 292485 694093 292497 694096
rect 292531 694093 292543 694127
rect 292485 694087 292543 694093
rect 302145 694127 302203 694133
rect 302145 694093 302157 694127
rect 302191 694124 302203 694127
rect 302237 694127 302295 694133
rect 302237 694124 302249 694127
rect 302191 694096 302249 694124
rect 302191 694093 302203 694096
rect 302145 694087 302203 694093
rect 302237 694093 302249 694096
rect 302283 694093 302295 694127
rect 578000 694096 582820 694192
rect 302237 694087 302295 694093
rect 1104 693552 6000 693648
rect 578000 693552 582820 693648
rect 3142 693336 3148 693388
rect 3200 693376 3206 693388
rect 6089 693379 6147 693385
rect 6089 693376 6101 693379
rect 3200 693348 6101 693376
rect 3200 693336 3206 693348
rect 6089 693345 6101 693348
rect 6135 693345 6147 693379
rect 6089 693339 6147 693345
rect 1104 693008 6000 693104
rect 578000 693008 582820 693104
rect 1104 692464 6000 692560
rect 578000 692464 582820 692560
rect 1104 691920 6000 692016
rect 578000 691920 582820 692016
rect 1104 691376 6000 691472
rect 578000 691376 582820 691472
rect 1104 690832 6000 690928
rect 578000 690832 582820 690928
rect 1104 690288 6000 690384
rect 578000 690288 582820 690384
rect 1104 689744 6000 689840
rect 578000 689744 582820 689840
rect 1104 689200 6000 689296
rect 578000 689200 582820 689296
rect 1104 688656 6000 688752
rect 578000 688656 582820 688752
rect 1104 688112 6000 688208
rect 578000 688112 582820 688208
rect 1104 687568 6000 687664
rect 578000 687568 582820 687664
rect 578786 687148 578792 687200
rect 578844 687188 578850 687200
rect 580902 687188 580908 687200
rect 578844 687160 580908 687188
rect 578844 687148 578850 687160
rect 580902 687148 580908 687160
rect 580960 687148 580966 687200
rect 1104 687024 6000 687120
rect 578000 687024 582820 687120
rect 1104 686480 6000 686576
rect 578000 686480 582820 686576
rect 1104 685936 6000 686032
rect 578000 685936 582820 686032
rect 1104 685392 6000 685488
rect 578000 685392 582820 685488
rect 1104 684848 6000 684944
rect 578000 684848 582820 684944
rect 1104 684304 6000 684400
rect 578000 684304 582820 684400
rect 1104 683760 6000 683856
rect 578000 683760 582820 683856
rect 1104 683216 6000 683312
rect 578000 683216 582820 683312
rect 1104 682672 6000 682768
rect 578000 682672 582820 682768
rect 2866 682320 2872 682372
rect 2924 682360 2930 682372
rect 5718 682360 5724 682372
rect 2924 682332 5724 682360
rect 2924 682320 2930 682332
rect 5718 682320 5724 682332
rect 5776 682320 5782 682372
rect 1104 682128 6000 682224
rect 578000 682128 582820 682224
rect 1104 681584 6000 681680
rect 578000 681584 582820 681680
rect 1104 681040 6000 681136
rect 578000 681040 582820 681136
rect 1104 680496 6000 680592
rect 578000 680496 582820 680592
rect 1104 679952 6000 680048
rect 578000 679952 582820 680048
rect 1104 679408 6000 679504
rect 578000 679408 582820 679504
rect 1104 678864 6000 678960
rect 578000 678864 582820 678960
rect 1104 678320 6000 678416
rect 578000 678320 582820 678416
rect 1104 677776 6000 677872
rect 578000 677776 582820 677872
rect 1104 677232 6000 677328
rect 578000 677232 582820 677328
rect 1104 676688 6000 676784
rect 578000 676688 582820 676784
rect 1104 676144 6000 676240
rect 578000 676144 582820 676240
rect 1104 675600 6000 675696
rect 578000 675600 582820 675696
rect 1104 675056 6000 675152
rect 578000 675056 582820 675152
rect 575474 674772 575480 674824
rect 575532 674812 575538 674824
rect 579798 674812 579804 674824
rect 575532 674784 579804 674812
rect 575532 674772 575538 674784
rect 579798 674772 579804 674784
rect 579856 674772 579862 674824
rect 1104 674512 6000 674608
rect 578000 674512 582820 674608
rect 1104 673968 6000 674064
rect 578000 673968 582820 674064
rect 1104 673424 6000 673520
rect 578000 673424 582820 673520
rect 1104 672880 6000 672976
rect 578000 672880 582820 672976
rect 1104 672336 6000 672432
rect 578000 672336 582820 672432
rect 1104 671792 6000 671888
rect 578000 671792 582820 671888
rect 1104 671248 6000 671344
rect 578000 671248 582820 671344
rect 1104 670704 6000 670800
rect 578000 670704 582820 670800
rect 1104 670160 6000 670256
rect 578000 670160 582820 670256
rect 1104 669616 6000 669712
rect 578000 669616 582820 669712
rect 1104 669072 6000 669168
rect 578000 669072 582820 669168
rect 1104 668528 6000 668624
rect 578000 668528 582820 668624
rect 2774 668108 2780 668160
rect 2832 668148 2838 668160
rect 4706 668148 4712 668160
rect 2832 668120 4712 668148
rect 2832 668108 2838 668120
rect 4706 668108 4712 668120
rect 4764 668108 4770 668160
rect 1104 667984 6000 668080
rect 578000 667984 582820 668080
rect 1104 667440 6000 667536
rect 578000 667440 582820 667536
rect 1104 666896 6000 666992
rect 578000 666896 582820 666992
rect 1104 666352 6000 666448
rect 578000 666352 582820 666448
rect 1104 665808 6000 665904
rect 578000 665808 582820 665904
rect 1104 665264 6000 665360
rect 578000 665264 582820 665360
rect 1104 664720 6000 664816
rect 578000 664720 582820 664816
rect 1104 664176 6000 664272
rect 578000 664176 582820 664272
rect 1104 663632 6000 663728
rect 578000 663632 582820 663728
rect 1104 663088 6000 663184
rect 578000 663088 582820 663184
rect 1104 662544 6000 662640
rect 578000 662544 582820 662640
rect 1104 662000 6000 662096
rect 578000 662000 582820 662096
rect 1104 661456 6000 661552
rect 578000 661456 582820 661552
rect 1104 660912 6000 661008
rect 578000 660912 582820 661008
rect 1104 660368 6000 660464
rect 578000 660368 582820 660464
rect 1104 659824 6000 659920
rect 578000 659824 582820 659920
rect 1104 659280 6000 659376
rect 578000 659280 582820 659376
rect 1104 658736 6000 658832
rect 578000 658736 582820 658832
rect 1104 658192 6000 658288
rect 578000 658192 582820 658288
rect 1104 657648 6000 657744
rect 578000 657648 582820 657744
rect 1104 657104 6000 657200
rect 578000 657104 582820 657200
rect 1104 656560 6000 656656
rect 578000 656560 582820 656656
rect 1104 656016 6000 656112
rect 578000 656016 582820 656112
rect 1104 655472 6000 655568
rect 578000 655472 582820 655568
rect 1104 654928 6000 655024
rect 578000 654928 582820 655024
rect 1104 654384 6000 654480
rect 578000 654384 582820 654480
rect 1104 653840 6000 653936
rect 578000 653840 582820 653936
rect 3050 653556 3056 653608
rect 3108 653596 3114 653608
rect 7190 653596 7196 653608
rect 3108 653568 7196 653596
rect 3108 653556 3114 653568
rect 7190 653556 7196 653568
rect 7248 653556 7254 653608
rect 1104 653296 6000 653392
rect 578000 653296 582820 653392
rect 1104 652752 6000 652848
rect 578000 652752 582820 652848
rect 1104 652208 6000 652304
rect 578000 652208 582820 652304
rect 1104 651664 6000 651760
rect 578000 651664 582820 651760
rect 577406 651312 577412 651364
rect 577464 651352 577470 651364
rect 579614 651352 579620 651364
rect 577464 651324 579620 651352
rect 577464 651312 577470 651324
rect 579614 651312 579620 651324
rect 579672 651312 579678 651364
rect 1104 651120 6000 651216
rect 578000 651120 582820 651216
rect 1104 650576 6000 650672
rect 578000 650576 582820 650672
rect 1104 650032 6000 650128
rect 578000 650032 582820 650128
rect 1104 649488 6000 649584
rect 578000 649488 582820 649584
rect 1104 648944 6000 649040
rect 578000 648944 582820 649040
rect 1104 648400 6000 648496
rect 578000 648400 582820 648496
rect 1104 647856 6000 647952
rect 578000 647856 582820 647952
rect 1104 647312 6000 647408
rect 578000 647312 582820 647408
rect 1104 646768 6000 646864
rect 578000 646768 582820 646864
rect 1104 646224 6000 646320
rect 578000 646224 582820 646320
rect 1104 645680 6000 645776
rect 578000 645680 582820 645776
rect 1104 645136 6000 645232
rect 578000 645136 582820 645232
rect 1104 644592 6000 644688
rect 578000 644592 582820 644688
rect 1104 644048 6000 644144
rect 578000 644048 582820 644144
rect 1104 643504 6000 643600
rect 578000 643504 582820 643600
rect 1104 642960 6000 643056
rect 578000 642960 582820 643056
rect 1104 642416 6000 642512
rect 578000 642416 582820 642512
rect 1104 641872 6000 641968
rect 578000 641872 582820 641968
rect 1104 641328 6000 641424
rect 578000 641328 582820 641424
rect 1104 640784 6000 640880
rect 578000 640784 582820 640880
rect 1104 640240 6000 640336
rect 578000 640240 582820 640336
rect 1104 639696 6000 639792
rect 578000 639696 582820 639792
rect 1104 639152 6000 639248
rect 578000 639152 582820 639248
rect 1104 638608 6000 638704
rect 578000 638608 582820 638704
rect 1104 638064 6000 638160
rect 578000 638064 582820 638160
rect 1104 637520 6000 637616
rect 578000 637520 582820 637616
rect 1104 636976 6000 637072
rect 578000 636976 582820 637072
rect 1104 636432 6000 636528
rect 578000 636432 582820 636528
rect 1104 635888 6000 635984
rect 578000 635888 582820 635984
rect 1104 635344 6000 635440
rect 578000 635344 582820 635440
rect 1104 634800 6000 634896
rect 578000 634800 582820 634896
rect 1104 634256 6000 634352
rect 578000 634256 582820 634352
rect 1104 633712 6000 633808
rect 578000 633712 582820 633808
rect 1104 633168 6000 633264
rect 578000 633168 582820 633264
rect 1104 632624 6000 632720
rect 578000 632624 582820 632720
rect 1104 632080 6000 632176
rect 578000 632080 582820 632176
rect 1104 631536 6000 631632
rect 578000 631536 582820 631632
rect 1104 630992 6000 631088
rect 578000 630992 582820 631088
rect 1104 630448 6000 630544
rect 578000 630448 582820 630544
rect 1104 629904 6000 630000
rect 578000 629904 582820 630000
rect 1104 629360 6000 629456
rect 578000 629360 582820 629456
rect 1104 628816 6000 628912
rect 578000 628816 582820 628912
rect 1104 628272 6000 628368
rect 578000 628272 582820 628368
rect 575474 627852 575480 627904
rect 575532 627892 575538 627904
rect 579798 627892 579804 627904
rect 575532 627864 579804 627892
rect 575532 627852 575538 627864
rect 579798 627852 579804 627864
rect 579856 627852 579862 627904
rect 1104 627728 6000 627824
rect 578000 627728 582820 627824
rect 1104 627184 6000 627280
rect 578000 627184 582820 627280
rect 1104 626640 6000 626736
rect 578000 626640 582820 626736
rect 1104 626096 6000 626192
rect 578000 626096 582820 626192
rect 1104 625552 6000 625648
rect 578000 625552 582820 625648
rect 1104 625008 6000 625104
rect 578000 625008 582820 625104
rect 2958 624860 2964 624912
rect 3016 624900 3022 624912
rect 5810 624900 5816 624912
rect 3016 624872 5816 624900
rect 3016 624860 3022 624872
rect 5810 624860 5816 624872
rect 5868 624860 5874 624912
rect 1104 624464 6000 624560
rect 578000 624464 582820 624560
rect 1104 623920 6000 624016
rect 578000 623920 582820 624016
rect 1104 623376 6000 623472
rect 578000 623376 582820 623472
rect 1104 622832 6000 622928
rect 578000 622832 582820 622928
rect 1104 622288 6000 622384
rect 578000 622288 582820 622384
rect 1104 621744 6000 621840
rect 578000 621744 582820 621840
rect 1104 621200 6000 621296
rect 578000 621200 582820 621296
rect 1104 620656 6000 620752
rect 578000 620656 582820 620752
rect 1104 620112 6000 620208
rect 578000 620112 582820 620208
rect 1104 619568 6000 619664
rect 578000 619568 582820 619664
rect 1104 619024 6000 619120
rect 578000 619024 582820 619120
rect 1104 618480 6000 618576
rect 578000 618480 582820 618576
rect 1104 617936 6000 618032
rect 578000 617936 582820 618032
rect 1104 617392 6000 617488
rect 578000 617392 582820 617488
rect 1104 616848 6000 616944
rect 578000 616848 582820 616944
rect 1104 616304 6000 616400
rect 578000 616304 582820 616400
rect 1104 615760 6000 615856
rect 578000 615760 582820 615856
rect 1104 615216 6000 615312
rect 578000 615216 582820 615312
rect 1104 614672 6000 614768
rect 578000 614672 582820 614768
rect 1104 614128 6000 614224
rect 578000 614128 582820 614224
rect 1104 613584 6000 613680
rect 578000 613584 582820 613680
rect 1104 613040 6000 613136
rect 578000 613040 582820 613136
rect 1104 612496 6000 612592
rect 578000 612496 582820 612592
rect 1104 611952 6000 612048
rect 578000 611952 582820 612048
rect 1104 611408 6000 611504
rect 578000 611408 582820 611504
rect 2774 610988 2780 611040
rect 2832 611028 2838 611040
rect 5442 611028 5448 611040
rect 2832 611000 5448 611028
rect 2832 610988 2838 611000
rect 5442 610988 5448 611000
rect 5500 610988 5506 611040
rect 1104 610864 6000 610960
rect 578000 610864 582820 610960
rect 1104 610320 6000 610416
rect 578000 610320 582820 610416
rect 1104 609776 6000 609872
rect 578000 609776 582820 609872
rect 1104 609232 6000 609328
rect 578000 609232 582820 609328
rect 1104 608688 6000 608784
rect 578000 608688 582820 608784
rect 1104 608144 6000 608240
rect 578000 608144 582820 608240
rect 1104 607600 6000 607696
rect 578000 607600 582820 607696
rect 1104 607056 6000 607152
rect 578000 607056 582820 607152
rect 1104 606512 6000 606608
rect 578000 606512 582820 606608
rect 1104 605968 6000 606064
rect 578000 605968 582820 606064
rect 1104 605424 6000 605520
rect 578000 605424 582820 605520
rect 1104 604880 6000 604976
rect 578000 604880 582820 604976
rect 1104 604336 6000 604432
rect 578000 604336 582820 604432
rect 578142 604256 578148 604308
rect 578200 604296 578206 604308
rect 579614 604296 579620 604308
rect 578200 604268 579620 604296
rect 578200 604256 578206 604268
rect 579614 604256 579620 604268
rect 579672 604256 579678 604308
rect 1104 603792 6000 603888
rect 578000 603792 582820 603888
rect 1104 603248 6000 603344
rect 578000 603248 582820 603344
rect 1104 602704 6000 602800
rect 578000 602704 582820 602800
rect 1104 602160 6000 602256
rect 578000 602160 582820 602256
rect 1104 601616 6000 601712
rect 578000 601616 582820 601712
rect 1104 601072 6000 601168
rect 578000 601072 582820 601168
rect 1104 600528 6000 600624
rect 578000 600528 582820 600624
rect 1104 599984 6000 600080
rect 578000 599984 582820 600080
rect 1104 599440 6000 599536
rect 578000 599440 582820 599536
rect 1104 598896 6000 598992
rect 578000 598896 582820 598992
rect 1104 598352 6000 598448
rect 578000 598352 582820 598448
rect 1104 597808 6000 597904
rect 578000 597808 582820 597904
rect 1104 597264 6000 597360
rect 578000 597264 582820 597360
rect 1104 596720 6000 596816
rect 578000 596720 582820 596816
rect 1104 596176 6000 596272
rect 578000 596176 582820 596272
rect 3050 596028 3056 596080
rect 3108 596068 3114 596080
rect 7282 596068 7288 596080
rect 3108 596040 7288 596068
rect 3108 596028 3114 596040
rect 7282 596028 7288 596040
rect 7340 596028 7346 596080
rect 1104 595632 6000 595728
rect 578000 595632 582820 595728
rect 1104 595088 6000 595184
rect 578000 595088 582820 595184
rect 1104 594544 6000 594640
rect 578000 594544 582820 594640
rect 1104 594000 6000 594096
rect 578000 594000 582820 594096
rect 1104 593456 6000 593552
rect 578000 593456 582820 593552
rect 1104 592912 6000 593008
rect 578000 592912 582820 593008
rect 1104 592368 6000 592464
rect 578000 592368 582820 592464
rect 1104 591824 6000 591920
rect 578000 591824 582820 591920
rect 1104 591280 6000 591376
rect 578000 591280 582820 591376
rect 1104 590736 6000 590832
rect 578000 590736 582820 590832
rect 1104 590192 6000 590288
rect 578000 590192 582820 590288
rect 1104 589648 6000 589744
rect 578000 589648 582820 589744
rect 1104 589104 6000 589200
rect 578000 589104 582820 589200
rect 1104 588560 6000 588656
rect 578000 588560 582820 588656
rect 1104 588016 6000 588112
rect 578000 588016 582820 588112
rect 1104 587472 6000 587568
rect 578000 587472 582820 587568
rect 1104 586928 6000 587024
rect 578000 586928 582820 587024
rect 1104 586384 6000 586480
rect 578000 586384 582820 586480
rect 1104 585840 6000 585936
rect 578000 585840 582820 585936
rect 1104 585296 6000 585392
rect 578000 585296 582820 585392
rect 1104 584752 6000 584848
rect 578000 584752 582820 584848
rect 1104 584208 6000 584304
rect 578000 584208 582820 584304
rect 1104 583664 6000 583760
rect 578000 583664 582820 583760
rect 1104 583120 6000 583216
rect 578000 583120 582820 583216
rect 1104 582576 6000 582672
rect 578000 582576 582820 582672
rect 1104 582032 6000 582128
rect 578000 582032 582820 582128
rect 1104 581488 6000 581584
rect 578000 581488 582820 581584
rect 1104 580944 6000 581040
rect 578000 580944 582820 581040
rect 575382 580864 575388 580916
rect 575440 580904 575446 580916
rect 580166 580904 580172 580916
rect 575440 580876 580172 580904
rect 575440 580864 575446 580876
rect 580166 580864 580172 580876
rect 580224 580864 580230 580916
rect 1104 580400 6000 580496
rect 578000 580400 582820 580496
rect 1104 579856 6000 579952
rect 578000 579856 582820 579952
rect 1104 579312 6000 579408
rect 578000 579312 582820 579408
rect 1104 578768 6000 578864
rect 578000 578768 582820 578864
rect 1104 578224 6000 578320
rect 578000 578224 582820 578320
rect 1104 577680 6000 577776
rect 578000 577680 582820 577776
rect 1104 577136 6000 577232
rect 578000 577136 582820 577232
rect 1104 576592 6000 576688
rect 578000 576592 582820 576688
rect 1104 576048 6000 576144
rect 578000 576048 582820 576144
rect 1104 575504 6000 575600
rect 578000 575504 582820 575600
rect 1104 574960 6000 575056
rect 578000 574960 582820 575056
rect 1104 574416 6000 574512
rect 578000 574416 582820 574512
rect 1104 573872 6000 573968
rect 578000 573872 582820 573968
rect 1104 573328 6000 573424
rect 578000 573328 582820 573424
rect 1104 572784 6000 572880
rect 578000 572784 582820 572880
rect 1104 572240 6000 572336
rect 578000 572240 582820 572336
rect 1104 571696 6000 571792
rect 578000 571696 582820 571792
rect 1104 571152 6000 571248
rect 578000 571152 582820 571248
rect 1104 570608 6000 570704
rect 578000 570608 582820 570704
rect 1104 570064 6000 570160
rect 578000 570064 582820 570160
rect 1104 569520 6000 569616
rect 578000 569520 582820 569616
rect 1104 568976 6000 569072
rect 578000 568976 582820 569072
rect 1104 568432 6000 568528
rect 578000 568432 582820 568528
rect 1104 567888 6000 567984
rect 578000 567888 582820 567984
rect 2958 567468 2964 567520
rect 3016 567508 3022 567520
rect 5902 567508 5908 567520
rect 3016 567480 5908 567508
rect 3016 567468 3022 567480
rect 5902 567468 5908 567480
rect 5960 567468 5966 567520
rect 1104 567344 6000 567440
rect 578000 567344 582820 567440
rect 1104 566800 6000 566896
rect 578000 566800 582820 566896
rect 1104 566256 6000 566352
rect 578000 566256 582820 566352
rect 1104 565712 6000 565808
rect 578000 565712 582820 565808
rect 1104 565168 6000 565264
rect 578000 565168 582820 565264
rect 1104 564624 6000 564720
rect 578000 564624 582820 564720
rect 1104 564080 6000 564176
rect 578000 564080 582820 564176
rect 1104 563536 6000 563632
rect 578000 563536 582820 563632
rect 1104 562992 6000 563088
rect 578000 562992 582820 563088
rect 1104 562448 6000 562544
rect 578000 562448 582820 562544
rect 1104 561904 6000 562000
rect 578000 561904 582820 562000
rect 1104 561360 6000 561456
rect 578000 561360 582820 561456
rect 1104 560816 6000 560912
rect 578000 560816 582820 560912
rect 1104 560272 6000 560368
rect 578000 560272 582820 560368
rect 1104 559728 6000 559824
rect 578000 559728 582820 559824
rect 1104 559184 6000 559280
rect 578000 559184 582820 559280
rect 1104 558640 6000 558736
rect 578000 558640 582820 558736
rect 1104 558096 6000 558192
rect 578000 558096 582820 558192
rect 1104 557552 6000 557648
rect 578000 557552 582820 557648
rect 578050 557336 578056 557388
rect 578108 557376 578114 557388
rect 579614 557376 579620 557388
rect 578108 557348 579620 557376
rect 578108 557336 578114 557348
rect 579614 557336 579620 557348
rect 579672 557336 579678 557388
rect 1104 557008 6000 557104
rect 578000 557008 582820 557104
rect 1104 556464 6000 556560
rect 578000 556464 582820 556560
rect 1104 555920 6000 556016
rect 578000 555920 582820 556016
rect 1104 555376 6000 555472
rect 578000 555376 582820 555472
rect 1104 554832 6000 554928
rect 578000 554832 582820 554928
rect 1104 554288 6000 554384
rect 578000 554288 582820 554384
rect 1104 553744 6000 553840
rect 578000 553744 582820 553840
rect 1104 553200 6000 553296
rect 578000 553200 582820 553296
rect 1104 552656 6000 552752
rect 578000 552656 582820 552752
rect 1104 552112 6000 552208
rect 578000 552112 582820 552208
rect 1104 551568 6000 551664
rect 578000 551568 582820 551664
rect 1104 551024 6000 551120
rect 578000 551024 582820 551120
rect 1104 550480 6000 550576
rect 578000 550480 582820 550576
rect 1104 549936 6000 550032
rect 578000 549936 582820 550032
rect 1104 549392 6000 549488
rect 578000 549392 582820 549488
rect 1104 548848 6000 548944
rect 578000 548848 582820 548944
rect 1104 548304 6000 548400
rect 578000 548304 582820 548400
rect 1104 547760 6000 547856
rect 578000 547760 582820 547856
rect 1104 547216 6000 547312
rect 578000 547216 582820 547312
rect 1104 546672 6000 546768
rect 578000 546672 582820 546768
rect 1104 546128 6000 546224
rect 578000 546128 582820 546224
rect 1104 545584 6000 545680
rect 578000 545584 582820 545680
rect 1104 545040 6000 545136
rect 578000 545040 582820 545136
rect 1104 544496 6000 544592
rect 578000 544496 582820 544592
rect 1104 543952 6000 544048
rect 578000 543952 582820 544048
rect 1104 543408 6000 543504
rect 578000 543408 582820 543504
rect 1104 542864 6000 542960
rect 578000 542864 582820 542960
rect 1104 542320 6000 542416
rect 578000 542320 582820 542416
rect 1104 541776 6000 541872
rect 578000 541776 582820 541872
rect 1104 541232 6000 541328
rect 578000 541232 582820 541328
rect 1104 540688 6000 540784
rect 578000 540688 582820 540784
rect 1104 540144 6000 540240
rect 578000 540144 582820 540240
rect 1104 539600 6000 539696
rect 578000 539600 582820 539696
rect 1104 539056 6000 539152
rect 578000 539056 582820 539152
rect 1104 538512 6000 538608
rect 578000 538512 582820 538608
rect 1104 537968 6000 538064
rect 578000 537968 582820 538064
rect 1104 537424 6000 537520
rect 578000 537424 582820 537520
rect 1104 536880 6000 536976
rect 578000 536880 582820 536976
rect 1104 536336 6000 536432
rect 578000 536336 582820 536432
rect 1104 535792 6000 535888
rect 578000 535792 582820 535888
rect 1104 535248 6000 535344
rect 578000 535248 582820 535344
rect 1104 534704 6000 534800
rect 578000 534704 582820 534800
rect 1104 534160 6000 534256
rect 578000 534160 582820 534256
rect 577958 534012 577964 534064
rect 578016 534052 578022 534064
rect 579706 534052 579712 534064
rect 578016 534024 579712 534052
rect 578016 534012 578022 534024
rect 579706 534012 579712 534024
rect 579764 534012 579770 534064
rect 1104 533616 6000 533712
rect 578000 533616 582820 533712
rect 1104 533072 6000 533168
rect 578000 533072 582820 533168
rect 1104 532528 6000 532624
rect 578000 532528 582820 532624
rect 1104 531984 6000 532080
rect 578000 531984 582820 532080
rect 1104 531440 6000 531536
rect 578000 531440 582820 531536
rect 1104 530896 6000 530992
rect 578000 530896 582820 530992
rect 1104 530352 6000 530448
rect 578000 530352 582820 530448
rect 1104 529808 6000 529904
rect 578000 529808 582820 529904
rect 1104 529264 6000 529360
rect 578000 529264 582820 529360
rect 1104 528720 6000 528816
rect 578000 528720 582820 528816
rect 1104 528176 6000 528272
rect 578000 528176 582820 528272
rect 1104 527632 6000 527728
rect 578000 527632 582820 527728
rect 1104 527088 6000 527184
rect 578000 527088 582820 527184
rect 1104 526544 6000 526640
rect 578000 526544 582820 526640
rect 1104 526000 6000 526096
rect 578000 526000 582820 526096
rect 1104 525456 6000 525552
rect 578000 525456 582820 525552
rect 1104 524912 6000 525008
rect 578000 524912 582820 525008
rect 1104 524368 6000 524464
rect 578000 524368 582820 524464
rect 1104 523824 6000 523920
rect 578000 523824 582820 523920
rect 1104 523280 6000 523376
rect 578000 523280 582820 523376
rect 1104 522736 6000 522832
rect 578000 522736 582820 522832
rect 1104 522192 6000 522288
rect 578000 522192 582820 522288
rect 1104 521648 6000 521744
rect 578000 521648 582820 521744
rect 1104 521104 6000 521200
rect 578000 521104 582820 521200
rect 1104 520560 6000 520656
rect 578000 520560 582820 520656
rect 1104 520016 6000 520112
rect 578000 520016 582820 520112
rect 1104 519472 6000 519568
rect 578000 519472 582820 519568
rect 1104 518928 6000 519024
rect 578000 518928 582820 519024
rect 1104 518384 6000 518480
rect 578000 518384 582820 518480
rect 1104 517840 6000 517936
rect 578000 517840 582820 517936
rect 1104 517296 6000 517392
rect 578000 517296 582820 517392
rect 1104 516752 6000 516848
rect 578000 516752 582820 516848
rect 1104 516208 6000 516304
rect 578000 516208 582820 516304
rect 1104 515664 6000 515760
rect 578000 515664 582820 515760
rect 1104 515120 6000 515216
rect 578000 515120 582820 515216
rect 1104 514576 6000 514672
rect 578000 514576 582820 514672
rect 1104 514032 6000 514128
rect 578000 514032 582820 514128
rect 1104 513488 6000 513584
rect 578000 513488 582820 513584
rect 1104 512944 6000 513040
rect 578000 512944 582820 513040
rect 1104 512400 6000 512496
rect 578000 512400 582820 512496
rect 1104 511856 6000 511952
rect 578000 511856 582820 511952
rect 1104 511312 6000 511408
rect 578000 511312 582820 511408
rect 1104 510768 6000 510864
rect 578000 510768 582820 510864
rect 576026 510552 576032 510604
rect 576084 510592 576090 510604
rect 580166 510592 580172 510604
rect 576084 510564 580172 510592
rect 576084 510552 576090 510564
rect 580166 510552 580172 510564
rect 580224 510552 580230 510604
rect 3050 510348 3056 510400
rect 3108 510388 3114 510400
rect 5994 510388 6000 510400
rect 3108 510360 6000 510388
rect 3108 510348 3114 510360
rect 5994 510348 6000 510360
rect 6052 510348 6058 510400
rect 1104 510224 6000 510320
rect 578000 510224 582820 510320
rect 1104 509680 6000 509776
rect 578000 509680 582820 509776
rect 1104 509136 6000 509232
rect 578000 509136 582820 509232
rect 1104 508592 6000 508688
rect 578000 508592 582820 508688
rect 1104 508048 6000 508144
rect 578000 508048 582820 508144
rect 1104 507504 6000 507600
rect 578000 507504 582820 507600
rect 1104 506960 6000 507056
rect 578000 506960 582820 507056
rect 1104 506416 6000 506512
rect 578000 506416 582820 506512
rect 1104 505872 6000 505968
rect 578000 505872 582820 505968
rect 1104 505328 6000 505424
rect 578000 505328 582820 505424
rect 1104 504784 6000 504880
rect 578000 504784 582820 504880
rect 1104 504240 6000 504336
rect 578000 504240 582820 504336
rect 1104 503696 6000 503792
rect 578000 503696 582820 503792
rect 1104 503152 6000 503248
rect 578000 503152 582820 503248
rect 1104 502608 6000 502704
rect 578000 502608 582820 502704
rect 1104 502064 6000 502160
rect 578000 502064 582820 502160
rect 1104 501520 6000 501616
rect 578000 501520 582820 501616
rect 1104 500976 6000 501072
rect 578000 500976 582820 501072
rect 1104 500432 6000 500528
rect 578000 500432 582820 500528
rect 1104 499888 6000 499984
rect 578000 499888 582820 499984
rect 1104 499344 6000 499440
rect 578000 499344 582820 499440
rect 577866 499060 577872 499112
rect 577924 499100 577930 499112
rect 580166 499100 580172 499112
rect 577924 499072 580172 499100
rect 577924 499060 577930 499072
rect 580166 499060 580172 499072
rect 580224 499060 580230 499112
rect 1104 498800 6000 498896
rect 578000 498800 582820 498896
rect 1104 498256 6000 498352
rect 578000 498256 582820 498352
rect 1104 497712 6000 497808
rect 578000 497712 582820 497808
rect 1104 497168 6000 497264
rect 578000 497168 582820 497264
rect 1104 496624 6000 496720
rect 578000 496624 582820 496720
rect 1104 496080 6000 496176
rect 578000 496080 582820 496176
rect 1104 495536 6000 495632
rect 578000 495536 582820 495632
rect 1104 494992 6000 495088
rect 578000 494992 582820 495088
rect 1104 494448 6000 494544
rect 578000 494448 582820 494544
rect 1104 493904 6000 494000
rect 578000 493904 582820 494000
rect 1104 493360 6000 493456
rect 578000 493360 582820 493456
rect 1104 492816 6000 492912
rect 578000 492816 582820 492912
rect 1104 492272 6000 492368
rect 578000 492272 582820 492368
rect 1104 491728 6000 491824
rect 578000 491728 582820 491824
rect 1104 491184 6000 491280
rect 578000 491184 582820 491280
rect 1104 490640 6000 490736
rect 578000 490640 582820 490736
rect 1104 490096 6000 490192
rect 578000 490096 582820 490192
rect 1104 489552 6000 489648
rect 578000 489552 582820 489648
rect 1104 489008 6000 489104
rect 578000 489008 582820 489104
rect 1104 488464 6000 488560
rect 578000 488464 582820 488560
rect 1104 487920 6000 488016
rect 578000 487920 582820 488016
rect 1104 487376 6000 487472
rect 578000 487376 582820 487472
rect 576762 487092 576768 487144
rect 576820 487132 576826 487144
rect 579982 487132 579988 487144
rect 576820 487104 579988 487132
rect 576820 487092 576826 487104
rect 579982 487092 579988 487104
rect 580040 487092 580046 487144
rect 1104 486832 6000 486928
rect 578000 486832 582820 486928
rect 1104 486288 6000 486384
rect 578000 486288 582820 486384
rect 1104 485744 6000 485840
rect 578000 485744 582820 485840
rect 1104 485200 6000 485296
rect 578000 485200 582820 485296
rect 1104 484656 6000 484752
rect 578000 484656 582820 484752
rect 1104 484112 6000 484208
rect 578000 484112 582820 484208
rect 1104 483568 6000 483664
rect 578000 483568 582820 483664
rect 1104 483024 6000 483120
rect 578000 483024 582820 483120
rect 1104 482480 6000 482576
rect 578000 482480 582820 482576
rect 1104 481936 6000 482032
rect 578000 481936 582820 482032
rect 1104 481392 6000 481488
rect 578000 481392 582820 481488
rect 3234 481108 3240 481160
rect 3292 481148 3298 481160
rect 7374 481148 7380 481160
rect 3292 481120 7380 481148
rect 3292 481108 3298 481120
rect 7374 481108 7380 481120
rect 7432 481108 7438 481160
rect 1104 480848 6000 480944
rect 578000 480848 582820 480944
rect 1104 480304 6000 480400
rect 578000 480304 582820 480400
rect 1104 479760 6000 479856
rect 578000 479760 582820 479856
rect 1104 479216 6000 479312
rect 578000 479216 582820 479312
rect 1104 478672 6000 478768
rect 578000 478672 582820 478768
rect 1104 478128 6000 478224
rect 578000 478128 582820 478224
rect 1104 477584 6000 477680
rect 578000 477584 582820 477680
rect 1104 477040 6000 477136
rect 578000 477040 582820 477136
rect 1104 476496 6000 476592
rect 578000 476496 582820 476592
rect 1104 475952 6000 476048
rect 578000 475952 582820 476048
rect 1104 475408 6000 475504
rect 578000 475408 582820 475504
rect 1104 474864 6000 474960
rect 578000 474864 582820 474960
rect 1104 474320 6000 474416
rect 578000 474320 582820 474416
rect 1104 473776 6000 473872
rect 578000 473776 582820 473872
rect 1104 473232 6000 473328
rect 578000 473232 582820 473328
rect 1104 472688 6000 472784
rect 578000 472688 582820 472784
rect 1104 472144 6000 472240
rect 578000 472144 582820 472240
rect 1104 471600 6000 471696
rect 578000 471600 582820 471696
rect 1104 471056 6000 471152
rect 578000 471056 582820 471152
rect 1104 470512 6000 470608
rect 578000 470512 582820 470608
rect 1104 469968 6000 470064
rect 578000 469968 582820 470064
rect 1104 469424 6000 469520
rect 578000 469424 582820 469520
rect 1104 468880 6000 468976
rect 578000 468880 582820 468976
rect 1104 468336 6000 468432
rect 578000 468336 582820 468432
rect 1104 467792 6000 467888
rect 578000 467792 582820 467888
rect 1104 467248 6000 467344
rect 578000 467248 582820 467344
rect 1104 466704 6000 466800
rect 578000 466704 582820 466800
rect 1104 466160 6000 466256
rect 578000 466160 582820 466256
rect 1104 465616 6000 465712
rect 578000 465616 582820 465712
rect 1104 465072 6000 465168
rect 578000 465072 582820 465168
rect 1104 464528 6000 464624
rect 578000 464528 582820 464624
rect 1104 463984 6000 464080
rect 578000 463984 582820 464080
rect 577774 463632 577780 463684
rect 577832 463672 577838 463684
rect 579614 463672 579620 463684
rect 577832 463644 579620 463672
rect 577832 463632 577838 463644
rect 579614 463632 579620 463644
rect 579672 463632 579678 463684
rect 1104 463440 6000 463536
rect 578000 463440 582820 463536
rect 1104 462896 6000 462992
rect 578000 462896 582820 462992
rect 1104 462352 6000 462448
rect 578000 462352 582820 462448
rect 1104 461808 6000 461904
rect 578000 461808 582820 461904
rect 1104 461264 6000 461360
rect 578000 461264 582820 461360
rect 1104 460720 6000 460816
rect 578000 460720 582820 460816
rect 1104 460176 6000 460272
rect 578000 460176 582820 460272
rect 1104 459632 6000 459728
rect 578000 459632 582820 459728
rect 1104 459088 6000 459184
rect 578000 459088 582820 459184
rect 1104 458544 6000 458640
rect 578000 458544 582820 458640
rect 1104 458000 6000 458096
rect 578000 458000 582820 458096
rect 1104 457456 6000 457552
rect 578000 457456 582820 457552
rect 1104 456912 6000 457008
rect 578000 456912 582820 457008
rect 1104 456368 6000 456464
rect 578000 456368 582820 456464
rect 1104 455824 6000 455920
rect 578000 455824 582820 455920
rect 1104 455280 6000 455376
rect 578000 455280 582820 455376
rect 1104 454736 6000 454832
rect 578000 454736 582820 454832
rect 1104 454192 6000 454288
rect 578000 454192 582820 454288
rect 1104 453648 6000 453744
rect 578000 453648 582820 453744
rect 1104 453104 6000 453200
rect 578000 453104 582820 453200
rect 1104 452560 6000 452656
rect 578000 452560 582820 452656
rect 3050 452412 3056 452464
rect 3108 452452 3114 452464
rect 6086 452452 6092 452464
rect 3108 452424 6092 452452
rect 3108 452412 3114 452424
rect 6086 452412 6092 452424
rect 6144 452412 6150 452464
rect 1104 452016 6000 452112
rect 578000 452016 582820 452112
rect 1104 451472 6000 451568
rect 578000 451472 582820 451568
rect 1104 450928 6000 451024
rect 578000 450928 582820 451024
rect 1104 450384 6000 450480
rect 578000 450384 582820 450480
rect 1104 449840 6000 449936
rect 578000 449840 582820 449936
rect 1104 449296 6000 449392
rect 578000 449296 582820 449392
rect 1104 448752 6000 448848
rect 578000 448752 582820 448848
rect 1104 448208 6000 448304
rect 578000 448208 582820 448304
rect 1104 447664 6000 447760
rect 578000 447664 582820 447760
rect 1104 447120 6000 447216
rect 578000 447120 582820 447216
rect 1104 446576 6000 446672
rect 578000 446576 582820 446672
rect 1104 446032 6000 446128
rect 578000 446032 582820 446128
rect 1104 445488 6000 445584
rect 578000 445488 582820 445584
rect 1104 444944 6000 445040
rect 578000 444944 582820 445040
rect 1104 444400 6000 444496
rect 578000 444400 582820 444496
rect 1104 443856 6000 443952
rect 578000 443856 582820 443952
rect 1104 443312 6000 443408
rect 578000 443312 582820 443408
rect 1104 442768 6000 442864
rect 578000 442768 582820 442864
rect 1104 442224 6000 442320
rect 578000 442224 582820 442320
rect 1104 441680 6000 441776
rect 578000 441680 582820 441776
rect 1104 441136 6000 441232
rect 578000 441136 582820 441232
rect 1104 440592 6000 440688
rect 578000 440592 582820 440688
rect 3970 440240 3976 440292
rect 4028 440280 4034 440292
rect 5350 440280 5356 440292
rect 4028 440252 5356 440280
rect 4028 440240 4034 440252
rect 5350 440240 5356 440252
rect 5408 440240 5414 440292
rect 576670 440172 576676 440224
rect 576728 440212 576734 440224
rect 579982 440212 579988 440224
rect 576728 440184 579988 440212
rect 576728 440172 576734 440184
rect 579982 440172 579988 440184
rect 580040 440172 580046 440224
rect 1104 440048 6000 440144
rect 578000 440048 582820 440144
rect 1104 439504 6000 439600
rect 578000 439504 582820 439600
rect 1104 438960 6000 439056
rect 578000 438960 582820 439056
rect 1104 438416 6000 438512
rect 578000 438416 582820 438512
rect 1104 437872 6000 437968
rect 578000 437872 582820 437968
rect 1104 437328 6000 437424
rect 578000 437328 582820 437424
rect 1104 436784 6000 436880
rect 578000 436784 582820 436880
rect 1104 436240 6000 436336
rect 578000 436240 582820 436336
rect 1104 435696 6000 435792
rect 578000 435696 582820 435792
rect 1104 435152 6000 435248
rect 578000 435152 582820 435248
rect 1104 434608 6000 434704
rect 578000 434608 582820 434704
rect 1104 434064 6000 434160
rect 578000 434064 582820 434160
rect 1104 433520 6000 433616
rect 578000 433520 582820 433616
rect 1104 432976 6000 433072
rect 578000 432976 582820 433072
rect 1104 432432 6000 432528
rect 578000 432432 582820 432528
rect 1104 431888 6000 431984
rect 578000 431888 582820 431984
rect 1104 431344 6000 431440
rect 578000 431344 582820 431440
rect 1104 430800 6000 430896
rect 578000 430800 582820 430896
rect 1104 430256 6000 430352
rect 578000 430256 582820 430352
rect 1104 429712 6000 429808
rect 578000 429712 582820 429808
rect 1104 429168 6000 429264
rect 578000 429168 582820 429264
rect 1104 428624 6000 428720
rect 578000 428624 582820 428720
rect 1104 428080 6000 428176
rect 578000 428080 582820 428176
rect 1104 427536 6000 427632
rect 578000 427536 582820 427632
rect 1104 426992 6000 427088
rect 578000 426992 582820 427088
rect 1104 426448 6000 426544
rect 578000 426448 582820 426544
rect 1104 425904 6000 426000
rect 578000 425904 582820 426000
rect 1104 425360 6000 425456
rect 578000 425360 582820 425456
rect 1104 424816 6000 424912
rect 578000 424816 582820 424912
rect 1104 424272 6000 424368
rect 578000 424272 582820 424368
rect 3326 423920 3332 423972
rect 3384 423960 3390 423972
rect 6822 423960 6828 423972
rect 3384 423932 6828 423960
rect 3384 423920 3390 423932
rect 6822 423920 6828 423932
rect 6880 423920 6886 423972
rect 1104 423728 6000 423824
rect 578000 423728 582820 423824
rect 1104 423184 6000 423280
rect 578000 423184 582820 423280
rect 1104 422640 6000 422736
rect 578000 422640 582820 422736
rect 1104 422096 6000 422192
rect 578000 422096 582820 422192
rect 1104 421552 6000 421648
rect 578000 421552 582820 421648
rect 1104 421008 6000 421104
rect 578000 421008 582820 421104
rect 1104 420464 6000 420560
rect 578000 420464 582820 420560
rect 1104 419920 6000 420016
rect 578000 419920 582820 420016
rect 1104 419376 6000 419472
rect 578000 419376 582820 419472
rect 1104 418832 6000 418928
rect 578000 418832 582820 418928
rect 1104 418288 6000 418384
rect 578000 418288 582820 418384
rect 1104 417744 6000 417840
rect 578000 417744 582820 417840
rect 1104 417200 6000 417296
rect 578000 417200 582820 417296
rect 1104 416656 6000 416752
rect 578000 416656 582820 416752
rect 576578 416576 576584 416628
rect 576636 416616 576642 416628
rect 580166 416616 580172 416628
rect 576636 416588 580172 416616
rect 576636 416576 576642 416588
rect 580166 416576 580172 416588
rect 580224 416576 580230 416628
rect 1104 416112 6000 416208
rect 578000 416112 582820 416208
rect 1104 415568 6000 415664
rect 578000 415568 582820 415664
rect 1104 415024 6000 415120
rect 578000 415024 582820 415120
rect 1104 414480 6000 414576
rect 578000 414480 582820 414576
rect 1104 413936 6000 414032
rect 578000 413936 582820 414032
rect 1104 413392 6000 413488
rect 578000 413392 582820 413488
rect 1104 412848 6000 412944
rect 578000 412848 582820 412944
rect 1104 412304 6000 412400
rect 578000 412304 582820 412400
rect 1104 411760 6000 411856
rect 578000 411760 582820 411856
rect 1104 411216 6000 411312
rect 578000 411216 582820 411312
rect 1104 410672 6000 410768
rect 578000 410672 582820 410768
rect 1104 410128 6000 410224
rect 578000 410128 582820 410224
rect 1104 409584 6000 409680
rect 578000 409584 582820 409680
rect 1104 409040 6000 409136
rect 578000 409040 582820 409136
rect 1104 408496 6000 408592
rect 578000 408496 582820 408592
rect 1104 407952 6000 408048
rect 578000 407952 582820 408048
rect 1104 407408 6000 407504
rect 578000 407408 582820 407504
rect 1104 406864 6000 406960
rect 578000 406864 582820 406960
rect 1104 406320 6000 406416
rect 578000 406320 582820 406416
rect 1104 405776 6000 405872
rect 578000 405776 582820 405872
rect 1104 405232 6000 405328
rect 578000 405232 582820 405328
rect 1104 404688 6000 404784
rect 578000 404688 582820 404784
rect 1104 404144 6000 404240
rect 578000 404144 582820 404240
rect 1104 403600 6000 403696
rect 578000 403600 582820 403696
rect 1104 403056 6000 403152
rect 578000 403056 582820 403152
rect 1104 402512 6000 402608
rect 578000 402512 582820 402608
rect 1104 401968 6000 402064
rect 578000 401968 582820 402064
rect 1104 401424 6000 401520
rect 578000 401424 582820 401520
rect 1104 400880 6000 400976
rect 578000 400880 582820 400976
rect 1104 400336 6000 400432
rect 578000 400336 582820 400432
rect 1104 399792 6000 399888
rect 578000 399792 582820 399888
rect 1104 399248 6000 399344
rect 578000 399248 582820 399344
rect 1104 398704 6000 398800
rect 578000 398704 582820 398800
rect 1104 398160 6000 398256
rect 578000 398160 582820 398256
rect 1104 397616 6000 397712
rect 578000 397616 582820 397712
rect 1104 397072 6000 397168
rect 578000 397072 582820 397168
rect 1104 396528 6000 396624
rect 578000 396528 582820 396624
rect 1104 395984 6000 396080
rect 578000 395984 582820 396080
rect 3326 395700 3332 395752
rect 3384 395740 3390 395752
rect 6730 395740 6736 395752
rect 3384 395712 6736 395740
rect 3384 395700 3390 395712
rect 6730 395700 6736 395712
rect 6788 395700 6794 395752
rect 1104 395440 6000 395536
rect 578000 395440 582820 395536
rect 1104 394896 6000 394992
rect 578000 394896 582820 394992
rect 1104 394352 6000 394448
rect 578000 394352 582820 394448
rect 1104 393808 6000 393904
rect 578000 393808 582820 393904
rect 1104 393264 6000 393360
rect 578000 393264 582820 393360
rect 1104 392720 6000 392816
rect 578000 392720 582820 392816
rect 1104 392176 6000 392272
rect 578000 392176 582820 392272
rect 1104 391632 6000 391728
rect 578000 391632 582820 391728
rect 1104 391088 6000 391184
rect 578000 391088 582820 391184
rect 1104 390544 6000 390640
rect 578000 390544 582820 390640
rect 1104 390000 6000 390096
rect 578000 390000 582820 390096
rect 1104 389456 6000 389552
rect 578000 389456 582820 389552
rect 1104 388912 6000 389008
rect 578000 388912 582820 389008
rect 1104 388368 6000 388464
rect 578000 388368 582820 388464
rect 1104 387824 6000 387920
rect 578000 387824 582820 387920
rect 1104 387280 6000 387376
rect 578000 387280 582820 387376
rect 1104 386736 6000 386832
rect 578000 386736 582820 386832
rect 1104 386192 6000 386288
rect 578000 386192 582820 386288
rect 1104 385648 6000 385744
rect 578000 385648 582820 385744
rect 1104 385104 6000 385200
rect 578000 385104 582820 385200
rect 1104 384560 6000 384656
rect 578000 384560 582820 384656
rect 1104 384016 6000 384112
rect 578000 384016 582820 384112
rect 1104 383472 6000 383568
rect 578000 383472 582820 383568
rect 1104 382928 6000 383024
rect 578000 382928 582820 383024
rect 1104 382384 6000 382480
rect 578000 382384 582820 382480
rect 1104 381840 6000 381936
rect 578000 381840 582820 381936
rect 1104 381296 6000 381392
rect 578000 381296 582820 381392
rect 1104 380752 6000 380848
rect 578000 380752 582820 380848
rect 1104 380208 6000 380304
rect 578000 380208 582820 380304
rect 1104 379664 6000 379760
rect 578000 379664 582820 379760
rect 1104 379120 6000 379216
rect 578000 379120 582820 379216
rect 1104 378576 6000 378672
rect 578000 378576 582820 378672
rect 4062 378428 4068 378480
rect 4120 378468 4126 378480
rect 5258 378468 5264 378480
rect 4120 378440 5264 378468
rect 4120 378428 4126 378440
rect 5258 378428 5264 378440
rect 5316 378428 5322 378480
rect 1104 378032 6000 378128
rect 578000 378032 582820 378128
rect 1104 377488 6000 377584
rect 578000 377488 582820 377584
rect 1104 376944 6000 377040
rect 578000 376944 582820 377040
rect 1104 376400 6000 376496
rect 578000 376400 582820 376496
rect 1104 375856 6000 375952
rect 578000 375856 582820 375952
rect 1104 375312 6000 375408
rect 578000 375312 582820 375408
rect 1104 374768 6000 374864
rect 578000 374768 582820 374864
rect 1104 374224 6000 374320
rect 578000 374224 582820 374320
rect 1104 373680 6000 373776
rect 578000 373680 582820 373776
rect 1104 373136 6000 373232
rect 578000 373136 582820 373232
rect 1104 372592 6000 372688
rect 578000 372592 582820 372688
rect 1104 372048 6000 372144
rect 578000 372048 582820 372144
rect 1104 371504 6000 371600
rect 578000 371504 582820 371600
rect 1104 370960 6000 371056
rect 578000 370960 582820 371056
rect 1104 370416 6000 370512
rect 578000 370416 582820 370512
rect 1104 369872 6000 369968
rect 578000 369872 582820 369968
rect 1104 369328 6000 369424
rect 578000 369328 582820 369424
rect 1104 368784 6000 368880
rect 578000 368784 582820 368880
rect 1104 368240 6000 368336
rect 578000 368240 582820 368336
rect 1104 367696 6000 367792
rect 578000 367696 582820 367792
rect 1104 367152 6000 367248
rect 578000 367152 582820 367248
rect 1104 366608 6000 366704
rect 578000 366608 582820 366704
rect 3326 366188 3332 366240
rect 3384 366228 3390 366240
rect 7466 366228 7472 366240
rect 3384 366200 7472 366228
rect 3384 366188 3390 366200
rect 7466 366188 7472 366200
rect 7524 366188 7530 366240
rect 1104 366064 6000 366160
rect 578000 366064 582820 366160
rect 1104 365520 6000 365616
rect 578000 365520 582820 365616
rect 1104 364976 6000 365072
rect 578000 364976 582820 365072
rect 1104 364432 6000 364528
rect 578000 364432 582820 364528
rect 1104 363888 6000 363984
rect 578000 363888 582820 363984
rect 1104 363344 6000 363440
rect 578000 363344 582820 363440
rect 1104 362800 6000 362896
rect 578000 362800 582820 362896
rect 1104 362256 6000 362352
rect 578000 362256 582820 362352
rect 1104 361712 6000 361808
rect 578000 361712 582820 361808
rect 1104 361168 6000 361264
rect 578000 361168 582820 361264
rect 1104 360624 6000 360720
rect 578000 360624 582820 360720
rect 1104 360080 6000 360176
rect 578000 360080 582820 360176
rect 1104 359536 6000 359632
rect 578000 359536 582820 359632
rect 1104 358992 6000 359088
rect 578000 358992 582820 359088
rect 577682 358708 577688 358760
rect 577740 358748 577746 358760
rect 580810 358748 580816 358760
rect 577740 358720 580816 358748
rect 577740 358708 577746 358720
rect 580810 358708 580816 358720
rect 580868 358708 580874 358760
rect 1104 358448 6000 358544
rect 578000 358448 582820 358544
rect 1104 357904 6000 358000
rect 578000 357904 582820 358000
rect 1104 357360 6000 357456
rect 578000 357360 582820 357456
rect 1104 356816 6000 356912
rect 578000 356816 582820 356912
rect 1104 356272 6000 356368
rect 578000 356272 582820 356368
rect 1104 355728 6000 355824
rect 578000 355728 582820 355824
rect 1104 355184 6000 355280
rect 578000 355184 582820 355280
rect 1104 354640 6000 354736
rect 578000 354640 582820 354736
rect 1104 354096 6000 354192
rect 578000 354096 582820 354192
rect 1104 353552 6000 353648
rect 578000 353552 582820 353648
rect 1104 353008 6000 353104
rect 578000 353008 582820 353104
rect 1104 352464 6000 352560
rect 578000 352464 582820 352560
rect 1104 351920 6000 352016
rect 578000 351920 582820 352016
rect 1104 351376 6000 351472
rect 578000 351376 582820 351472
rect 1104 350832 6000 350928
rect 578000 350832 582820 350928
rect 1104 350288 6000 350384
rect 578000 350288 582820 350384
rect 1104 349744 6000 349840
rect 578000 349744 582820 349840
rect 1104 349200 6000 349296
rect 578000 349200 582820 349296
rect 1104 348656 6000 348752
rect 578000 348656 582820 348752
rect 1104 348112 6000 348208
rect 578000 348112 582820 348208
rect 1104 347568 6000 347664
rect 578000 347568 582820 347664
rect 1104 347024 6000 347120
rect 578000 347024 582820 347120
rect 1104 346480 6000 346576
rect 578000 346480 582820 346576
rect 576486 346332 576492 346384
rect 576544 346372 576550 346384
rect 579982 346372 579988 346384
rect 576544 346344 579988 346372
rect 576544 346332 576550 346344
rect 579982 346332 579988 346344
rect 580040 346332 580046 346384
rect 1104 345936 6000 346032
rect 578000 345936 582820 346032
rect 1104 345392 6000 345488
rect 578000 345392 582820 345488
rect 1104 344848 6000 344944
rect 578000 344848 582820 344944
rect 1104 344304 6000 344400
rect 578000 344304 582820 344400
rect 1104 343760 6000 343856
rect 578000 343760 582820 343856
rect 1104 343216 6000 343312
rect 578000 343216 582820 343312
rect 1104 342672 6000 342768
rect 578000 342672 582820 342768
rect 1104 342128 6000 342224
rect 578000 342128 582820 342224
rect 1104 341584 6000 341680
rect 578000 341584 582820 341680
rect 1104 341040 6000 341136
rect 578000 341040 582820 341136
rect 1104 340496 6000 340592
rect 578000 340496 582820 340592
rect 1104 339952 6000 340048
rect 578000 339952 582820 340048
rect 1104 339408 6000 339504
rect 578000 339408 582820 339504
rect 1104 338864 6000 338960
rect 578000 338864 582820 338960
rect 1104 338320 6000 338416
rect 578000 338320 582820 338416
rect 3326 337900 3332 337952
rect 3384 337940 3390 337952
rect 6638 337940 6644 337952
rect 3384 337912 6644 337940
rect 3384 337900 3390 337912
rect 6638 337900 6644 337912
rect 6696 337900 6702 337952
rect 1104 337776 6000 337872
rect 578000 337776 582820 337872
rect 1104 337232 6000 337328
rect 578000 337232 582820 337328
rect 1104 336688 6000 336784
rect 578000 336688 582820 336784
rect 1104 336144 6000 336240
rect 578000 336144 582820 336240
rect 1104 335600 6000 335696
rect 578000 335600 582820 335696
rect 1104 335056 6000 335152
rect 578000 335056 582820 335152
rect 1104 334512 6000 334608
rect 578000 334512 582820 334608
rect 1104 333968 6000 334064
rect 578000 333968 582820 334064
rect 1104 333424 6000 333520
rect 578000 333424 582820 333520
rect 1104 332880 6000 332976
rect 578000 332880 582820 332976
rect 1104 332336 6000 332432
rect 578000 332336 582820 332432
rect 1104 331792 6000 331888
rect 578000 331792 582820 331888
rect 1104 331248 6000 331344
rect 578000 331248 582820 331344
rect 1104 330704 6000 330800
rect 578000 330704 582820 330800
rect 1104 330160 6000 330256
rect 578000 330160 582820 330256
rect 1104 329616 6000 329712
rect 578000 329616 582820 329712
rect 1104 329072 6000 329168
rect 578000 329072 582820 329168
rect 1104 328528 6000 328624
rect 578000 328528 582820 328624
rect 1104 327984 6000 328080
rect 578000 327984 582820 328080
rect 1104 327440 6000 327536
rect 578000 327440 582820 327536
rect 1104 326896 6000 326992
rect 578000 326896 582820 326992
rect 1104 326352 6000 326448
rect 578000 326352 582820 326448
rect 1104 325808 6000 325904
rect 578000 325808 582820 325904
rect 1104 325264 6000 325360
rect 578000 325264 582820 325360
rect 1104 324720 6000 324816
rect 578000 324720 582820 324816
rect 1104 324176 6000 324272
rect 578000 324176 582820 324272
rect 2774 323892 2780 323944
rect 2832 323932 2838 323944
rect 5166 323932 5172 323944
rect 2832 323904 5172 323932
rect 2832 323892 2838 323904
rect 5166 323892 5172 323904
rect 5224 323892 5230 323944
rect 1104 323632 6000 323728
rect 578000 323632 582820 323728
rect 1104 323088 6000 323184
rect 578000 323088 582820 323184
rect 1104 322544 6000 322640
rect 578000 322544 582820 322640
rect 1104 322000 6000 322096
rect 578000 322000 582820 322096
rect 1104 321456 6000 321552
rect 578000 321456 582820 321552
rect 1104 320912 6000 321008
rect 578000 320912 582820 321008
rect 1104 320368 6000 320464
rect 578000 320368 582820 320464
rect 1104 319824 6000 319920
rect 578000 319824 582820 319920
rect 1104 319280 6000 319376
rect 578000 319280 582820 319376
rect 1104 318736 6000 318832
rect 578000 318736 582820 318832
rect 1104 318192 6000 318288
rect 578000 318192 582820 318288
rect 1104 317648 6000 317744
rect 578000 317648 582820 317744
rect 1104 317104 6000 317200
rect 578000 317104 582820 317200
rect 1104 316560 6000 316656
rect 578000 316560 582820 316656
rect 1104 316016 6000 316112
rect 578000 316016 582820 316112
rect 1104 315472 6000 315568
rect 578000 315472 582820 315568
rect 1104 314928 6000 315024
rect 578000 314928 582820 315024
rect 1104 314384 6000 314480
rect 578000 314384 582820 314480
rect 1104 313840 6000 313936
rect 578000 313840 582820 313936
rect 1104 313296 6000 313392
rect 578000 313296 582820 313392
rect 1104 312752 6000 312848
rect 578000 312752 582820 312848
rect 1104 312208 6000 312304
rect 578000 312208 582820 312304
rect 577590 311788 577596 311840
rect 577648 311828 577654 311840
rect 580810 311828 580816 311840
rect 577648 311800 580816 311828
rect 577648 311788 577654 311800
rect 580810 311788 580816 311800
rect 580868 311788 580874 311840
rect 1104 311664 6000 311760
rect 578000 311664 582820 311760
rect 1104 311120 6000 311216
rect 578000 311120 582820 311216
rect 1104 310576 6000 310672
rect 578000 310576 582820 310672
rect 1104 310032 6000 310128
rect 578000 310032 582820 310128
rect 1104 309488 6000 309584
rect 578000 309488 582820 309584
rect 1104 308944 6000 309040
rect 578000 308944 582820 309040
rect 1104 308400 6000 308496
rect 578000 308400 582820 308496
rect 1104 307856 6000 307952
rect 578000 307856 582820 307952
rect 1104 307312 6000 307408
rect 578000 307312 582820 307408
rect 1104 306768 6000 306864
rect 578000 306768 582820 306864
rect 1104 306224 6000 306320
rect 578000 306224 582820 306320
rect 1104 305680 6000 305776
rect 578000 305680 582820 305776
rect 1104 305136 6000 305232
rect 578000 305136 582820 305232
rect 1104 304592 6000 304688
rect 578000 304592 582820 304688
rect 1104 304048 6000 304144
rect 578000 304048 582820 304144
rect 1104 303504 6000 303600
rect 578000 303504 582820 303600
rect 1104 302960 6000 303056
rect 578000 302960 582820 303056
rect 1104 302416 6000 302512
rect 578000 302416 582820 302512
rect 1104 301872 6000 301968
rect 578000 301872 582820 301968
rect 1104 301328 6000 301424
rect 578000 301328 582820 301424
rect 1104 300784 6000 300880
rect 578000 300784 582820 300880
rect 1104 300240 6000 300336
rect 578000 300240 582820 300336
rect 1104 299696 6000 299792
rect 578000 299696 582820 299792
rect 575290 299412 575296 299464
rect 575348 299452 575354 299464
rect 579614 299452 579620 299464
rect 575348 299424 579620 299452
rect 575348 299412 575354 299424
rect 579614 299412 579620 299424
rect 579672 299412 579678 299464
rect 1104 299152 6000 299248
rect 578000 299152 582820 299248
rect 1104 298608 6000 298704
rect 578000 298608 582820 298704
rect 1104 298064 6000 298160
rect 578000 298064 582820 298160
rect 1104 297520 6000 297616
rect 578000 297520 582820 297616
rect 1104 296976 6000 297072
rect 578000 296976 582820 297072
rect 1104 296432 6000 296528
rect 578000 296432 582820 296528
rect 1104 295888 6000 295984
rect 578000 295888 582820 295984
rect 1104 295344 6000 295440
rect 578000 295344 582820 295440
rect 3326 295060 3332 295112
rect 3384 295100 3390 295112
rect 6546 295100 6552 295112
rect 3384 295072 6552 295100
rect 3384 295060 3390 295072
rect 6546 295060 6552 295072
rect 6604 295060 6610 295112
rect 1104 294800 6000 294896
rect 578000 294800 582820 294896
rect 1104 294256 6000 294352
rect 578000 294256 582820 294352
rect 1104 293712 6000 293808
rect 578000 293712 582820 293808
rect 1104 293168 6000 293264
rect 578000 293168 582820 293264
rect 1104 292624 6000 292720
rect 578000 292624 582820 292720
rect 1104 292080 6000 292176
rect 578000 292080 582820 292176
rect 1104 291536 6000 291632
rect 578000 291536 582820 291632
rect 1104 290992 6000 291088
rect 578000 290992 582820 291088
rect 1104 290448 6000 290544
rect 578000 290448 582820 290544
rect 1104 289904 6000 290000
rect 578000 289904 582820 290000
rect 1104 289360 6000 289456
rect 578000 289360 582820 289456
rect 1104 288816 6000 288912
rect 578000 288816 582820 288912
rect 1104 288272 6000 288368
rect 578000 288272 582820 288368
rect 1104 287728 6000 287824
rect 578000 287728 582820 287824
rect 1104 287184 6000 287280
rect 578000 287184 582820 287280
rect 1104 286640 6000 286736
rect 578000 286640 582820 286736
rect 1104 286096 6000 286192
rect 578000 286096 582820 286192
rect 1104 285552 6000 285648
rect 578000 285552 582820 285648
rect 1104 285008 6000 285104
rect 578000 285008 582820 285104
rect 1104 284464 6000 284560
rect 578000 284464 582820 284560
rect 1104 283920 6000 284016
rect 578000 283920 582820 284016
rect 1104 283376 6000 283472
rect 578000 283376 582820 283472
rect 1104 282832 6000 282928
rect 578000 282832 582820 282928
rect 1104 282288 6000 282384
rect 578000 282288 582820 282384
rect 1104 281744 6000 281840
rect 578000 281744 582820 281840
rect 1104 281200 6000 281296
rect 578000 281200 582820 281296
rect 1104 280656 6000 280752
rect 578000 280656 582820 280752
rect 1104 280112 6000 280208
rect 578000 280112 582820 280208
rect 2774 280032 2780 280084
rect 2832 280072 2838 280084
rect 5074 280072 5080 280084
rect 2832 280044 5080 280072
rect 2832 280032 2838 280044
rect 5074 280032 5080 280044
rect 5132 280032 5138 280084
rect 1104 279568 6000 279664
rect 578000 279568 582820 279664
rect 1104 279024 6000 279120
rect 578000 279024 582820 279120
rect 1104 278480 6000 278576
rect 578000 278480 582820 278576
rect 1104 277936 6000 278032
rect 578000 277936 582820 278032
rect 1104 277392 6000 277488
rect 578000 277392 582820 277488
rect 1104 276848 6000 276944
rect 578000 276848 582820 276944
rect 1104 276304 6000 276400
rect 578000 276304 582820 276400
rect 1104 275760 6000 275856
rect 578000 275760 582820 275856
rect 1104 275216 6000 275312
rect 578000 275216 582820 275312
rect 1104 274672 6000 274768
rect 578000 274672 582820 274768
rect 1104 274128 6000 274224
rect 578000 274128 582820 274224
rect 1104 273584 6000 273680
rect 578000 273584 582820 273680
rect 1104 273040 6000 273136
rect 578000 273040 582820 273136
rect 1104 272496 6000 272592
rect 578000 272496 582820 272592
rect 1104 271952 6000 272048
rect 578000 271952 582820 272048
rect 1104 271408 6000 271504
rect 578000 271408 582820 271504
rect 1104 270864 6000 270960
rect 578000 270864 582820 270960
rect 1104 270320 6000 270416
rect 578000 270320 582820 270416
rect 1104 269776 6000 269872
rect 578000 269776 582820 269872
rect 1104 269232 6000 269328
rect 578000 269232 582820 269328
rect 1104 268688 6000 268784
rect 578000 268688 582820 268784
rect 1104 268144 6000 268240
rect 578000 268144 582820 268240
rect 1104 267600 6000 267696
rect 578000 267600 582820 267696
rect 1104 267056 6000 267152
rect 578000 267056 582820 267152
rect 1104 266512 6000 266608
rect 578000 266512 582820 266608
rect 3142 266228 3148 266280
rect 3200 266268 3206 266280
rect 6454 266268 6460 266280
rect 3200 266240 6460 266268
rect 3200 266228 3206 266240
rect 6454 266228 6460 266240
rect 6512 266228 6518 266280
rect 1104 265968 6000 266064
rect 578000 265968 582820 266064
rect 1104 265424 6000 265520
rect 578000 265424 582820 265520
rect 1104 264880 6000 264976
rect 578000 264880 582820 264976
rect 576394 264800 576400 264852
rect 576452 264840 576458 264852
rect 580166 264840 580172 264852
rect 576452 264812 580172 264840
rect 576452 264800 576458 264812
rect 580166 264800 580172 264812
rect 580224 264800 580230 264852
rect 1104 264336 6000 264432
rect 578000 264336 582820 264432
rect 1104 263792 6000 263888
rect 578000 263792 582820 263888
rect 1104 263248 6000 263344
rect 578000 263248 582820 263344
rect 1104 262704 6000 262800
rect 578000 262704 582820 262800
rect 1104 262160 6000 262256
rect 578000 262160 582820 262256
rect 1104 261616 6000 261712
rect 578000 261616 582820 261712
rect 1104 261072 6000 261168
rect 578000 261072 582820 261168
rect 1104 260528 6000 260624
rect 578000 260528 582820 260624
rect 1104 259984 6000 260080
rect 578000 259984 582820 260080
rect 1104 259440 6000 259536
rect 578000 259440 582820 259536
rect 1104 258896 6000 258992
rect 578000 258896 582820 258992
rect 1104 258352 6000 258448
rect 578000 258352 582820 258448
rect 1104 257808 6000 257904
rect 578000 257808 582820 257904
rect 1104 257264 6000 257360
rect 578000 257264 582820 257360
rect 1104 256720 6000 256816
rect 578000 256720 582820 256816
rect 1104 256176 6000 256272
rect 578000 256176 582820 256272
rect 1104 255632 6000 255728
rect 578000 255632 582820 255728
rect 1104 255088 6000 255184
rect 578000 255088 582820 255184
rect 1104 254544 6000 254640
rect 578000 254544 582820 254640
rect 1104 254000 6000 254096
rect 578000 254000 582820 254096
rect 1104 253456 6000 253552
rect 578000 253456 582820 253552
rect 1104 252912 6000 253008
rect 578000 252912 582820 253008
rect 3234 252492 3240 252544
rect 3292 252532 3298 252544
rect 6362 252532 6368 252544
rect 3292 252504 6368 252532
rect 3292 252492 3298 252504
rect 6362 252492 6368 252504
rect 6420 252492 6426 252544
rect 575198 252492 575204 252544
rect 575256 252532 575262 252544
rect 580166 252532 580172 252544
rect 575256 252504 580172 252532
rect 575256 252492 575262 252504
rect 580166 252492 580172 252504
rect 580224 252492 580230 252544
rect 1104 252368 6000 252464
rect 578000 252368 582820 252464
rect 1104 251824 6000 251920
rect 578000 251824 582820 251920
rect 1104 251280 6000 251376
rect 578000 251280 582820 251376
rect 1104 250736 6000 250832
rect 578000 250736 582820 250832
rect 1104 250192 6000 250288
rect 578000 250192 582820 250288
rect 1104 249648 6000 249744
rect 578000 249648 582820 249744
rect 1104 249104 6000 249200
rect 578000 249104 582820 249200
rect 1104 248560 6000 248656
rect 578000 248560 582820 248656
rect 1104 248016 6000 248112
rect 578000 248016 582820 248112
rect 1104 247472 6000 247568
rect 578000 247472 582820 247568
rect 1104 246928 6000 247024
rect 578000 246928 582820 247024
rect 1104 246384 6000 246480
rect 578000 246384 582820 246480
rect 1104 245840 6000 245936
rect 578000 245840 582820 245936
rect 1104 245296 6000 245392
rect 578000 245296 582820 245392
rect 1104 244752 6000 244848
rect 578000 244752 582820 244848
rect 1104 244208 6000 244304
rect 578000 244208 582820 244304
rect 1104 243664 6000 243760
rect 578000 243664 582820 243760
rect 1104 243120 6000 243216
rect 578000 243120 582820 243216
rect 1104 242576 6000 242672
rect 578000 242576 582820 242672
rect 1104 242032 6000 242128
rect 578000 242032 582820 242128
rect 1104 241488 6000 241584
rect 578000 241488 582820 241584
rect 1104 240944 6000 241040
rect 578000 240944 582820 241040
rect 1104 240400 6000 240496
rect 578000 240400 582820 240496
rect 1104 239856 6000 239952
rect 578000 239856 582820 239952
rect 1104 239312 6000 239408
rect 578000 239312 582820 239408
rect 1104 238768 6000 238864
rect 578000 238768 582820 238864
rect 1104 238224 6000 238320
rect 578000 238224 582820 238320
rect 1104 237680 6000 237776
rect 578000 237680 582820 237776
rect 1104 237136 6000 237232
rect 578000 237136 582820 237232
rect 1104 236592 6000 236688
rect 578000 236592 582820 236688
rect 1104 236048 6000 236144
rect 578000 236048 582820 236144
rect 1104 235504 6000 235600
rect 578000 235504 582820 235600
rect 1104 234960 6000 235056
rect 578000 234960 582820 235056
rect 1104 234416 6000 234512
rect 578000 234416 582820 234512
rect 1104 233872 6000 233968
rect 578000 233872 582820 233968
rect 1104 233328 6000 233424
rect 578000 233328 582820 233424
rect 1104 232784 6000 232880
rect 578000 232784 582820 232880
rect 1104 232240 6000 232336
rect 578000 232240 582820 232336
rect 1104 231696 6000 231792
rect 578000 231696 582820 231792
rect 1104 231152 6000 231248
rect 578000 231152 582820 231248
rect 1104 230608 6000 230704
rect 578000 230608 582820 230704
rect 1104 230064 6000 230160
rect 578000 230064 582820 230160
rect 1104 229520 6000 229616
rect 578000 229520 582820 229616
rect 1104 228976 6000 229072
rect 578000 228976 582820 229072
rect 1104 228432 6000 228528
rect 578000 228432 582820 228528
rect 1104 227888 6000 227984
rect 578000 227888 582820 227984
rect 1104 227344 6000 227440
rect 578000 227344 582820 227440
rect 1104 226800 6000 226896
rect 578000 226800 582820 226896
rect 1104 226256 6000 226352
rect 578000 226256 582820 226352
rect 1104 225712 6000 225808
rect 578000 225712 582820 225808
rect 1104 225168 6000 225264
rect 578000 225168 582820 225264
rect 1104 224624 6000 224720
rect 578000 224624 582820 224720
rect 1104 224080 6000 224176
rect 578000 224080 582820 224176
rect 1104 223536 6000 223632
rect 578000 223536 582820 223632
rect 1104 222992 6000 223088
rect 578000 222992 582820 223088
rect 1104 222448 6000 222544
rect 578000 222448 582820 222544
rect 1104 221904 6000 222000
rect 578000 221904 582820 222000
rect 1104 221360 6000 221456
rect 578000 221360 582820 221456
rect 1104 220816 6000 220912
rect 578000 220816 582820 220912
rect 1104 220272 6000 220368
rect 578000 220272 582820 220368
rect 1104 219728 6000 219824
rect 578000 219728 582820 219824
rect 1104 219184 6000 219280
rect 578000 219184 582820 219280
rect 1104 218640 6000 218736
rect 578000 218640 582820 218736
rect 1104 218096 6000 218192
rect 578000 218096 582820 218192
rect 1104 217552 6000 217648
rect 578000 217552 582820 217648
rect 1104 217008 6000 217104
rect 578000 217008 582820 217104
rect 1104 216464 6000 216560
rect 578000 216464 582820 216560
rect 1104 215920 6000 216016
rect 578000 215920 582820 216016
rect 1104 215376 6000 215472
rect 578000 215376 582820 215472
rect 1104 214832 6000 214928
rect 578000 214832 582820 214928
rect 1104 214288 6000 214384
rect 578000 214288 582820 214384
rect 1104 213744 6000 213840
rect 578000 213744 582820 213840
rect 1104 213200 6000 213296
rect 578000 213200 582820 213296
rect 1104 212656 6000 212752
rect 578000 212656 582820 212752
rect 1104 212112 6000 212208
rect 578000 212112 582820 212208
rect 1104 211568 6000 211664
rect 578000 211568 582820 211664
rect 1104 211024 6000 211120
rect 578000 211024 582820 211120
rect 1104 210480 6000 210576
rect 578000 210480 582820 210576
rect 1104 209936 6000 210032
rect 578000 209936 582820 210032
rect 1104 209392 6000 209488
rect 578000 209392 582820 209488
rect 1104 208848 6000 208944
rect 578000 208848 582820 208944
rect 1104 208304 6000 208400
rect 578000 208304 582820 208400
rect 3142 208156 3148 208208
rect 3200 208196 3206 208208
rect 6270 208196 6276 208208
rect 3200 208168 6276 208196
rect 3200 208156 3206 208168
rect 6270 208156 6276 208168
rect 6328 208156 6334 208208
rect 1104 207760 6000 207856
rect 578000 207760 582820 207856
rect 1104 207216 6000 207312
rect 578000 207216 582820 207312
rect 1104 206672 6000 206768
rect 578000 206672 582820 206768
rect 1104 206128 6000 206224
rect 578000 206128 582820 206224
rect 1104 205584 6000 205680
rect 578000 205584 582820 205680
rect 575106 205504 575112 205556
rect 575164 205544 575170 205556
rect 580166 205544 580172 205556
rect 575164 205516 580172 205544
rect 575164 205504 575170 205516
rect 580166 205504 580172 205516
rect 580224 205504 580230 205556
rect 1104 205040 6000 205136
rect 578000 205040 582820 205136
rect 1104 204496 6000 204592
rect 578000 204496 582820 204592
rect 1104 203952 6000 204048
rect 578000 203952 582820 204048
rect 1104 203408 6000 203504
rect 578000 203408 582820 203504
rect 1104 202864 6000 202960
rect 578000 202864 582820 202960
rect 1104 202320 6000 202416
rect 578000 202320 582820 202416
rect 1104 201776 6000 201872
rect 578000 201776 582820 201872
rect 1104 201232 6000 201328
rect 578000 201232 582820 201328
rect 1104 200688 6000 200784
rect 578000 200688 582820 200784
rect 1104 200144 6000 200240
rect 578000 200144 582820 200240
rect 1104 199600 6000 199696
rect 578000 199600 582820 199696
rect 1104 199056 6000 199152
rect 578000 199056 582820 199152
rect 1104 198512 6000 198608
rect 578000 198512 582820 198608
rect 1104 197968 6000 198064
rect 578000 197968 582820 198064
rect 1104 197424 6000 197520
rect 578000 197424 582820 197520
rect 1104 196880 6000 196976
rect 578000 196880 582820 196976
rect 1104 196336 6000 196432
rect 578000 196336 582820 196432
rect 1104 195792 6000 195888
rect 578000 195792 582820 195888
rect 1104 195248 6000 195344
rect 578000 195248 582820 195344
rect 1104 194704 6000 194800
rect 578000 194704 582820 194800
rect 2774 194420 2780 194472
rect 2832 194460 2838 194472
rect 4982 194460 4988 194472
rect 2832 194432 4988 194460
rect 2832 194420 2838 194432
rect 4982 194420 4988 194432
rect 5040 194420 5046 194472
rect 1104 194160 6000 194256
rect 578000 194160 582820 194256
rect 1104 193616 6000 193712
rect 578000 193616 582820 193712
rect 1104 193072 6000 193168
rect 578000 193072 582820 193168
rect 1104 192528 6000 192624
rect 578000 192528 582820 192624
rect 1104 191984 6000 192080
rect 578000 191984 582820 192080
rect 1104 191440 6000 191536
rect 578000 191440 582820 191536
rect 1104 190896 6000 190992
rect 578000 190896 582820 190992
rect 1104 190352 6000 190448
rect 578000 190352 582820 190448
rect 1104 189808 6000 189904
rect 578000 189808 582820 189904
rect 1104 189264 6000 189360
rect 578000 189264 582820 189360
rect 1104 188720 6000 188816
rect 578000 188720 582820 188816
rect 1104 188176 6000 188272
rect 578000 188176 582820 188272
rect 1104 187632 6000 187728
rect 578000 187632 582820 187728
rect 1104 187088 6000 187184
rect 578000 187088 582820 187184
rect 1104 186544 6000 186640
rect 578000 186544 582820 186640
rect 1104 186000 6000 186096
rect 578000 186000 582820 186096
rect 1104 185456 6000 185552
rect 578000 185456 582820 185552
rect 1104 184912 6000 185008
rect 578000 184912 582820 185008
rect 1104 184368 6000 184464
rect 578000 184368 582820 184464
rect 1104 183824 6000 183920
rect 578000 183824 582820 183920
rect 1104 183280 6000 183376
rect 578000 183280 582820 183376
rect 1104 182736 6000 182832
rect 578000 182736 582820 182832
rect 1104 182192 6000 182288
rect 578000 182192 582820 182288
rect 575014 182112 575020 182164
rect 575072 182152 575078 182164
rect 580166 182152 580172 182164
rect 575072 182124 580172 182152
rect 575072 182112 575078 182124
rect 580166 182112 580172 182124
rect 580224 182112 580230 182164
rect 1104 181648 6000 181744
rect 578000 181648 582820 181744
rect 1104 181104 6000 181200
rect 578000 181104 582820 181200
rect 1104 180560 6000 180656
rect 578000 180560 582820 180656
rect 1104 180016 6000 180112
rect 578000 180016 582820 180112
rect 1104 179472 6000 179568
rect 578000 179472 582820 179568
rect 1104 178928 6000 179024
rect 578000 178928 582820 179024
rect 1104 178384 6000 178480
rect 578000 178384 582820 178480
rect 1104 177840 6000 177936
rect 578000 177840 582820 177936
rect 1104 177296 6000 177392
rect 578000 177296 582820 177392
rect 1104 176752 6000 176848
rect 578000 176752 582820 176848
rect 1104 176208 6000 176304
rect 578000 176208 582820 176304
rect 1104 175664 6000 175760
rect 578000 175664 582820 175760
rect 1104 175120 6000 175216
rect 578000 175120 582820 175216
rect 1104 174576 6000 174672
rect 578000 174576 582820 174672
rect 1104 174032 6000 174128
rect 578000 174032 582820 174128
rect 1104 173488 6000 173584
rect 578000 173488 582820 173584
rect 1104 172944 6000 173040
rect 578000 172944 582820 173040
rect 1104 172400 6000 172496
rect 578000 172400 582820 172496
rect 1104 171856 6000 171952
rect 578000 171856 582820 171952
rect 1104 171312 6000 171408
rect 578000 171312 582820 171408
rect 576302 171028 576308 171080
rect 576360 171068 576366 171080
rect 579614 171068 579620 171080
rect 576360 171040 579620 171068
rect 576360 171028 576366 171040
rect 579614 171028 579620 171040
rect 579672 171028 579678 171080
rect 1104 170768 6000 170864
rect 578000 170768 582820 170864
rect 1104 170224 6000 170320
rect 578000 170224 582820 170320
rect 1104 169680 6000 169776
rect 578000 169680 582820 169776
rect 1104 169136 6000 169232
rect 578000 169136 582820 169232
rect 1104 168592 6000 168688
rect 578000 168592 582820 168688
rect 1104 168048 6000 168144
rect 578000 168048 582820 168144
rect 1104 167504 6000 167600
rect 578000 167504 582820 167600
rect 1104 166960 6000 167056
rect 578000 166960 582820 167056
rect 1104 166416 6000 166512
rect 578000 166416 582820 166512
rect 1104 165872 6000 165968
rect 578000 165872 582820 165968
rect 1118 165656 1124 165708
rect 1176 165696 1182 165708
rect 7926 165696 7932 165708
rect 1176 165668 7932 165696
rect 1176 165656 1182 165668
rect 7926 165656 7932 165668
rect 7984 165656 7990 165708
rect 1104 165328 6000 165424
rect 578000 165328 582820 165424
rect 1104 164784 6000 164880
rect 578000 164784 582820 164880
rect 1104 164240 6000 164336
rect 578000 164240 582820 164336
rect 1104 163696 6000 163792
rect 578000 163696 582820 163792
rect 1104 163152 6000 163248
rect 578000 163152 582820 163248
rect 1104 162608 6000 162704
rect 578000 162608 582820 162704
rect 1104 162064 6000 162160
rect 578000 162064 582820 162160
rect 1104 161520 6000 161616
rect 578000 161520 582820 161616
rect 1104 160976 6000 161072
rect 578000 160976 582820 161072
rect 1104 160432 6000 160528
rect 578000 160432 582820 160528
rect 1104 159888 6000 159984
rect 578000 159888 582820 159984
rect 1104 159344 6000 159440
rect 578000 159344 582820 159440
rect 1104 158800 6000 158896
rect 578000 158800 582820 158896
rect 577498 158652 577504 158704
rect 577556 158692 577562 158704
rect 580626 158692 580632 158704
rect 577556 158664 580632 158692
rect 577556 158652 577562 158664
rect 580626 158652 580632 158664
rect 580684 158652 580690 158704
rect 1104 158256 6000 158352
rect 578000 158256 582820 158352
rect 1104 157712 6000 157808
rect 578000 157712 582820 157808
rect 1104 157168 6000 157264
rect 578000 157168 582820 157264
rect 1104 156624 6000 156720
rect 578000 156624 582820 156720
rect 1104 156080 6000 156176
rect 578000 156080 582820 156176
rect 1104 155536 6000 155632
rect 578000 155536 582820 155632
rect 1104 154992 6000 155088
rect 578000 154992 582820 155088
rect 1104 154448 6000 154544
rect 578000 154448 582820 154544
rect 1104 153904 6000 154000
rect 578000 153904 582820 154000
rect 1104 153360 6000 153456
rect 578000 153360 582820 153456
rect 1104 152816 6000 152912
rect 578000 152816 582820 152912
rect 1104 152272 6000 152368
rect 578000 152272 582820 152368
rect 1104 151728 6000 151824
rect 578000 151728 582820 151824
rect 1104 151184 6000 151280
rect 578000 151184 582820 151280
rect 2774 150832 2780 150884
rect 2832 150872 2838 150884
rect 4890 150872 4896 150884
rect 2832 150844 4896 150872
rect 2832 150832 2838 150844
rect 4890 150832 4896 150844
rect 4948 150832 4954 150884
rect 1104 150640 6000 150736
rect 578000 150640 582820 150736
rect 1104 150096 6000 150192
rect 578000 150096 582820 150192
rect 1104 149552 6000 149648
rect 578000 149552 582820 149648
rect 1104 149008 6000 149104
rect 578000 149008 582820 149104
rect 1104 148464 6000 148560
rect 578000 148464 582820 148560
rect 1104 147920 6000 148016
rect 578000 147920 582820 148016
rect 1104 147376 6000 147472
rect 578000 147376 582820 147472
rect 1104 146832 6000 146928
rect 578000 146832 582820 146928
rect 1104 146288 6000 146384
rect 578000 146288 582820 146384
rect 1104 145744 6000 145840
rect 578000 145744 582820 145840
rect 1104 145200 6000 145296
rect 578000 145200 582820 145296
rect 1104 144656 6000 144752
rect 578000 144656 582820 144752
rect 1104 144112 6000 144208
rect 578000 144112 582820 144208
rect 1104 143568 6000 143664
rect 578000 143568 582820 143664
rect 1104 143024 6000 143120
rect 578000 143024 582820 143120
rect 1104 142480 6000 142576
rect 578000 142480 582820 142576
rect 1104 141936 6000 142032
rect 578000 141936 582820 142032
rect 1104 141392 6000 141488
rect 578000 141392 582820 141488
rect 1104 140848 6000 140944
rect 578000 140848 582820 140944
rect 1104 140304 6000 140400
rect 578000 140304 582820 140400
rect 1104 139760 6000 139856
rect 578000 139760 582820 139856
rect 1104 139216 6000 139312
rect 578000 139216 582820 139312
rect 1104 138672 6000 138768
rect 578000 138672 582820 138768
rect 1104 138128 6000 138224
rect 578000 138128 582820 138224
rect 1104 137584 6000 137680
rect 578000 137584 582820 137680
rect 1104 137040 6000 137136
rect 578000 137040 582820 137136
rect 1104 136496 6000 136592
rect 578000 136496 582820 136592
rect 3326 136348 3332 136400
rect 3384 136388 3390 136400
rect 7834 136388 7840 136400
rect 3384 136360 7840 136388
rect 3384 136348 3390 136360
rect 7834 136348 7840 136360
rect 7892 136348 7898 136400
rect 1104 135952 6000 136048
rect 578000 135952 582820 136048
rect 1104 135408 6000 135504
rect 578000 135408 582820 135504
rect 1104 134864 6000 134960
rect 578000 134864 582820 134960
rect 1104 134320 6000 134416
rect 578000 134320 582820 134416
rect 1104 133776 6000 133872
rect 578000 133776 582820 133872
rect 1104 133232 6000 133328
rect 578000 133232 582820 133328
rect 1104 132688 6000 132784
rect 578000 132688 582820 132784
rect 1104 132144 6000 132240
rect 578000 132144 582820 132240
rect 1104 131600 6000 131696
rect 578000 131600 582820 131696
rect 1104 131056 6000 131152
rect 578000 131056 582820 131152
rect 1104 130512 6000 130608
rect 578000 130512 582820 130608
rect 1104 129968 6000 130064
rect 578000 129968 582820 130064
rect 1104 129424 6000 129520
rect 578000 129424 582820 129520
rect 1104 128880 6000 128976
rect 578000 128880 582820 128976
rect 1104 128336 6000 128432
rect 578000 128336 582820 128432
rect 1104 127792 6000 127888
rect 578000 127792 582820 127888
rect 1104 127248 6000 127344
rect 578000 127248 582820 127344
rect 1104 126704 6000 126800
rect 578000 126704 582820 126800
rect 1104 126160 6000 126256
rect 578000 126160 582820 126256
rect 1104 125616 6000 125712
rect 578000 125616 582820 125712
rect 1104 125072 6000 125168
rect 578000 125072 582820 125168
rect 1104 124528 6000 124624
rect 578000 124528 582820 124624
rect 1104 123984 6000 124080
rect 578000 123984 582820 124080
rect 1104 123440 6000 123536
rect 578000 123440 582820 123536
rect 1104 122896 6000 122992
rect 578000 122896 582820 122992
rect 1104 122352 6000 122448
rect 578000 122352 582820 122448
rect 3326 122068 3332 122120
rect 3384 122108 3390 122120
rect 7742 122108 7748 122120
rect 3384 122080 7748 122108
rect 3384 122068 3390 122080
rect 7742 122068 7748 122080
rect 7800 122068 7806 122120
rect 1104 121808 6000 121904
rect 578000 121808 582820 121904
rect 1104 121264 6000 121360
rect 578000 121264 582820 121360
rect 1104 120720 6000 120816
rect 578000 120720 582820 120816
rect 1104 120176 6000 120272
rect 578000 120176 582820 120272
rect 1104 119632 6000 119728
rect 578000 119632 582820 119728
rect 1104 119088 6000 119184
rect 578000 119088 582820 119184
rect 1104 118544 6000 118640
rect 578000 118544 582820 118640
rect 1104 118000 6000 118096
rect 578000 118000 582820 118096
rect 1104 117456 6000 117552
rect 578000 117456 582820 117552
rect 1104 116912 6000 117008
rect 578000 116912 582820 117008
rect 1104 116368 6000 116464
rect 578000 116368 582820 116464
rect 1104 115824 6000 115920
rect 578000 115824 582820 115920
rect 1104 115280 6000 115376
rect 578000 115280 582820 115376
rect 1104 114736 6000 114832
rect 578000 114736 582820 114832
rect 1104 114192 6000 114288
rect 578000 114192 582820 114288
rect 1104 113648 6000 113744
rect 578000 113648 582820 113744
rect 1104 113104 6000 113200
rect 578000 113104 582820 113200
rect 1104 112560 6000 112656
rect 578000 112560 582820 112656
rect 1104 112016 6000 112112
rect 578000 112016 582820 112112
rect 574922 111732 574928 111784
rect 574980 111772 574986 111784
rect 579614 111772 579620 111784
rect 574980 111744 579620 111772
rect 574980 111732 574986 111744
rect 579614 111732 579620 111744
rect 579672 111732 579678 111784
rect 1104 111472 6000 111568
rect 578000 111472 582820 111568
rect 1104 110928 6000 111024
rect 578000 110928 582820 111024
rect 1104 110384 6000 110480
rect 578000 110384 582820 110480
rect 1104 109840 6000 109936
rect 578000 109840 582820 109936
rect 1104 109296 6000 109392
rect 578000 109296 582820 109392
rect 1104 108752 6000 108848
rect 578000 108752 582820 108848
rect 1104 108208 6000 108304
rect 578000 108208 582820 108304
rect 1104 107664 6000 107760
rect 578000 107664 582820 107760
rect 1104 107120 6000 107216
rect 578000 107120 582820 107216
rect 1104 106576 6000 106672
rect 578000 106576 582820 106672
rect 1104 106032 6000 106128
rect 578000 106032 582820 106128
rect 1104 105488 6000 105584
rect 578000 105488 582820 105584
rect 1104 104944 6000 105040
rect 578000 104944 582820 105040
rect 1104 104400 6000 104496
rect 578000 104400 582820 104496
rect 1104 103856 6000 103952
rect 578000 103856 582820 103952
rect 1104 103312 6000 103408
rect 578000 103312 582820 103408
rect 1104 102768 6000 102864
rect 578000 102768 582820 102864
rect 1104 102224 6000 102320
rect 578000 102224 582820 102320
rect 1104 101680 6000 101776
rect 578000 101680 582820 101776
rect 1104 101136 6000 101232
rect 578000 101136 582820 101232
rect 1104 100592 6000 100688
rect 578000 100592 582820 100688
rect 1104 100048 6000 100144
rect 578000 100048 582820 100144
rect 1104 99504 6000 99600
rect 578000 99504 582820 99600
rect 1104 98960 6000 99056
rect 578000 98960 582820 99056
rect 1104 98416 6000 98512
rect 578000 98416 582820 98512
rect 1104 97872 6000 97968
rect 578000 97872 582820 97968
rect 1104 97328 6000 97424
rect 578000 97328 582820 97424
rect 1104 96784 6000 96880
rect 578000 96784 582820 96880
rect 1104 96240 6000 96336
rect 578000 96240 582820 96336
rect 1104 95696 6000 95792
rect 578000 95696 582820 95792
rect 1104 95152 6000 95248
rect 578000 95152 582820 95248
rect 1104 94608 6000 94704
rect 578000 94608 582820 94704
rect 1104 94064 6000 94160
rect 578000 94064 582820 94160
rect 1104 93520 6000 93616
rect 578000 93520 582820 93616
rect 1104 92976 6000 93072
rect 578000 92976 582820 93072
rect 1104 92432 6000 92528
rect 578000 92432 582820 92528
rect 1104 91888 6000 91984
rect 578000 91888 582820 91984
rect 1104 91344 6000 91440
rect 578000 91344 582820 91440
rect 1104 90800 6000 90896
rect 578000 90800 582820 90896
rect 1104 90256 6000 90352
rect 578000 90256 582820 90352
rect 1104 89712 6000 89808
rect 578000 89712 582820 89808
rect 1104 89168 6000 89264
rect 578000 89168 582820 89264
rect 1104 88624 6000 88720
rect 578000 88624 582820 88720
rect 1104 88080 6000 88176
rect 578000 88080 582820 88176
rect 1104 87536 6000 87632
rect 578000 87536 582820 87632
rect 1104 86992 6000 87088
rect 578000 86992 582820 87088
rect 1104 86448 6000 86544
rect 578000 86448 582820 86544
rect 1104 85904 6000 86000
rect 578000 85904 582820 86000
rect 1104 85360 6000 85456
rect 578000 85360 582820 85456
rect 1104 84816 6000 84912
rect 578000 84816 582820 84912
rect 1104 84272 6000 84368
rect 578000 84272 582820 84368
rect 1104 83728 6000 83824
rect 578000 83728 582820 83824
rect 1104 83184 6000 83280
rect 578000 83184 582820 83280
rect 1104 82640 6000 82736
rect 578000 82640 582820 82736
rect 1104 82096 6000 82192
rect 578000 82096 582820 82192
rect 1104 81552 6000 81648
rect 578000 81552 582820 81648
rect 1104 81008 6000 81104
rect 578000 81008 582820 81104
rect 1104 80464 6000 80560
rect 578000 80464 582820 80560
rect 1104 79920 6000 80016
rect 578000 79920 582820 80016
rect 3050 79840 3056 79892
rect 3108 79880 3114 79892
rect 7650 79880 7656 79892
rect 3108 79852 7656 79880
rect 3108 79840 3114 79852
rect 7650 79840 7656 79852
rect 7708 79840 7714 79892
rect 1104 79376 6000 79472
rect 578000 79376 582820 79472
rect 1104 78832 6000 78928
rect 578000 78832 582820 78928
rect 1104 78288 6000 78384
rect 578000 78288 582820 78384
rect 1104 77744 6000 77840
rect 578000 77744 582820 77840
rect 1104 77200 6000 77296
rect 578000 77200 582820 77296
rect 1104 76656 6000 76752
rect 578000 76656 582820 76752
rect 1104 76112 6000 76208
rect 578000 76112 582820 76208
rect 1104 75568 6000 75664
rect 578000 75568 582820 75664
rect 1104 75024 6000 75120
rect 578000 75024 582820 75120
rect 1104 74480 6000 74576
rect 578000 74480 582820 74576
rect 1104 73936 6000 74032
rect 578000 73936 582820 74032
rect 1104 73392 6000 73488
rect 578000 73392 582820 73488
rect 1104 72848 6000 72944
rect 578000 72848 582820 72944
rect 1104 72304 6000 72400
rect 578000 72304 582820 72400
rect 1104 71760 6000 71856
rect 578000 71760 582820 71856
rect 1104 71216 6000 71312
rect 578000 71216 582820 71312
rect 1104 70672 6000 70768
rect 578000 70672 582820 70768
rect 1104 70128 6000 70224
rect 578000 70128 582820 70224
rect 1104 69584 6000 69680
rect 578000 69584 582820 69680
rect 1104 69040 6000 69136
rect 578000 69040 582820 69136
rect 1104 68496 6000 68592
rect 578000 68496 582820 68592
rect 1104 67952 6000 68048
rect 578000 67952 582820 68048
rect 1104 67408 6000 67504
rect 578000 67408 582820 67504
rect 1104 66864 6000 66960
rect 578000 66864 582820 66960
rect 1104 66320 6000 66416
rect 578000 66320 582820 66416
rect 1104 65776 6000 65872
rect 578000 65776 582820 65872
rect 1104 65232 6000 65328
rect 578000 65232 582820 65328
rect 576210 64812 576216 64864
rect 576268 64852 576274 64864
rect 579798 64852 579804 64864
rect 576268 64824 579804 64852
rect 576268 64812 576274 64824
rect 579798 64812 579804 64824
rect 579856 64812 579862 64864
rect 1104 64688 6000 64784
rect 578000 64688 582820 64784
rect 2774 64540 2780 64592
rect 2832 64580 2838 64592
rect 4798 64580 4804 64592
rect 2832 64552 4804 64580
rect 2832 64540 2838 64552
rect 4798 64540 4804 64552
rect 4856 64540 4862 64592
rect 1104 64144 6000 64240
rect 578000 64144 582820 64240
rect 1104 63600 6000 63696
rect 578000 63600 582820 63696
rect 1104 63056 6000 63152
rect 578000 63056 582820 63152
rect 1104 62512 6000 62608
rect 578000 62512 582820 62608
rect 1104 61968 6000 62064
rect 578000 61968 582820 62064
rect 1104 61424 6000 61520
rect 578000 61424 582820 61520
rect 1104 60880 6000 60976
rect 578000 60880 582820 60976
rect 1104 60336 6000 60432
rect 578000 60336 582820 60432
rect 1104 59792 6000 59888
rect 578000 59792 582820 59888
rect 1104 59248 6000 59344
rect 578000 59248 582820 59344
rect 1104 58704 6000 58800
rect 578000 58704 582820 58800
rect 1104 58160 6000 58256
rect 578000 58160 582820 58256
rect 1104 57616 6000 57712
rect 578000 57616 582820 57712
rect 1104 57072 6000 57168
rect 578000 57072 582820 57168
rect 1104 56528 6000 56624
rect 578000 56528 582820 56624
rect 1104 55984 6000 56080
rect 578000 55984 582820 56080
rect 1104 55440 6000 55536
rect 578000 55440 582820 55536
rect 1104 54896 6000 54992
rect 578000 54896 582820 54992
rect 1104 54352 6000 54448
rect 578000 54352 582820 54448
rect 1104 53808 6000 53904
rect 578000 53808 582820 53904
rect 1104 53264 6000 53360
rect 578000 53264 582820 53360
rect 1104 52720 6000 52816
rect 578000 52720 582820 52816
rect 1104 52176 6000 52272
rect 578000 52176 582820 52272
rect 1104 51632 6000 51728
rect 578000 51632 582820 51728
rect 1104 51088 6000 51184
rect 578000 51088 582820 51184
rect 1104 50544 6000 50640
rect 578000 50544 582820 50640
rect 1104 50000 6000 50096
rect 578000 50000 582820 50096
rect 1104 49456 6000 49552
rect 578000 49456 582820 49552
rect 1104 48912 6000 49008
rect 578000 48912 582820 49008
rect 1104 48368 6000 48464
rect 578000 48368 582820 48464
rect 1104 47824 6000 47920
rect 578000 47824 582820 47920
rect 1104 47280 6000 47376
rect 578000 47280 582820 47376
rect 1104 46736 6000 46832
rect 578000 46736 582820 46832
rect 1104 46192 6000 46288
rect 578000 46192 582820 46288
rect 1104 45648 6000 45744
rect 578000 45648 582820 45744
rect 1104 45104 6000 45200
rect 578000 45104 582820 45200
rect 1104 44560 6000 44656
rect 578000 44560 582820 44656
rect 1104 44016 6000 44112
rect 578000 44016 582820 44112
rect 1104 43472 6000 43568
rect 578000 43472 582820 43568
rect 1104 42928 6000 43024
rect 578000 42928 582820 43024
rect 1104 42384 6000 42480
rect 578000 42384 582820 42480
rect 1104 41840 6000 41936
rect 578000 41840 582820 41936
rect 1104 41296 6000 41392
rect 578000 41296 582820 41392
rect 575014 41216 575020 41268
rect 575072 41256 575078 41268
rect 580166 41256 580172 41268
rect 575072 41228 580172 41256
rect 575072 41216 575078 41228
rect 580166 41216 580172 41228
rect 580224 41216 580230 41268
rect 1104 40752 6000 40848
rect 578000 40752 582820 40848
rect 1104 40208 6000 40304
rect 578000 40208 582820 40304
rect 1104 39664 6000 39760
rect 578000 39664 582820 39760
rect 1104 39120 6000 39216
rect 578000 39120 582820 39216
rect 1104 38576 6000 38672
rect 578000 38576 582820 38672
rect 1104 38032 6000 38128
rect 578000 38032 582820 38128
rect 1104 37488 6000 37584
rect 578000 37488 582820 37584
rect 1104 36944 6000 37040
rect 578000 36944 582820 37040
rect 1104 36400 6000 36496
rect 578000 36400 582820 36496
rect 1104 35856 6000 35952
rect 578000 35856 582820 35952
rect 3510 35776 3516 35828
rect 3568 35816 3574 35828
rect 7558 35816 7564 35828
rect 3568 35788 7564 35816
rect 3568 35776 3574 35788
rect 7558 35776 7564 35788
rect 7616 35776 7622 35828
rect 1104 35312 6000 35408
rect 578000 35312 582820 35408
rect 1104 34768 6000 34864
rect 578000 34768 582820 34864
rect 1104 34224 6000 34320
rect 578000 34224 582820 34320
rect 1104 33680 6000 33776
rect 578000 33680 582820 33776
rect 1104 33136 6000 33232
rect 578000 33136 582820 33232
rect 1104 32592 6000 32688
rect 578000 32592 582820 32688
rect 1104 32048 6000 32144
rect 578000 32048 582820 32144
rect 1104 31504 6000 31600
rect 578000 31504 582820 31600
rect 1104 30960 6000 31056
rect 578000 30960 582820 31056
rect 1104 30416 6000 30512
rect 578000 30416 582820 30512
rect 576118 30268 576124 30320
rect 576176 30308 576182 30320
rect 580166 30308 580172 30320
rect 576176 30280 580172 30308
rect 576176 30268 576182 30280
rect 580166 30268 580172 30280
rect 580224 30268 580230 30320
rect 1104 29872 6000 29968
rect 578000 29872 582820 29968
rect 1104 29328 6000 29424
rect 578000 29328 582820 29424
rect 1104 28784 6000 28880
rect 578000 28784 582820 28880
rect 1104 28240 6000 28336
rect 578000 28240 582820 28336
rect 1104 27696 6000 27792
rect 578000 27696 582820 27792
rect 1104 27152 6000 27248
rect 578000 27152 582820 27248
rect 1104 26608 6000 26704
rect 578000 26608 582820 26704
rect 1104 26064 6000 26160
rect 578000 26064 582820 26160
rect 1104 25520 6000 25616
rect 578000 25520 582820 25616
rect 1104 24976 6000 25072
rect 578000 24976 582820 25072
rect 1104 24432 6000 24528
rect 578000 24432 582820 24528
rect 1104 23888 6000 23984
rect 578000 23888 582820 23984
rect 1104 23344 6000 23440
rect 578000 23344 582820 23440
rect 1104 22800 6000 22896
rect 578000 22800 582820 22896
rect 1104 22256 6000 22352
rect 578000 22256 582820 22352
rect 1104 21712 6000 21808
rect 578000 21712 582820 21808
rect 1104 21168 6000 21264
rect 578000 21168 582820 21264
rect 1104 20624 6000 20720
rect 578000 20624 582820 20720
rect 1104 20080 6000 20176
rect 578000 20080 582820 20176
rect 1104 19536 6000 19632
rect 578000 19536 582820 19632
rect 1104 18992 6000 19088
rect 578000 18992 582820 19088
rect 1104 18448 6000 18544
rect 578000 18448 582820 18544
rect 1104 17904 6000 18000
rect 578000 17904 582820 18000
rect 575014 17824 575020 17876
rect 575072 17864 575078 17876
rect 580166 17864 580172 17876
rect 575072 17836 580172 17864
rect 575072 17824 575078 17836
rect 580166 17824 580172 17836
rect 580224 17824 580230 17876
rect 1104 17360 6000 17456
rect 578000 17360 582820 17456
rect 1104 16816 6000 16912
rect 578000 16816 582820 16912
rect 1104 16272 6000 16368
rect 578000 16272 582820 16368
rect 1104 15728 6000 15824
rect 578000 15728 582820 15824
rect 1104 15184 6000 15280
rect 578000 15184 582820 15280
rect 1104 14640 6000 14736
rect 578000 14640 582820 14736
rect 1104 14096 6000 14192
rect 578000 14096 582820 14192
rect 1104 13552 6000 13648
rect 578000 13552 582820 13648
rect 1104 13008 6000 13104
rect 578000 13008 582820 13104
rect 1104 12464 6000 12560
rect 578000 12464 582820 12560
rect 1104 11920 6000 12016
rect 578000 11920 582820 12016
rect 1104 11376 6000 11472
rect 578000 11376 582820 11472
rect 1104 10832 6000 10928
rect 578000 10832 582820 10928
rect 1104 10288 6000 10384
rect 578000 10288 582820 10384
rect 1104 9744 6000 9840
rect 578000 9744 582820 9840
rect 1104 9200 6000 9296
rect 578000 9200 582820 9296
rect 1104 8656 6000 8752
rect 578000 8656 582820 8752
rect 1104 8112 6000 8208
rect 578000 8112 582820 8208
rect 1104 7568 6000 7664
rect 578000 7568 582820 7664
rect 3142 7148 3148 7200
rect 3200 7188 3206 7200
rect 6178 7188 6184 7200
rect 3200 7160 6184 7188
rect 3200 7148 3206 7160
rect 6178 7148 6184 7160
rect 6236 7148 6242 7200
rect 1104 7024 6000 7120
rect 578000 7024 582820 7120
rect 484946 6808 484952 6860
rect 485004 6848 485010 6860
rect 495342 6848 495348 6860
rect 485004 6820 495348 6848
rect 485004 6808 485010 6820
rect 495342 6808 495348 6820
rect 495400 6808 495406 6860
rect 506658 6808 506664 6860
rect 506716 6848 506722 6860
rect 516134 6848 516140 6860
rect 506716 6820 516140 6848
rect 506716 6808 506722 6820
rect 516134 6808 516140 6820
rect 516192 6808 516198 6860
rect 519262 6808 519268 6860
rect 519320 6848 519326 6860
rect 531038 6848 531044 6860
rect 519320 6820 531044 6848
rect 519320 6808 519326 6820
rect 531038 6808 531044 6820
rect 531096 6808 531102 6860
rect 538766 6808 538772 6860
rect 538824 6848 538830 6860
rect 549530 6848 549536 6860
rect 538824 6820 549536 6848
rect 538824 6808 538830 6820
rect 549530 6808 549536 6820
rect 549588 6808 549594 6860
rect 560478 6808 560484 6860
rect 560536 6848 560542 6860
rect 570138 6848 570144 6860
rect 560536 6820 570144 6848
rect 560536 6808 560542 6820
rect 570138 6808 570144 6820
rect 570196 6808 570202 6860
rect 450538 6740 450544 6792
rect 450596 6780 450602 6792
rect 459646 6780 459652 6792
rect 450596 6752 459652 6780
rect 450596 6740 450602 6752
rect 459646 6740 459652 6752
rect 459704 6740 459710 6792
rect 494054 6740 494060 6792
rect 494112 6780 494118 6792
rect 504726 6780 504732 6792
rect 494112 6752 504732 6780
rect 494112 6740 494118 6752
rect 504726 6740 504732 6752
rect 504784 6740 504790 6792
rect 507854 6740 507860 6792
rect 507912 6780 507918 6792
rect 519078 6780 519084 6792
rect 507912 6752 519084 6780
rect 507912 6740 507918 6752
rect 519078 6740 519084 6752
rect 519136 6740 519142 6792
rect 520458 6740 520464 6792
rect 520516 6780 520522 6792
rect 532234 6780 532240 6792
rect 520516 6752 532240 6780
rect 520516 6740 520522 6752
rect 532234 6740 532240 6752
rect 532292 6740 532298 6792
rect 535270 6740 535276 6792
rect 535328 6780 535334 6792
rect 545114 6780 545120 6792
rect 535328 6752 545120 6780
rect 535328 6740 535334 6752
rect 545114 6740 545120 6752
rect 545172 6740 545178 6792
rect 546770 6740 546776 6792
rect 546828 6780 546834 6792
rect 556154 6780 556160 6792
rect 546828 6752 556160 6780
rect 546828 6740 546834 6752
rect 556154 6740 556160 6752
rect 556212 6740 556218 6792
rect 561674 6740 561680 6792
rect 561732 6780 561738 6792
rect 571334 6780 571340 6792
rect 561732 6752 571340 6780
rect 561732 6740 561738 6752
rect 571334 6740 571340 6752
rect 571392 6740 571398 6792
rect 458542 6672 458548 6724
rect 458600 6712 458606 6724
rect 467926 6712 467932 6724
rect 458600 6684 467932 6712
rect 458600 6672 458606 6684
rect 467926 6672 467932 6684
rect 467984 6672 467990 6724
rect 476942 6672 476948 6724
rect 477000 6712 477006 6724
rect 486694 6712 486700 6724
rect 477000 6684 486700 6712
rect 477000 6672 477006 6684
rect 486694 6672 486700 6684
rect 486752 6672 486758 6724
rect 492950 6672 492956 6724
rect 493008 6712 493014 6724
rect 503622 6712 503628 6724
rect 493008 6684 503628 6712
rect 493008 6672 493014 6684
rect 503622 6672 503628 6684
rect 503680 6672 503686 6724
rect 511258 6672 511264 6724
rect 511316 6712 511322 6724
rect 522666 6712 522672 6724
rect 511316 6684 522672 6712
rect 511316 6672 511322 6684
rect 522666 6672 522672 6684
rect 522724 6672 522730 6724
rect 527266 6672 527272 6724
rect 527324 6712 527330 6724
rect 539318 6712 539324 6724
rect 527324 6684 539324 6712
rect 527324 6672 527330 6684
rect 539318 6672 539324 6684
rect 539376 6672 539382 6724
rect 545574 6672 545580 6724
rect 545632 6712 545638 6724
rect 556246 6712 556252 6724
rect 545632 6684 556252 6712
rect 545632 6672 545638 6684
rect 556246 6672 556252 6684
rect 556304 6672 556310 6724
rect 558178 6672 558184 6724
rect 558236 6712 558242 6724
rect 568206 6712 568212 6724
rect 558236 6684 568212 6712
rect 558236 6672 558242 6684
rect 568206 6672 568212 6684
rect 568264 6672 568270 6724
rect 470042 6604 470048 6656
rect 470100 6644 470106 6656
rect 479886 6644 479892 6656
rect 470100 6616 479892 6644
rect 470100 6604 470106 6616
rect 479886 6604 479892 6616
rect 479944 6604 479950 6656
rect 486050 6604 486056 6656
rect 486108 6644 486114 6656
rect 496538 6644 496544 6656
rect 486108 6616 496544 6644
rect 486108 6604 486114 6616
rect 496538 6604 496544 6616
rect 496596 6604 496602 6656
rect 505554 6604 505560 6656
rect 505612 6644 505618 6656
rect 516778 6644 516784 6656
rect 505612 6616 516784 6644
rect 505612 6604 505618 6616
rect 516778 6604 516784 6616
rect 516836 6604 516842 6656
rect 526162 6604 526168 6656
rect 526220 6644 526226 6656
rect 538122 6644 538128 6656
rect 526220 6616 538128 6644
rect 526220 6604 526226 6616
rect 538122 6604 538128 6616
rect 538180 6604 538186 6656
rect 541066 6604 541072 6656
rect 541124 6644 541130 6656
rect 553302 6644 553308 6656
rect 541124 6616 553308 6644
rect 541124 6604 541130 6616
rect 553302 6604 553308 6616
rect 553360 6604 553366 6656
rect 557074 6604 557080 6656
rect 557132 6644 557138 6656
rect 568390 6644 568396 6656
rect 557132 6616 568396 6644
rect 557132 6604 557138 6616
rect 568390 6604 568396 6616
rect 568448 6604 568454 6656
rect 1104 6480 6000 6576
rect 468846 6536 468852 6588
rect 468904 6576 468910 6588
rect 478690 6576 478696 6588
rect 468904 6548 478696 6576
rect 468904 6536 468910 6548
rect 478690 6536 478696 6548
rect 478748 6536 478754 6588
rect 479150 6536 479156 6588
rect 479208 6576 479214 6588
rect 489362 6576 489368 6588
rect 479208 6548 489368 6576
rect 479208 6536 479214 6548
rect 489362 6536 489368 6548
rect 489420 6536 489426 6588
rect 490650 6536 490656 6588
rect 490708 6576 490714 6588
rect 501230 6576 501236 6588
rect 490708 6548 501236 6576
rect 490708 6536 490714 6548
rect 501230 6536 501236 6548
rect 501288 6536 501294 6588
rect 504358 6536 504364 6588
rect 504416 6576 504422 6588
rect 515582 6576 515588 6588
rect 504416 6548 515588 6576
rect 504416 6536 504422 6548
rect 515582 6536 515588 6548
rect 515640 6536 515646 6588
rect 521562 6536 521568 6588
rect 521620 6576 521626 6588
rect 531314 6576 531320 6588
rect 521620 6548 531320 6576
rect 521620 6536 521626 6548
rect 531314 6536 531320 6548
rect 531372 6536 531378 6588
rect 543366 6536 543372 6588
rect 543424 6576 543430 6588
rect 553394 6576 553400 6588
rect 543424 6548 553400 6576
rect 543424 6536 543430 6548
rect 553394 6536 553400 6548
rect 553452 6536 553458 6588
rect 559374 6536 559380 6588
rect 559432 6576 559438 6588
rect 572622 6576 572628 6588
rect 559432 6548 572628 6576
rect 559432 6536 559438 6548
rect 572622 6536 572628 6548
rect 572680 6536 572686 6588
rect 119430 6468 119436 6520
rect 119488 6508 119494 6520
rect 123018 6508 123024 6520
rect 119488 6480 123024 6508
rect 119488 6468 119494 6480
rect 123018 6468 123024 6480
rect 123076 6468 123082 6520
rect 407022 6468 407028 6520
rect 407080 6508 407086 6520
rect 408494 6508 408500 6520
rect 407080 6480 408500 6508
rect 407080 6468 407086 6480
rect 408494 6468 408500 6480
rect 408552 6468 408558 6520
rect 466638 6468 466644 6520
rect 466696 6508 466702 6520
rect 476298 6508 476304 6520
rect 466696 6480 476304 6508
rect 466696 6468 466702 6480
rect 476298 6468 476304 6480
rect 476356 6468 476362 6520
rect 483750 6468 483756 6520
rect 483808 6508 483814 6520
rect 494146 6508 494152 6520
rect 483808 6480 494152 6508
rect 483808 6468 483814 6480
rect 494146 6468 494152 6480
rect 494204 6468 494210 6520
rect 495250 6468 495256 6520
rect 495308 6508 495314 6520
rect 506014 6508 506020 6520
rect 495308 6480 506020 6508
rect 495308 6468 495314 6480
rect 506014 6468 506020 6480
rect 506072 6468 506078 6520
rect 510154 6468 510160 6520
rect 510212 6508 510218 6520
rect 521470 6508 521476 6520
rect 510212 6480 521476 6508
rect 510212 6468 510218 6480
rect 521470 6468 521476 6480
rect 521528 6468 521534 6520
rect 524966 6468 524972 6520
rect 525024 6508 525030 6520
rect 536742 6508 536748 6520
rect 525024 6480 536748 6508
rect 525024 6468 525030 6480
rect 536742 6468 536748 6480
rect 536800 6468 536806 6520
rect 537570 6468 537576 6520
rect 537628 6508 537634 6520
rect 546586 6508 546592 6520
rect 537628 6480 546592 6508
rect 537628 6468 537634 6480
rect 546586 6468 546592 6480
rect 546644 6468 546650 6520
rect 550174 6468 550180 6520
rect 550232 6508 550238 6520
rect 560386 6508 560392 6520
rect 550232 6480 560392 6508
rect 550232 6468 550238 6480
rect 560386 6468 560392 6480
rect 560444 6468 560450 6520
rect 563974 6468 563980 6520
rect 564032 6508 564038 6520
rect 575474 6508 575480 6520
rect 564032 6480 575480 6508
rect 564032 6468 564038 6480
rect 575474 6468 575480 6480
rect 575532 6468 575538 6520
rect 578000 6480 582820 6576
rect 88518 6400 88524 6452
rect 88576 6440 88582 6452
rect 93302 6440 93308 6452
rect 88576 6412 93308 6440
rect 88576 6400 88582 6412
rect 93302 6400 93308 6412
rect 93360 6400 93366 6452
rect 102778 6400 102784 6452
rect 102836 6440 102842 6452
rect 107010 6440 107016 6452
rect 102836 6412 107016 6440
rect 102836 6400 102842 6412
rect 107010 6400 107016 6412
rect 107068 6400 107074 6452
rect 120626 6400 120632 6452
rect 120684 6440 120690 6452
rect 124214 6440 124220 6452
rect 120684 6412 124220 6440
rect 120684 6400 120690 6412
rect 124214 6400 124220 6412
rect 124272 6400 124278 6452
rect 464338 6400 464344 6452
rect 464396 6440 464402 6452
rect 473906 6440 473912 6452
rect 464396 6412 473912 6440
rect 464396 6400 464402 6412
rect 473906 6400 473912 6412
rect 473964 6400 473970 6452
rect 475746 6400 475752 6452
rect 475804 6440 475810 6452
rect 485682 6440 485688 6452
rect 475804 6412 485688 6440
rect 475804 6400 475810 6412
rect 485682 6400 485688 6412
rect 485740 6400 485746 6452
rect 502058 6400 502064 6452
rect 502116 6440 502122 6452
rect 510982 6440 510988 6452
rect 502116 6412 510988 6440
rect 502116 6400 502122 6412
rect 510982 6400 510988 6412
rect 511040 6400 511046 6452
rect 512362 6400 512368 6452
rect 512420 6440 512426 6452
rect 523862 6440 523868 6452
rect 512420 6412 523868 6440
rect 512420 6400 512426 6412
rect 523862 6400 523868 6412
rect 523920 6400 523926 6452
rect 530762 6400 530768 6452
rect 530820 6440 530826 6452
rect 541526 6440 541532 6452
rect 530820 6412 541532 6440
rect 530820 6400 530826 6412
rect 541526 6400 541532 6412
rect 541584 6400 541590 6452
rect 544470 6400 544476 6452
rect 544528 6440 544534 6452
rect 554866 6440 554872 6452
rect 544528 6412 554872 6440
rect 544528 6400 544534 6412
rect 554866 6400 554872 6412
rect 554924 6400 554930 6452
rect 565078 6400 565084 6452
rect 565136 6440 565142 6452
rect 577682 6440 577688 6452
rect 565136 6412 577688 6440
rect 565136 6400 565142 6412
rect 577682 6400 577688 6412
rect 577740 6400 577746 6452
rect 151538 6332 151544 6384
rect 151596 6372 151602 6384
rect 153930 6372 153936 6384
rect 151596 6344 153936 6372
rect 151596 6332 151602 6344
rect 153930 6332 153936 6344
rect 153988 6332 153994 6384
rect 313182 6332 313188 6384
rect 313240 6372 313246 6384
rect 314654 6372 314660 6384
rect 313240 6344 314660 6372
rect 313240 6332 313246 6344
rect 314654 6332 314660 6344
rect 314712 6332 314718 6384
rect 340598 6332 340604 6384
rect 340656 6372 340662 6384
rect 342714 6372 342720 6384
rect 340656 6344 342720 6372
rect 340656 6332 340662 6344
rect 342714 6332 342720 6344
rect 342772 6332 342778 6384
rect 370406 6332 370412 6384
rect 370464 6372 370470 6384
rect 372614 6372 372620 6384
rect 370464 6344 372620 6372
rect 370464 6332 370470 6344
rect 372614 6332 372620 6344
rect 372672 6332 372678 6384
rect 379606 6332 379612 6384
rect 379664 6372 379670 6384
rect 382366 6372 382372 6384
rect 379664 6344 382372 6372
rect 379664 6332 379670 6344
rect 382366 6332 382372 6344
rect 382424 6332 382430 6384
rect 416222 6332 416228 6384
rect 416280 6372 416286 6384
rect 418154 6372 418160 6384
rect 416280 6344 418160 6372
rect 416280 6332 416286 6344
rect 418154 6332 418160 6344
rect 418212 6332 418218 6384
rect 442534 6332 442540 6384
rect 442592 6372 442598 6384
rect 445478 6372 445484 6384
rect 442592 6344 445484 6372
rect 442592 6332 442598 6344
rect 445478 6332 445484 6344
rect 445536 6332 445542 6384
rect 449434 6332 449440 6384
rect 449492 6372 449498 6384
rect 458450 6372 458456 6384
rect 449492 6344 458456 6372
rect 449492 6332 449498 6344
rect 458450 6332 458456 6344
rect 458508 6332 458514 6384
rect 463142 6332 463148 6384
rect 463200 6372 463206 6384
rect 472710 6372 472716 6384
rect 463200 6344 472716 6372
rect 463200 6332 463206 6344
rect 472710 6332 472716 6344
rect 472768 6332 472774 6384
rect 474642 6332 474648 6384
rect 474700 6372 474706 6384
rect 484578 6372 484584 6384
rect 474700 6344 484584 6372
rect 474700 6332 474706 6344
rect 484578 6332 484584 6344
rect 484636 6332 484642 6384
rect 489454 6332 489460 6384
rect 489512 6372 489518 6384
rect 500126 6372 500132 6384
rect 489512 6344 500132 6372
rect 489512 6332 489518 6344
rect 500126 6332 500132 6344
rect 500184 6332 500190 6384
rect 500218 6332 500224 6384
rect 500276 6372 500282 6384
rect 510798 6372 510804 6384
rect 500276 6344 510804 6372
rect 500276 6332 500282 6344
rect 510798 6332 510804 6344
rect 510856 6332 510862 6384
rect 513558 6332 513564 6384
rect 513616 6372 513622 6384
rect 525058 6372 525064 6384
rect 513616 6344 525064 6372
rect 513616 6332 513622 6344
rect 525058 6332 525064 6344
rect 525116 6332 525122 6384
rect 529566 6332 529572 6384
rect 529624 6372 529630 6384
rect 539962 6372 539968 6384
rect 529624 6344 539968 6372
rect 529624 6332 529630 6344
rect 539962 6332 539968 6344
rect 540020 6332 540026 6384
rect 542170 6332 542176 6384
rect 542228 6372 542234 6384
rect 552014 6372 552020 6384
rect 542228 6344 552020 6372
rect 542228 6332 542234 6344
rect 552014 6332 552020 6344
rect 552072 6332 552078 6384
rect 562778 6332 562784 6384
rect 562836 6372 562842 6384
rect 576210 6372 576216 6384
rect 562836 6344 576216 6372
rect 562836 6332 562842 6344
rect 576210 6332 576216 6344
rect 576268 6332 576274 6384
rect 93302 6264 93308 6316
rect 93360 6304 93366 6316
rect 97810 6304 97816 6316
rect 93360 6276 97816 6304
rect 93360 6264 93366 6276
rect 97810 6264 97816 6276
rect 97868 6264 97874 6316
rect 418522 6264 418528 6316
rect 418580 6304 418586 6316
rect 420914 6304 420920 6316
rect 418580 6276 420920 6304
rect 418580 6264 418586 6276
rect 420914 6264 420920 6276
rect 420972 6264 420978 6316
rect 465442 6264 465448 6316
rect 465500 6304 465506 6316
rect 475102 6304 475108 6316
rect 465500 6276 475108 6304
rect 465500 6264 465506 6276
rect 475102 6264 475108 6276
rect 475160 6264 475166 6316
rect 481450 6264 481456 6316
rect 481508 6304 481514 6316
rect 491754 6304 491760 6316
rect 481508 6276 491760 6304
rect 481508 6264 481514 6276
rect 491754 6264 491760 6276
rect 491812 6264 491818 6316
rect 496354 6264 496360 6316
rect 496412 6304 496418 6316
rect 507210 6304 507216 6316
rect 496412 6276 507216 6304
rect 496412 6264 496418 6276
rect 507210 6264 507216 6276
rect 507268 6264 507274 6316
rect 514662 6264 514668 6316
rect 514720 6304 514726 6316
rect 524414 6304 524420 6316
rect 514720 6276 524420 6304
rect 514720 6264 514726 6276
rect 524414 6264 524420 6276
rect 524472 6264 524478 6316
rect 528462 6264 528468 6316
rect 528520 6304 528526 6316
rect 539410 6304 539416 6316
rect 528520 6276 539416 6304
rect 528520 6264 528526 6276
rect 539410 6264 539416 6276
rect 539468 6264 539474 6316
rect 539870 6264 539876 6316
rect 539928 6304 539934 6316
rect 550634 6304 550640 6316
rect 539928 6276 550640 6304
rect 539928 6264 539934 6276
rect 550634 6264 550640 6276
rect 550692 6264 550698 6316
rect 554774 6264 554780 6316
rect 554832 6304 554838 6316
rect 564434 6304 564440 6316
rect 554832 6276 564440 6304
rect 554832 6264 554838 6276
rect 564434 6264 564440 6276
rect 564492 6264 564498 6316
rect 566182 6264 566188 6316
rect 566240 6304 566246 6316
rect 579798 6304 579804 6316
rect 566240 6276 579804 6304
rect 566240 6264 566246 6276
rect 579798 6264 579804 6276
rect 579856 6264 579862 6316
rect 161106 6196 161112 6248
rect 161164 6236 161170 6248
rect 163130 6236 163136 6248
rect 161164 6208 163136 6236
rect 161164 6196 161170 6208
rect 163130 6196 163136 6208
rect 163188 6196 163194 6248
rect 361206 6196 361212 6248
rect 361264 6236 361270 6248
rect 362954 6236 362960 6248
rect 361264 6208 362960 6236
rect 361264 6196 361270 6208
rect 362954 6196 362960 6208
rect 363012 6196 363018 6248
rect 415026 6196 415032 6248
rect 415084 6236 415090 6248
rect 416958 6236 416964 6248
rect 415084 6208 416964 6236
rect 415084 6196 415090 6208
rect 416958 6196 416964 6208
rect 417016 6196 417022 6248
rect 427630 6196 427636 6248
rect 427688 6236 427694 6248
rect 429838 6236 429844 6248
rect 427688 6208 429844 6236
rect 427688 6196 427694 6208
rect 429838 6196 429844 6208
rect 429896 6196 429902 6248
rect 433426 6196 433432 6248
rect 433484 6236 433490 6248
rect 436094 6236 436100 6248
rect 433484 6208 436100 6236
rect 433484 6196 433490 6208
rect 436094 6196 436100 6208
rect 436152 6196 436158 6248
rect 437934 6196 437940 6248
rect 437992 6236 437998 6248
rect 440326 6236 440332 6248
rect 437992 6208 440332 6236
rect 437992 6196 437998 6208
rect 440326 6196 440332 6208
rect 440384 6196 440390 6248
rect 448238 6196 448244 6248
rect 448296 6236 448302 6248
rect 457254 6236 457260 6248
rect 448296 6208 457260 6236
rect 448296 6196 448302 6208
rect 457254 6196 457260 6208
rect 457312 6196 457318 6248
rect 462038 6196 462044 6248
rect 462096 6236 462102 6248
rect 471514 6236 471520 6248
rect 462096 6208 471520 6236
rect 462096 6196 462102 6208
rect 471514 6196 471520 6208
rect 471572 6196 471578 6248
rect 473446 6196 473452 6248
rect 473504 6236 473510 6248
rect 483474 6236 483480 6248
rect 473504 6208 483480 6236
rect 473504 6196 473510 6208
rect 483474 6196 483480 6208
rect 483532 6196 483538 6248
rect 487246 6196 487252 6248
rect 487304 6236 487310 6248
rect 490742 6236 490748 6248
rect 487304 6208 490748 6236
rect 487304 6196 487310 6208
rect 490742 6196 490748 6208
rect 490800 6196 490806 6248
rect 497550 6196 497556 6248
rect 497608 6236 497614 6248
rect 508406 6236 508412 6248
rect 497608 6208 508412 6236
rect 497608 6196 497614 6208
rect 508406 6196 508412 6208
rect 508464 6196 508470 6248
rect 508958 6196 508964 6248
rect 509016 6236 509022 6248
rect 520182 6236 520188 6248
rect 509016 6208 520188 6236
rect 509016 6196 509022 6208
rect 520182 6196 520188 6208
rect 520240 6196 520246 6248
rect 524138 6196 524144 6248
rect 524196 6236 524202 6248
rect 535362 6236 535368 6248
rect 524196 6208 535368 6236
rect 524196 6196 524202 6208
rect 535362 6196 535368 6208
rect 535420 6196 535426 6248
rect 536466 6196 536472 6248
rect 536524 6236 536530 6248
rect 546494 6236 546500 6248
rect 536524 6208 546500 6236
rect 536524 6196 536530 6208
rect 546494 6196 546500 6208
rect 546552 6196 546558 6248
rect 551370 6196 551376 6248
rect 551428 6236 551434 6248
rect 561766 6236 561772 6248
rect 551428 6208 561772 6236
rect 551428 6196 551434 6208
rect 561766 6196 561772 6208
rect 561824 6196 561830 6248
rect 567378 6196 567384 6248
rect 567436 6236 567442 6248
rect 580994 6236 581000 6248
rect 567436 6208 581000 6236
rect 567436 6196 567442 6208
rect 580994 6196 581000 6208
rect 581052 6196 581058 6248
rect 5534 6128 5540 6180
rect 5592 6168 5598 6180
rect 10778 6168 10784 6180
rect 5592 6140 10784 6168
rect 5592 6128 5598 6140
rect 10778 6128 10784 6140
rect 10836 6128 10842 6180
rect 17586 6128 17592 6180
rect 17644 6168 17650 6180
rect 18874 6168 18880 6180
rect 17644 6140 18880 6168
rect 17644 6128 17650 6140
rect 18874 6128 18880 6140
rect 18932 6128 18938 6180
rect 86126 6128 86132 6180
rect 86184 6168 86190 6180
rect 91002 6168 91008 6180
rect 86184 6140 91008 6168
rect 86184 6128 86190 6140
rect 91002 6128 91008 6140
rect 91060 6128 91066 6180
rect 112346 6128 112352 6180
rect 112404 6168 112410 6180
rect 116210 6168 116216 6180
rect 112404 6140 116216 6168
rect 112404 6128 112410 6140
rect 116210 6128 116216 6140
rect 116268 6128 116274 6180
rect 270770 6128 270776 6180
rect 270828 6168 270834 6180
rect 272886 6168 272892 6180
rect 270828 6140 272892 6168
rect 270828 6128 270834 6140
rect 272886 6128 272892 6140
rect 272944 6128 272950 6180
rect 307386 6128 307392 6180
rect 307444 6168 307450 6180
rect 309134 6168 309140 6180
rect 307444 6140 309140 6168
rect 307444 6128 307450 6140
rect 309134 6128 309140 6140
rect 309192 6128 309198 6180
rect 322290 6128 322296 6180
rect 322348 6168 322354 6180
rect 324314 6168 324320 6180
rect 322348 6140 324320 6168
rect 322348 6128 322354 6140
rect 324314 6128 324320 6140
rect 324372 6128 324378 6180
rect 342898 6128 342904 6180
rect 342956 6168 342962 6180
rect 346118 6168 346124 6180
rect 342956 6140 346124 6168
rect 342956 6128 342962 6140
rect 346118 6128 346124 6140
rect 346176 6128 346182 6180
rect 434530 6128 434536 6180
rect 434588 6168 434594 6180
rect 442994 6168 443000 6180
rect 434588 6140 443000 6168
rect 434588 6128 434594 6140
rect 442994 6128 443000 6140
rect 443052 6128 443058 6180
rect 455138 6128 455144 6180
rect 455196 6168 455202 6180
rect 464430 6168 464436 6180
rect 455196 6140 464436 6168
rect 455196 6128 455202 6140
rect 464430 6128 464436 6140
rect 464488 6128 464494 6180
rect 467742 6128 467748 6180
rect 467800 6168 467806 6180
rect 477494 6168 477500 6180
rect 467800 6140 477500 6168
rect 467800 6128 467806 6140
rect 477494 6128 477500 6140
rect 477552 6128 477558 6180
rect 482646 6128 482652 6180
rect 482704 6168 482710 6180
rect 492950 6168 492956 6180
rect 482704 6140 492956 6168
rect 482704 6128 482710 6140
rect 492950 6128 492956 6140
rect 493008 6128 493014 6180
rect 498654 6128 498660 6180
rect 498712 6168 498718 6180
rect 509602 6168 509608 6180
rect 498712 6140 509608 6168
rect 498712 6128 498718 6140
rect 509602 6128 509608 6140
rect 509660 6128 509666 6180
rect 515858 6128 515864 6180
rect 515916 6168 515922 6180
rect 527082 6168 527088 6180
rect 515916 6140 527088 6168
rect 515916 6128 515922 6140
rect 527082 6128 527088 6140
rect 527140 6128 527146 6180
rect 534166 6128 534172 6180
rect 534224 6168 534230 6180
rect 546402 6168 546408 6180
rect 534224 6140 546408 6168
rect 534224 6128 534230 6140
rect 546402 6128 546408 6140
rect 546460 6128 546466 6180
rect 553670 6128 553676 6180
rect 553728 6168 553734 6180
rect 564618 6168 564624 6180
rect 553728 6140 564624 6168
rect 553728 6128 553734 6140
rect 564618 6128 564624 6140
rect 564676 6128 564682 6180
rect 568482 6128 568488 6180
rect 568540 6168 568546 6180
rect 582190 6168 582196 6180
rect 568540 6140 582196 6168
rect 568540 6128 568546 6140
rect 582190 6128 582196 6140
rect 582248 6128 582254 6180
rect 341794 6060 341800 6112
rect 341852 6100 341858 6112
rect 343634 6100 343640 6112
rect 341852 6072 343640 6100
rect 341852 6060 341858 6072
rect 343634 6060 343640 6072
rect 343692 6060 343698 6112
rect 350902 6060 350908 6112
rect 350960 6100 350966 6112
rect 353294 6100 353300 6112
rect 350960 6072 353300 6100
rect 350960 6060 350966 6072
rect 353294 6060 353300 6072
rect 353352 6060 353358 6112
rect 355502 6060 355508 6112
rect 355560 6100 355566 6112
rect 358170 6100 358176 6112
rect 355560 6072 358176 6100
rect 355560 6060 355566 6072
rect 358170 6060 358176 6072
rect 358228 6060 358234 6112
rect 360102 6060 360108 6112
rect 360160 6100 360166 6112
rect 362218 6100 362224 6112
rect 360160 6072 362224 6100
rect 360160 6060 360166 6072
rect 362218 6060 362224 6072
rect 362276 6060 362282 6112
rect 369210 6060 369216 6112
rect 369268 6100 369274 6112
rect 371602 6100 371608 6112
rect 369268 6072 371608 6100
rect 369268 6060 369274 6072
rect 371602 6060 371608 6072
rect 371660 6060 371666 6112
rect 388714 6060 388720 6112
rect 388772 6100 388778 6112
rect 391106 6100 391112 6112
rect 388772 6072 391112 6100
rect 388772 6060 388778 6072
rect 391106 6060 391112 6072
rect 391164 6060 391170 6112
rect 419626 6060 419632 6112
rect 419684 6100 419690 6112
rect 423582 6100 423588 6112
rect 419684 6072 423588 6100
rect 419684 6060 419690 6072
rect 423582 6060 423588 6072
rect 423640 6060 423646 6112
rect 436830 6060 436836 6112
rect 436888 6100 436894 6112
rect 439222 6100 439228 6112
rect 436888 6072 439228 6100
rect 436888 6060 436894 6072
rect 439222 6060 439228 6072
rect 439280 6060 439286 6112
rect 447134 6060 447140 6112
rect 447192 6100 447198 6112
rect 449894 6100 449900 6112
rect 447192 6072 449900 6100
rect 447192 6060 447198 6072
rect 449894 6060 449900 6072
rect 449952 6060 449958 6112
rect 454034 6060 454040 6112
rect 454092 6100 454098 6112
rect 457530 6100 457536 6112
rect 454092 6072 457536 6100
rect 454092 6060 454098 6072
rect 457530 6060 457536 6072
rect 457588 6060 457594 6112
rect 460842 6060 460848 6112
rect 460900 6100 460906 6112
rect 470318 6100 470324 6112
rect 460900 6072 470324 6100
rect 460900 6060 460906 6072
rect 470318 6060 470324 6072
rect 470376 6060 470382 6112
rect 478046 6060 478052 6112
rect 478104 6100 478110 6112
rect 488166 6100 488172 6112
rect 478104 6072 488172 6100
rect 478104 6060 478110 6072
rect 488166 6060 488172 6072
rect 488224 6060 488230 6112
rect 500954 6060 500960 6112
rect 501012 6100 501018 6112
rect 511902 6100 511908 6112
rect 501012 6072 511908 6100
rect 501012 6060 501018 6072
rect 511902 6060 511908 6072
rect 511960 6060 511966 6112
rect 522574 6060 522580 6112
rect 522632 6100 522638 6112
rect 531498 6100 531504 6112
rect 522632 6072 531504 6100
rect 522632 6060 522638 6072
rect 531498 6060 531504 6072
rect 531556 6060 531562 6112
rect 552474 6060 552480 6112
rect 552532 6100 552538 6112
rect 561674 6100 561680 6112
rect 552532 6072 561680 6100
rect 552532 6060 552538 6072
rect 561674 6060 561680 6072
rect 561732 6060 561738 6112
rect 1104 6010 582820 6032
rect 1104 5958 18822 6010
rect 18874 5958 18886 6010
rect 18938 5958 18950 6010
rect 19002 5958 19014 6010
rect 19066 5958 19078 6010
rect 19130 5958 19142 6010
rect 19194 5958 19206 6010
rect 19258 5958 19270 6010
rect 19322 5958 19334 6010
rect 19386 5958 54822 6010
rect 54874 5958 54886 6010
rect 54938 5958 54950 6010
rect 55002 5958 55014 6010
rect 55066 5958 55078 6010
rect 55130 5958 55142 6010
rect 55194 5958 55206 6010
rect 55258 5958 55270 6010
rect 55322 5958 55334 6010
rect 55386 5958 90822 6010
rect 90874 5958 90886 6010
rect 90938 5958 90950 6010
rect 91002 5958 91014 6010
rect 91066 5958 91078 6010
rect 91130 5958 91142 6010
rect 91194 5958 91206 6010
rect 91258 5958 91270 6010
rect 91322 5958 91334 6010
rect 91386 5958 126822 6010
rect 126874 5958 126886 6010
rect 126938 5958 126950 6010
rect 127002 5958 127014 6010
rect 127066 5958 127078 6010
rect 127130 5958 127142 6010
rect 127194 5958 127206 6010
rect 127258 5958 127270 6010
rect 127322 5958 127334 6010
rect 127386 5958 162822 6010
rect 162874 5958 162886 6010
rect 162938 5958 162950 6010
rect 163002 5958 163014 6010
rect 163066 5958 163078 6010
rect 163130 5958 163142 6010
rect 163194 5958 163206 6010
rect 163258 5958 163270 6010
rect 163322 5958 163334 6010
rect 163386 5958 198822 6010
rect 198874 5958 198886 6010
rect 198938 5958 198950 6010
rect 199002 5958 199014 6010
rect 199066 5958 199078 6010
rect 199130 5958 199142 6010
rect 199194 5958 199206 6010
rect 199258 5958 199270 6010
rect 199322 5958 199334 6010
rect 199386 5958 234822 6010
rect 234874 5958 234886 6010
rect 234938 5958 234950 6010
rect 235002 5958 235014 6010
rect 235066 5958 235078 6010
rect 235130 5958 235142 6010
rect 235194 5958 235206 6010
rect 235258 5958 235270 6010
rect 235322 5958 235334 6010
rect 235386 5958 270822 6010
rect 270874 5958 270886 6010
rect 270938 5958 270950 6010
rect 271002 5958 271014 6010
rect 271066 5958 271078 6010
rect 271130 5958 271142 6010
rect 271194 5958 271206 6010
rect 271258 5958 271270 6010
rect 271322 5958 271334 6010
rect 271386 5958 306822 6010
rect 306874 5958 306886 6010
rect 306938 5958 306950 6010
rect 307002 5958 307014 6010
rect 307066 5958 307078 6010
rect 307130 5958 307142 6010
rect 307194 5958 307206 6010
rect 307258 5958 307270 6010
rect 307322 5958 307334 6010
rect 307386 5958 342822 6010
rect 342874 5958 342886 6010
rect 342938 5958 342950 6010
rect 343002 5958 343014 6010
rect 343066 5958 343078 6010
rect 343130 5958 343142 6010
rect 343194 5958 343206 6010
rect 343258 5958 343270 6010
rect 343322 5958 343334 6010
rect 343386 5958 378822 6010
rect 378874 5958 378886 6010
rect 378938 5958 378950 6010
rect 379002 5958 379014 6010
rect 379066 5958 379078 6010
rect 379130 5958 379142 6010
rect 379194 5958 379206 6010
rect 379258 5958 379270 6010
rect 379322 5958 379334 6010
rect 379386 5958 414822 6010
rect 414874 5958 414886 6010
rect 414938 5958 414950 6010
rect 415002 5958 415014 6010
rect 415066 5958 415078 6010
rect 415130 5958 415142 6010
rect 415194 5958 415206 6010
rect 415258 5958 415270 6010
rect 415322 5958 415334 6010
rect 415386 5958 450822 6010
rect 450874 5958 450886 6010
rect 450938 5958 450950 6010
rect 451002 5958 451014 6010
rect 451066 5958 451078 6010
rect 451130 5958 451142 6010
rect 451194 5958 451206 6010
rect 451258 5958 451270 6010
rect 451322 5958 451334 6010
rect 451386 5958 486822 6010
rect 486874 5958 486886 6010
rect 486938 5958 486950 6010
rect 487002 5958 487014 6010
rect 487066 5958 487078 6010
rect 487130 5958 487142 6010
rect 487194 5958 487206 6010
rect 487258 5958 487270 6010
rect 487322 5958 487334 6010
rect 487386 5958 522822 6010
rect 522874 5958 522886 6010
rect 522938 5958 522950 6010
rect 523002 5958 523014 6010
rect 523066 5958 523078 6010
rect 523130 5958 523142 6010
rect 523194 5958 523206 6010
rect 523258 5958 523270 6010
rect 523322 5958 523334 6010
rect 523386 5958 558822 6010
rect 558874 5958 558886 6010
rect 558938 5958 558950 6010
rect 559002 5958 559014 6010
rect 559066 5958 559078 6010
rect 559130 5958 559142 6010
rect 559194 5958 559206 6010
rect 559258 5958 559270 6010
rect 559322 5958 559334 6010
rect 559386 5958 582820 6010
rect 1104 5936 582820 5958
rect 331490 5856 331496 5908
rect 331548 5896 331554 5908
rect 333974 5896 333980 5908
rect 331548 5868 333980 5896
rect 331548 5856 331554 5868
rect 333974 5856 333980 5868
rect 334032 5856 334038 5908
rect 402422 5856 402428 5908
rect 402480 5896 402486 5908
rect 405642 5896 405648 5908
rect 402480 5868 405648 5896
rect 402480 5856 402486 5868
rect 405642 5856 405648 5868
rect 405700 5856 405706 5908
rect 410518 5856 410524 5908
rect 410576 5896 410582 5908
rect 413738 5896 413744 5908
rect 410576 5868 413744 5896
rect 410576 5856 410582 5868
rect 413738 5856 413744 5868
rect 413796 5856 413802 5908
rect 421926 5856 421932 5908
rect 421984 5896 421990 5908
rect 424502 5896 424508 5908
rect 421984 5868 424508 5896
rect 421984 5856 421990 5868
rect 424502 5856 424508 5868
rect 424560 5856 424566 5908
rect 431126 5856 431132 5908
rect 431184 5896 431190 5908
rect 434162 5896 434168 5908
rect 431184 5868 434168 5896
rect 431184 5856 431190 5868
rect 434162 5856 434168 5868
rect 434220 5856 434226 5908
rect 440234 5856 440240 5908
rect 440292 5896 440298 5908
rect 443822 5896 443828 5908
rect 440292 5868 443828 5896
rect 440292 5856 440298 5868
rect 443822 5856 443828 5868
rect 443880 5856 443886 5908
rect 480346 5856 480352 5908
rect 480404 5896 480410 5908
rect 490558 5896 490564 5908
rect 480404 5868 490564 5896
rect 480404 5856 480410 5868
rect 490558 5856 490564 5868
rect 490616 5856 490622 5908
rect 491662 5856 491668 5908
rect 491720 5896 491726 5908
rect 502242 5896 502248 5908
rect 491720 5868 502248 5896
rect 491720 5856 491726 5868
rect 502242 5856 502248 5868
rect 502300 5856 502306 5908
rect 516962 5856 516968 5908
rect 517020 5896 517026 5908
rect 525794 5896 525800 5908
rect 517020 5868 525800 5896
rect 517020 5856 517026 5868
rect 525794 5856 525800 5868
rect 525852 5856 525858 5908
rect 531866 5856 531872 5908
rect 531924 5896 531930 5908
rect 541434 5896 541440 5908
rect 531924 5868 541440 5896
rect 531924 5856 531930 5868
rect 541434 5856 541440 5868
rect 541492 5856 541498 5908
rect 555878 5856 555884 5908
rect 555936 5896 555942 5908
rect 564526 5896 564532 5908
rect 555936 5868 564532 5896
rect 555936 5856 555942 5868
rect 564526 5856 564532 5868
rect 564584 5856 564590 5908
rect 105170 5788 105176 5840
rect 105228 5828 105234 5840
rect 109310 5828 109316 5840
rect 105228 5800 109316 5828
rect 105228 5788 105234 5800
rect 109310 5788 109316 5800
rect 109368 5788 109374 5840
rect 283374 5788 283380 5840
rect 283432 5828 283438 5840
rect 285950 5828 285956 5840
rect 283432 5800 285956 5828
rect 283432 5788 283438 5800
rect 285950 5788 285956 5800
rect 286008 5788 286014 5840
rect 292574 5788 292580 5840
rect 292632 5828 292638 5840
rect 295518 5828 295524 5840
rect 292632 5800 295524 5828
rect 292632 5788 292638 5800
rect 295518 5788 295524 5800
rect 295576 5788 295582 5840
rect 306282 5788 306288 5840
rect 306340 5828 306346 5840
rect 307938 5828 307944 5840
rect 306340 5800 307944 5828
rect 306340 5788 306346 5800
rect 307938 5788 307944 5800
rect 307996 5788 308002 5840
rect 321186 5788 321192 5840
rect 321244 5828 321250 5840
rect 324130 5828 324136 5840
rect 321244 5800 324136 5828
rect 321244 5788 321250 5800
rect 324130 5788 324136 5800
rect 324188 5788 324194 5840
rect 324590 5788 324596 5840
rect 324648 5828 324654 5840
rect 327166 5828 327172 5840
rect 324648 5800 327172 5828
rect 324648 5788 324654 5800
rect 327166 5788 327172 5800
rect 327224 5788 327230 5840
rect 333790 5788 333796 5840
rect 333848 5828 333854 5840
rect 336642 5828 336648 5840
rect 333848 5800 336648 5828
rect 333848 5788 333854 5800
rect 336642 5788 336648 5800
rect 336700 5788 336706 5840
rect 339494 5788 339500 5840
rect 339552 5828 339558 5840
rect 342254 5828 342260 5840
rect 339552 5800 342260 5828
rect 339552 5788 339558 5800
rect 342254 5788 342260 5800
rect 342312 5788 342318 5840
rect 349798 5788 349804 5840
rect 349856 5828 349862 5840
rect 352282 5828 352288 5840
rect 349856 5800 352288 5828
rect 349856 5788 349862 5800
rect 352282 5788 352288 5800
rect 352340 5788 352346 5840
rect 353202 5788 353208 5840
rect 353260 5828 353266 5840
rect 355502 5828 355508 5840
rect 353260 5800 355508 5828
rect 353260 5788 353266 5800
rect 355502 5788 355508 5800
rect 355560 5788 355566 5840
rect 368106 5788 368112 5840
rect 368164 5828 368170 5840
rect 371050 5828 371056 5840
rect 368164 5800 371056 5828
rect 368164 5788 368170 5800
rect 371050 5788 371056 5800
rect 371108 5788 371114 5840
rect 373810 5788 373816 5840
rect 373868 5828 373874 5840
rect 376662 5828 376668 5840
rect 373868 5800 376668 5828
rect 373868 5788 373874 5800
rect 376662 5788 376668 5800
rect 376720 5788 376726 5840
rect 380710 5788 380716 5840
rect 380768 5828 380774 5840
rect 382274 5828 382280 5840
rect 380768 5800 382280 5828
rect 380768 5788 380774 5800
rect 382274 5788 382280 5800
rect 382332 5788 382338 5840
rect 383010 5788 383016 5840
rect 383068 5828 383074 5840
rect 386138 5828 386144 5840
rect 383068 5800 386144 5828
rect 383068 5788 383074 5800
rect 386138 5788 386144 5800
rect 386196 5788 386202 5840
rect 387610 5788 387616 5840
rect 387668 5828 387674 5840
rect 389174 5828 389180 5840
rect 387668 5800 389180 5828
rect 387668 5788 387674 5800
rect 389174 5788 389180 5800
rect 389232 5788 389238 5840
rect 392118 5788 392124 5840
rect 392176 5828 392182 5840
rect 395338 5828 395344 5840
rect 392176 5800 395344 5828
rect 392176 5788 392182 5800
rect 395338 5788 395344 5800
rect 395396 5788 395402 5840
rect 396718 5788 396724 5840
rect 396776 5828 396782 5840
rect 399846 5828 399852 5840
rect 396776 5800 399852 5828
rect 396776 5788 396782 5800
rect 399846 5788 399852 5800
rect 399904 5788 399910 5840
rect 401318 5788 401324 5840
rect 401376 5828 401382 5840
rect 403894 5828 403900 5840
rect 401376 5800 403900 5828
rect 401376 5788 401382 5800
rect 403894 5788 403900 5800
rect 403952 5788 403958 5840
rect 408218 5788 408224 5840
rect 408276 5828 408282 5840
rect 410426 5828 410432 5840
rect 408276 5800 410432 5828
rect 408276 5788 408282 5800
rect 410426 5788 410432 5800
rect 410484 5788 410490 5840
rect 420822 5788 420828 5840
rect 420880 5828 420886 5840
rect 423306 5828 423312 5840
rect 420880 5800 423312 5828
rect 420880 5788 420886 5800
rect 423306 5788 423312 5800
rect 423364 5788 423370 5840
rect 425330 5788 425336 5840
rect 425388 5828 425394 5840
rect 427814 5828 427820 5840
rect 425388 5800 427820 5828
rect 425388 5788 425394 5800
rect 427814 5788 427820 5800
rect 427872 5788 427878 5840
rect 441430 5788 441436 5840
rect 441488 5828 441494 5840
rect 443454 5828 443460 5840
rect 441488 5800 443460 5828
rect 441488 5788 441494 5800
rect 443454 5788 443460 5800
rect 443512 5788 443518 5840
rect 443730 5788 443736 5840
rect 443788 5828 443794 5840
rect 445846 5828 445852 5840
rect 443788 5800 445852 5828
rect 443788 5788 443794 5800
rect 445846 5788 445852 5800
rect 445904 5788 445910 5840
rect 445938 5788 445944 5840
rect 445996 5828 446002 5840
rect 448606 5828 448612 5840
rect 445996 5800 448612 5828
rect 445996 5788 446002 5800
rect 448606 5788 448612 5800
rect 448664 5788 448670 5840
rect 456334 5788 456340 5840
rect 456392 5828 456398 5840
rect 458634 5828 458640 5840
rect 456392 5800 458640 5828
rect 456392 5788 456398 5800
rect 458634 5788 458640 5800
rect 458692 5788 458698 5840
rect 12526 5720 12532 5772
rect 12584 5760 12590 5772
rect 13814 5760 13820 5772
rect 12584 5732 13820 5760
rect 12584 5720 12590 5732
rect 13814 5720 13820 5732
rect 13872 5720 13878 5772
rect 94498 5720 94504 5772
rect 94556 5760 94562 5772
rect 99006 5760 99012 5772
rect 94556 5732 99012 5760
rect 94556 5720 94562 5732
rect 99006 5720 99012 5732
rect 99064 5720 99070 5772
rect 107562 5720 107568 5772
rect 107620 5760 107626 5772
rect 111610 5760 111616 5772
rect 107620 5732 111616 5760
rect 107620 5720 107626 5732
rect 111610 5720 111616 5732
rect 111668 5720 111674 5772
rect 113542 5720 113548 5772
rect 113600 5760 113606 5772
rect 117314 5760 117320 5772
rect 113600 5732 117320 5760
rect 113600 5720 113606 5732
rect 117314 5720 117320 5732
rect 117372 5720 117378 5772
rect 118234 5720 118240 5772
rect 118292 5760 118298 5772
rect 121914 5760 121920 5772
rect 118292 5732 121920 5760
rect 118292 5720 118298 5732
rect 121914 5720 121920 5732
rect 121972 5720 121978 5772
rect 123018 5720 123024 5772
rect 123076 5760 123082 5772
rect 126514 5760 126520 5772
rect 123076 5732 126520 5760
rect 123076 5720 123082 5732
rect 126514 5720 126520 5732
rect 126572 5720 126578 5772
rect 143258 5720 143264 5772
rect 143316 5760 143322 5772
rect 145926 5760 145932 5772
rect 143316 5732 145932 5760
rect 143316 5720 143322 5732
rect 145926 5720 145932 5732
rect 145984 5720 145990 5772
rect 152734 5720 152740 5772
rect 152792 5760 152798 5772
rect 155126 5760 155132 5772
rect 152792 5732 155132 5760
rect 152792 5720 152798 5732
rect 155126 5720 155132 5732
rect 155184 5720 155190 5772
rect 277670 5720 277676 5772
rect 277728 5760 277734 5772
rect 280062 5760 280068 5772
rect 277728 5732 280068 5760
rect 277728 5720 277734 5732
rect 280062 5720 280068 5732
rect 280120 5720 280126 5772
rect 282178 5720 282184 5772
rect 282236 5760 282242 5772
rect 284754 5760 284760 5772
rect 282236 5732 284760 5760
rect 282236 5720 282242 5732
rect 284754 5720 284760 5732
rect 284812 5720 284818 5772
rect 291378 5720 291384 5772
rect 291436 5760 291442 5772
rect 294322 5760 294328 5772
rect 291436 5732 294328 5760
rect 291436 5720 291442 5732
rect 294322 5720 294328 5732
rect 294380 5720 294386 5772
rect 297082 5720 297088 5772
rect 297140 5760 297146 5772
rect 300302 5760 300308 5772
rect 297140 5732 300308 5760
rect 297140 5720 297146 5732
rect 300302 5720 300308 5732
rect 300360 5720 300366 5772
rect 302878 5720 302884 5772
rect 302936 5760 302942 5772
rect 306190 5760 306196 5772
rect 302936 5732 306196 5760
rect 302936 5720 302942 5732
rect 306190 5720 306196 5732
rect 306248 5720 306254 5772
rect 308582 5720 308588 5772
rect 308640 5760 308646 5772
rect 311802 5760 311808 5772
rect 308640 5732 311808 5760
rect 308640 5720 308646 5732
rect 311802 5720 311808 5732
rect 311860 5720 311866 5772
rect 317690 5720 317696 5772
rect 317748 5760 317754 5772
rect 321462 5760 321468 5772
rect 317748 5732 321468 5760
rect 317748 5720 317754 5732
rect 321462 5720 321468 5732
rect 321520 5720 321526 5772
rect 332594 5720 332600 5772
rect 332652 5760 332658 5772
rect 335814 5760 335820 5772
rect 332652 5732 335820 5760
rect 332652 5720 332658 5732
rect 335814 5720 335820 5732
rect 335872 5720 335878 5772
rect 338298 5720 338304 5772
rect 338356 5760 338362 5772
rect 340874 5760 340880 5772
rect 338356 5732 340880 5760
rect 338356 5720 338362 5732
rect 340874 5720 340880 5732
rect 340932 5720 340938 5772
rect 365806 5720 365812 5772
rect 365864 5760 365870 5772
rect 368658 5760 368664 5772
rect 365864 5732 368664 5760
rect 365864 5720 365870 5732
rect 368658 5720 368664 5732
rect 368716 5720 368722 5772
rect 399018 5720 399024 5772
rect 399076 5760 399082 5772
rect 401594 5760 401600 5772
rect 399076 5732 401600 5760
rect 399076 5720 399082 5732
rect 401594 5720 401600 5732
rect 401652 5720 401658 5772
rect 12434 5652 12440 5704
rect 12492 5692 12498 5704
rect 15378 5692 15384 5704
rect 12492 5664 15384 5692
rect 12492 5652 12498 5664
rect 15378 5652 15384 5664
rect 15436 5652 15442 5704
rect 18690 5652 18696 5704
rect 18748 5692 18754 5704
rect 21082 5692 21088 5704
rect 18748 5664 21088 5692
rect 18748 5652 18754 5664
rect 21082 5652 21088 5664
rect 21140 5652 21146 5704
rect 22094 5652 22100 5704
rect 22152 5692 22158 5704
rect 24578 5692 24584 5704
rect 22152 5664 24584 5692
rect 22152 5652 22158 5664
rect 24578 5652 24584 5664
rect 24636 5652 24642 5704
rect 28994 5652 29000 5704
rect 29052 5692 29058 5704
rect 31386 5692 31392 5704
rect 29052 5664 31392 5692
rect 29052 5652 29058 5664
rect 31386 5652 31392 5664
rect 31444 5652 31450 5704
rect 79042 5652 79048 5704
rect 79100 5692 79106 5704
rect 84102 5692 84108 5704
rect 79100 5664 84108 5692
rect 79100 5652 79106 5664
rect 84102 5652 84108 5664
rect 84160 5652 84166 5704
rect 96890 5652 96896 5704
rect 96948 5692 96954 5704
rect 101306 5692 101312 5704
rect 96948 5664 101312 5692
rect 96948 5652 96954 5664
rect 101306 5652 101312 5664
rect 101364 5652 101370 5704
rect 101582 5652 101588 5704
rect 101640 5692 101646 5704
rect 105906 5692 105912 5704
rect 101640 5664 105912 5692
rect 101640 5652 101646 5664
rect 105906 5652 105912 5664
rect 105964 5652 105970 5704
rect 109954 5652 109960 5704
rect 110012 5692 110018 5704
rect 113910 5692 113916 5704
rect 110012 5664 113916 5692
rect 110012 5652 110018 5664
rect 113910 5652 113916 5664
rect 113968 5652 113974 5704
rect 114738 5652 114744 5704
rect 114796 5692 114802 5704
rect 118418 5692 118424 5704
rect 114796 5664 118424 5692
rect 114796 5652 114802 5664
rect 118418 5652 118424 5664
rect 118476 5652 118482 5704
rect 125410 5652 125416 5704
rect 125468 5692 125474 5704
rect 128722 5692 128728 5704
rect 125468 5664 128728 5692
rect 125468 5652 125474 5664
rect 128722 5652 128728 5664
rect 128780 5652 128786 5704
rect 128998 5652 129004 5704
rect 129056 5692 129062 5704
rect 132218 5692 132224 5704
rect 129056 5664 132224 5692
rect 129056 5652 129062 5664
rect 132218 5652 132224 5664
rect 132276 5652 132282 5704
rect 132586 5652 132592 5704
rect 132644 5692 132650 5704
rect 135622 5692 135628 5704
rect 132644 5664 135628 5692
rect 132644 5652 132650 5664
rect 135622 5652 135628 5664
rect 135680 5652 135686 5704
rect 136082 5652 136088 5704
rect 136140 5692 136146 5704
rect 139118 5692 139124 5704
rect 136140 5664 139124 5692
rect 136140 5652 136146 5664
rect 139118 5652 139124 5664
rect 139176 5652 139182 5704
rect 139670 5652 139676 5704
rect 139728 5692 139734 5704
rect 142522 5692 142528 5704
rect 139728 5664 142528 5692
rect 139728 5652 139734 5664
rect 142522 5652 142528 5664
rect 142580 5652 142586 5704
rect 144454 5652 144460 5704
rect 144512 5692 144518 5704
rect 147122 5692 147128 5704
rect 144512 5664 147128 5692
rect 144512 5652 144518 5664
rect 147122 5652 147128 5664
rect 147180 5652 147186 5704
rect 148042 5652 148048 5704
rect 148100 5692 148106 5704
rect 150526 5692 150532 5704
rect 148100 5664 150532 5692
rect 148100 5652 148106 5664
rect 150526 5652 150532 5664
rect 150584 5652 150590 5704
rect 157518 5652 157524 5704
rect 157576 5692 157582 5704
rect 159726 5692 159732 5704
rect 157576 5664 159732 5692
rect 157576 5652 157582 5664
rect 159726 5652 159732 5664
rect 159784 5652 159790 5704
rect 171778 5652 171784 5704
rect 171836 5692 171842 5704
rect 173434 5692 173440 5704
rect 171836 5664 173440 5692
rect 171836 5652 171842 5664
rect 173434 5652 173440 5664
rect 173492 5652 173498 5704
rect 184750 5652 184756 5704
rect 184808 5692 184814 5704
rect 186038 5692 186044 5704
rect 184808 5664 186044 5692
rect 184808 5652 184814 5664
rect 186038 5652 186044 5664
rect 186096 5652 186102 5704
rect 248966 5652 248972 5704
rect 249024 5692 249030 5704
rect 250346 5692 250352 5704
rect 249024 5664 250352 5692
rect 249024 5652 249030 5664
rect 250346 5652 250352 5664
rect 250404 5652 250410 5704
rect 266170 5652 266176 5704
rect 266228 5692 266234 5704
rect 268102 5692 268108 5704
rect 266228 5664 268108 5692
rect 266228 5652 266234 5664
rect 268102 5652 268108 5664
rect 268160 5652 268166 5704
rect 276474 5652 276480 5704
rect 276532 5692 276538 5704
rect 278866 5692 278872 5704
rect 276532 5664 278872 5692
rect 276532 5652 276538 5664
rect 278866 5652 278872 5664
rect 278924 5652 278930 5704
rect 281074 5652 281080 5704
rect 281132 5692 281138 5704
rect 283650 5692 283656 5704
rect 281132 5664 283656 5692
rect 281132 5652 281138 5664
rect 283650 5652 283656 5664
rect 283708 5652 283714 5704
rect 286778 5652 286784 5704
rect 286836 5692 286842 5704
rect 289538 5692 289544 5704
rect 286836 5664 289544 5692
rect 286836 5652 286842 5664
rect 289538 5652 289544 5664
rect 289596 5652 289602 5704
rect 290274 5652 290280 5704
rect 290332 5692 290338 5704
rect 293126 5692 293132 5704
rect 290332 5664 293132 5692
rect 290332 5652 290338 5664
rect 293126 5652 293132 5664
rect 293184 5652 293190 5704
rect 295978 5652 295984 5704
rect 296036 5692 296042 5704
rect 299106 5692 299112 5704
rect 296036 5664 299112 5692
rect 296036 5652 296042 5664
rect 299106 5652 299112 5664
rect 299164 5652 299170 5704
rect 300578 5652 300584 5704
rect 300636 5692 300642 5704
rect 303522 5692 303528 5704
rect 300636 5664 303528 5692
rect 300636 5652 300642 5664
rect 303522 5652 303528 5664
rect 303580 5652 303586 5704
rect 311986 5652 311992 5704
rect 312044 5692 312050 5704
rect 315758 5692 315764 5704
rect 312044 5664 315764 5692
rect 312044 5652 312050 5664
rect 315758 5652 315764 5664
rect 315816 5652 315822 5704
rect 319990 5652 319996 5704
rect 320048 5692 320054 5704
rect 322014 5692 322020 5704
rect 320048 5664 322020 5692
rect 320048 5652 320054 5664
rect 322014 5652 322020 5664
rect 322072 5652 322078 5704
rect 327994 5652 328000 5704
rect 328052 5692 328058 5704
rect 330110 5692 330116 5704
rect 328052 5664 330116 5692
rect 328052 5652 328058 5664
rect 330110 5652 330116 5664
rect 330168 5652 330174 5704
rect 337194 5652 337200 5704
rect 337252 5692 337258 5704
rect 339494 5692 339500 5704
rect 337252 5664 339500 5692
rect 337252 5652 337258 5664
rect 339494 5652 339500 5664
rect 339552 5652 339558 5704
rect 345198 5652 345204 5704
rect 345256 5692 345262 5704
rect 347774 5692 347780 5704
rect 345256 5664 347780 5692
rect 345256 5652 345262 5664
rect 347774 5652 347780 5664
rect 347832 5652 347838 5704
rect 348602 5652 348608 5704
rect 348660 5692 348666 5704
rect 351086 5692 351092 5704
rect 348660 5664 351092 5692
rect 348660 5652 348666 5664
rect 351086 5652 351092 5664
rect 351144 5652 351150 5704
rect 354398 5652 354404 5704
rect 354456 5692 354462 5704
rect 357250 5692 357256 5704
rect 354456 5664 357256 5692
rect 354456 5652 354462 5664
rect 357250 5652 357256 5664
rect 357308 5652 357314 5704
rect 358906 5652 358912 5704
rect 358964 5692 358970 5704
rect 361574 5692 361580 5704
rect 358964 5664 361580 5692
rect 358964 5652 358970 5664
rect 361574 5652 361580 5664
rect 361632 5652 361638 5704
rect 363506 5652 363512 5704
rect 363564 5692 363570 5704
rect 366542 5692 366548 5704
rect 363564 5664 366548 5692
rect 363564 5652 363570 5664
rect 366542 5652 366548 5664
rect 366600 5652 366606 5704
rect 372706 5652 372712 5704
rect 372764 5692 372770 5704
rect 375834 5692 375840 5704
rect 372764 5664 375840 5692
rect 372764 5652 372770 5664
rect 375834 5652 375840 5664
rect 375892 5652 375898 5704
rect 376110 5652 376116 5704
rect 376168 5692 376174 5704
rect 379422 5692 379428 5704
rect 376168 5664 379428 5692
rect 376168 5652 376174 5664
rect 379422 5652 379428 5664
rect 379480 5652 379486 5704
rect 386414 5652 386420 5704
rect 386472 5692 386478 5704
rect 389634 5692 389640 5704
rect 386472 5664 389640 5692
rect 386472 5652 386478 5664
rect 389634 5652 389640 5664
rect 389692 5652 389698 5704
rect 395614 5652 395620 5704
rect 395672 5692 395678 5704
rect 398742 5692 398748 5704
rect 395672 5664 398748 5692
rect 395672 5652 395678 5664
rect 398742 5652 398748 5664
rect 398800 5652 398806 5704
rect 405918 5652 405924 5704
rect 405976 5692 405982 5704
rect 409414 5692 409420 5704
rect 405976 5664 409420 5692
rect 405976 5652 405982 5664
rect 409414 5652 409420 5664
rect 409472 5652 409478 5704
rect 413922 5652 413928 5704
rect 413980 5692 413986 5704
rect 416682 5692 416688 5704
rect 413980 5664 416688 5692
rect 413980 5652 413986 5664
rect 416682 5652 416688 5664
rect 416740 5652 416746 5704
rect 428826 5652 428832 5704
rect 428884 5692 428890 5704
rect 430574 5692 430580 5704
rect 428884 5664 430580 5692
rect 428884 5652 428890 5664
rect 430574 5652 430580 5664
rect 430632 5652 430638 5704
rect 444834 5652 444840 5704
rect 444892 5692 444898 5704
rect 448054 5692 448060 5704
rect 444892 5664 448060 5692
rect 444892 5652 444898 5664
rect 448054 5652 448060 5664
rect 448112 5652 448118 5704
rect 457438 5652 457444 5704
rect 457496 5692 457502 5704
rect 459554 5692 459560 5704
rect 457496 5664 459560 5692
rect 457496 5652 457502 5664
rect 459554 5652 459560 5664
rect 459612 5652 459618 5704
rect 471146 5652 471152 5704
rect 471204 5692 471210 5704
rect 473354 5692 473360 5704
rect 471204 5664 473360 5692
rect 471204 5652 471210 5664
rect 473354 5652 473360 5664
rect 473412 5652 473418 5704
rect 488350 5652 488356 5704
rect 488408 5692 488414 5704
rect 490374 5692 490380 5704
rect 488408 5664 490380 5692
rect 488408 5652 488414 5664
rect 490374 5652 490380 5664
rect 490432 5652 490438 5704
rect 13814 5584 13820 5636
rect 13872 5624 13878 5636
rect 16574 5624 16580 5636
rect 13872 5596 16580 5624
rect 13872 5584 13878 5596
rect 16574 5584 16580 5596
rect 16632 5584 16638 5636
rect 19426 5584 19432 5636
rect 19484 5624 19490 5636
rect 22278 5624 22284 5636
rect 19484 5596 22284 5624
rect 19484 5584 19490 5596
rect 22278 5584 22284 5596
rect 22336 5584 22342 5636
rect 28258 5584 28264 5636
rect 28316 5624 28322 5636
rect 30282 5624 30288 5636
rect 28316 5596 30288 5624
rect 28316 5584 28322 5596
rect 30282 5584 30288 5596
rect 30340 5584 30346 5636
rect 31754 5584 31760 5636
rect 31812 5624 31818 5636
rect 33134 5624 33140 5636
rect 31812 5596 33140 5624
rect 31812 5584 31818 5596
rect 33134 5584 33140 5596
rect 33192 5584 33198 5636
rect 34514 5584 34520 5636
rect 34572 5624 34578 5636
rect 37182 5624 37188 5636
rect 34572 5596 37188 5624
rect 34572 5584 34578 5596
rect 37182 5584 37188 5596
rect 37240 5584 37246 5636
rect 37642 5584 37648 5636
rect 37700 5624 37706 5636
rect 39482 5624 39488 5636
rect 37700 5596 39488 5624
rect 37700 5584 37706 5596
rect 39482 5584 39488 5596
rect 39540 5584 39546 5636
rect 44174 5584 44180 5636
rect 44232 5624 44238 5636
rect 46290 5624 46296 5636
rect 44232 5596 46296 5624
rect 44232 5584 44238 5596
rect 46290 5584 46296 5596
rect 46348 5584 46354 5636
rect 81434 5584 81440 5636
rect 81492 5624 81498 5636
rect 86402 5624 86408 5636
rect 81492 5596 86408 5624
rect 81492 5584 81498 5596
rect 86402 5584 86408 5596
rect 86460 5584 86466 5636
rect 87322 5584 87328 5636
rect 87380 5624 87386 5636
rect 92106 5624 92112 5636
rect 87380 5596 92112 5624
rect 87380 5584 87386 5596
rect 92106 5584 92112 5596
rect 92164 5584 92170 5636
rect 98086 5584 98092 5636
rect 98144 5624 98150 5636
rect 102410 5624 102416 5636
rect 98144 5596 102416 5624
rect 98144 5584 98150 5596
rect 102410 5584 102416 5596
rect 102468 5584 102474 5636
rect 103974 5584 103980 5636
rect 104032 5624 104038 5636
rect 108114 5624 108120 5636
rect 104032 5596 108120 5624
rect 104032 5584 104038 5596
rect 108114 5584 108120 5596
rect 108172 5584 108178 5636
rect 108666 5584 108672 5636
rect 108724 5624 108730 5636
rect 112714 5624 112720 5636
rect 108724 5596 112720 5624
rect 108724 5584 108730 5596
rect 112714 5584 112720 5596
rect 112772 5584 112778 5636
rect 115934 5584 115940 5636
rect 115992 5624 115998 5636
rect 119614 5624 119620 5636
rect 115992 5596 119620 5624
rect 115992 5584 115998 5596
rect 119614 5584 119620 5596
rect 119672 5584 119678 5636
rect 124214 5584 124220 5636
rect 124272 5624 124278 5636
rect 127618 5624 127624 5636
rect 124272 5596 127624 5624
rect 124272 5584 124278 5596
rect 127618 5584 127624 5596
rect 127676 5584 127682 5636
rect 127802 5584 127808 5636
rect 127860 5624 127866 5636
rect 131022 5624 131028 5636
rect 127860 5596 131028 5624
rect 127860 5584 127866 5596
rect 131022 5584 131028 5596
rect 131080 5584 131086 5636
rect 131390 5584 131396 5636
rect 131448 5624 131454 5636
rect 134518 5624 134524 5636
rect 131448 5596 134524 5624
rect 131448 5584 131454 5596
rect 134518 5584 134524 5596
rect 134576 5584 134582 5636
rect 134886 5584 134892 5636
rect 134944 5624 134950 5636
rect 137922 5624 137928 5636
rect 134944 5596 137928 5624
rect 134944 5584 134950 5596
rect 137922 5584 137928 5596
rect 137980 5584 137986 5636
rect 138474 5584 138480 5636
rect 138532 5624 138538 5636
rect 141326 5624 141332 5636
rect 138532 5596 141332 5624
rect 138532 5584 138538 5596
rect 141326 5584 141332 5596
rect 141384 5584 141390 5636
rect 142062 5584 142068 5636
rect 142120 5624 142126 5636
rect 144822 5624 144828 5636
rect 142120 5596 144828 5624
rect 142120 5584 142126 5596
rect 144822 5584 144828 5596
rect 144880 5584 144886 5636
rect 146846 5584 146852 5636
rect 146904 5624 146910 5636
rect 149422 5624 149428 5636
rect 146904 5596 149428 5624
rect 146904 5584 146910 5596
rect 149422 5584 149428 5596
rect 149480 5584 149486 5636
rect 150434 5584 150440 5636
rect 150492 5624 150498 5636
rect 152826 5624 152832 5636
rect 150492 5596 152832 5624
rect 150492 5584 150498 5596
rect 152826 5584 152832 5596
rect 152884 5584 152890 5636
rect 155126 5584 155132 5636
rect 155184 5624 155190 5636
rect 157426 5624 157432 5636
rect 155184 5596 157432 5624
rect 155184 5584 155190 5596
rect 157426 5584 157432 5596
rect 157484 5584 157490 5636
rect 158714 5584 158720 5636
rect 158772 5624 158778 5636
rect 160830 5624 160836 5636
rect 158772 5596 160836 5624
rect 158772 5584 158778 5596
rect 160830 5584 160836 5596
rect 160888 5584 160894 5636
rect 163498 5584 163504 5636
rect 163556 5624 163562 5636
rect 165430 5624 165436 5636
rect 163556 5596 165436 5624
rect 163556 5584 163562 5596
rect 165430 5584 165436 5596
rect 165488 5584 165494 5636
rect 165890 5584 165896 5636
rect 165948 5624 165954 5636
rect 167730 5624 167736 5636
rect 165948 5596 167736 5624
rect 165948 5584 165954 5596
rect 167730 5584 167736 5596
rect 167788 5584 167794 5636
rect 168190 5584 168196 5636
rect 168248 5624 168254 5636
rect 170030 5624 170036 5636
rect 168248 5596 170036 5624
rect 168248 5584 168254 5596
rect 170030 5584 170036 5596
rect 170088 5584 170094 5636
rect 170582 5584 170588 5636
rect 170640 5624 170646 5636
rect 172330 5624 172336 5636
rect 170640 5596 172336 5624
rect 170640 5584 170646 5596
rect 172330 5584 172336 5596
rect 172388 5584 172394 5636
rect 174170 5584 174176 5636
rect 174228 5624 174234 5636
rect 175734 5624 175740 5636
rect 174228 5596 175740 5624
rect 174228 5584 174234 5596
rect 175734 5584 175740 5596
rect 175792 5584 175798 5636
rect 176562 5584 176568 5636
rect 176620 5624 176626 5636
rect 178034 5624 178040 5636
rect 176620 5596 178040 5624
rect 176620 5584 176626 5596
rect 178034 5584 178040 5596
rect 178092 5584 178098 5636
rect 178954 5584 178960 5636
rect 179012 5624 179018 5636
rect 180334 5624 180340 5636
rect 179012 5596 180340 5624
rect 179012 5584 179018 5596
rect 180334 5584 180340 5596
rect 180392 5584 180398 5636
rect 181530 5584 181536 5636
rect 181588 5624 181594 5636
rect 182634 5624 182640 5636
rect 181588 5596 182640 5624
rect 181588 5584 181594 5596
rect 182634 5584 182640 5596
rect 182692 5584 182698 5636
rect 247862 5584 247868 5636
rect 247920 5624 247926 5636
rect 249150 5624 249156 5636
rect 247920 5596 249156 5624
rect 247920 5584 247926 5596
rect 249150 5584 249156 5596
rect 249208 5584 249214 5636
rect 251266 5584 251272 5636
rect 251324 5624 251330 5636
rect 252646 5624 252652 5636
rect 251324 5596 252652 5624
rect 251324 5584 251330 5596
rect 252646 5584 252652 5596
rect 252704 5584 252710 5636
rect 253566 5584 253572 5636
rect 253624 5624 253630 5636
rect 255038 5624 255044 5636
rect 253624 5596 255044 5624
rect 253624 5584 253630 5596
rect 255038 5584 255044 5596
rect 255096 5584 255102 5636
rect 255866 5584 255872 5636
rect 255924 5624 255930 5636
rect 257430 5624 257436 5636
rect 255924 5596 257436 5624
rect 255924 5584 255930 5596
rect 257430 5584 257436 5596
rect 257488 5584 257494 5636
rect 258166 5584 258172 5636
rect 258224 5624 258230 5636
rect 259822 5624 259828 5636
rect 258224 5596 259828 5624
rect 258224 5584 258230 5596
rect 259822 5584 259828 5596
rect 259880 5584 259886 5636
rect 260466 5584 260472 5636
rect 260524 5624 260530 5636
rect 262214 5624 262220 5636
rect 260524 5596 262220 5624
rect 260524 5584 260530 5596
rect 262214 5584 262220 5596
rect 262272 5584 262278 5636
rect 262766 5584 262772 5636
rect 262824 5624 262830 5636
rect 264606 5624 264612 5636
rect 262824 5596 264612 5624
rect 262824 5584 262830 5596
rect 264606 5584 264612 5596
rect 264664 5584 264670 5636
rect 265066 5584 265072 5636
rect 265124 5624 265130 5636
rect 266998 5624 267004 5636
rect 265124 5596 267004 5624
rect 265124 5584 265130 5596
rect 266998 5584 267004 5596
rect 267056 5584 267062 5636
rect 268470 5584 268476 5636
rect 268528 5624 268534 5636
rect 270494 5624 270500 5636
rect 268528 5596 270500 5624
rect 268528 5584 268534 5596
rect 270494 5584 270500 5596
rect 270552 5584 270558 5636
rect 273070 5584 273076 5636
rect 273128 5624 273134 5636
rect 275278 5624 275284 5636
rect 273128 5596 275284 5624
rect 273128 5584 273134 5596
rect 275278 5584 275284 5596
rect 275336 5584 275342 5636
rect 275370 5584 275376 5636
rect 275428 5624 275434 5636
rect 277670 5624 277676 5636
rect 275428 5596 277676 5624
rect 275428 5584 275434 5596
rect 277670 5584 277676 5596
rect 277728 5584 277734 5636
rect 279970 5584 279976 5636
rect 280028 5624 280034 5636
rect 282454 5624 282460 5636
rect 280028 5596 282460 5624
rect 280028 5584 280034 5596
rect 282454 5584 282460 5596
rect 282512 5584 282518 5636
rect 285674 5584 285680 5636
rect 285732 5624 285738 5636
rect 288342 5624 288348 5636
rect 285732 5596 288348 5624
rect 285732 5584 285738 5596
rect 288342 5584 288348 5596
rect 288400 5584 288406 5636
rect 289078 5584 289084 5636
rect 289136 5624 289142 5636
rect 291930 5624 291936 5636
rect 289136 5596 291936 5624
rect 289136 5584 289142 5596
rect 291930 5584 291936 5596
rect 291988 5584 291994 5636
rect 294782 5584 294788 5636
rect 294840 5624 294846 5636
rect 297910 5624 297916 5636
rect 294840 5596 297916 5624
rect 294840 5584 294846 5596
rect 297910 5584 297916 5596
rect 297968 5584 297974 5636
rect 299382 5584 299388 5636
rect 299440 5624 299446 5636
rect 301038 5624 301044 5636
rect 299440 5596 301044 5624
rect 299440 5584 299446 5596
rect 301038 5584 301044 5596
rect 301096 5584 301102 5636
rect 301682 5584 301688 5636
rect 301740 5624 301746 5636
rect 304902 5624 304908 5636
rect 301740 5596 304908 5624
rect 301740 5584 301746 5596
rect 304902 5584 304908 5596
rect 304960 5584 304966 5636
rect 305086 5584 305092 5636
rect 305144 5624 305150 5636
rect 308582 5624 308588 5636
rect 305144 5596 308588 5624
rect 305144 5584 305150 5596
rect 308582 5584 308588 5596
rect 308640 5584 308646 5636
rect 310882 5584 310888 5636
rect 310940 5624 310946 5636
rect 314562 5624 314568 5636
rect 310940 5596 314568 5624
rect 310940 5584 310946 5596
rect 314562 5584 314568 5596
rect 314620 5584 314626 5636
rect 315390 5584 315396 5636
rect 315448 5624 315454 5636
rect 317690 5624 317696 5636
rect 315448 5596 317696 5624
rect 315448 5584 315454 5596
rect 317690 5584 317696 5596
rect 317748 5584 317754 5636
rect 318886 5584 318892 5636
rect 318944 5624 318950 5636
rect 322842 5624 322848 5636
rect 318944 5596 322848 5624
rect 318944 5584 318950 5596
rect 322842 5584 322848 5596
rect 322900 5584 322906 5636
rect 325694 5584 325700 5636
rect 325752 5624 325758 5636
rect 329742 5624 329748 5636
rect 325752 5596 329748 5624
rect 325752 5584 325758 5596
rect 329742 5584 329748 5596
rect 329800 5584 329806 5636
rect 330294 5584 330300 5636
rect 330352 5624 330358 5636
rect 332594 5624 332600 5636
rect 330352 5596 332600 5624
rect 330352 5584 330358 5596
rect 332594 5584 332600 5596
rect 332652 5584 332658 5636
rect 334894 5584 334900 5636
rect 334952 5624 334958 5636
rect 337286 5624 337292 5636
rect 334952 5596 337292 5624
rect 334952 5584 334958 5596
rect 337286 5584 337292 5596
rect 337344 5584 337350 5636
rect 346394 5584 346400 5636
rect 346452 5624 346458 5636
rect 349154 5624 349160 5636
rect 346452 5596 349160 5624
rect 346452 5584 346458 5596
rect 349154 5584 349160 5596
rect 349212 5584 349218 5636
rect 352098 5584 352104 5636
rect 352156 5624 352162 5636
rect 355594 5624 355600 5636
rect 352156 5596 355600 5624
rect 352156 5584 352162 5596
rect 355594 5584 355600 5596
rect 355652 5584 355658 5636
rect 357802 5584 357808 5636
rect 357860 5624 357866 5636
rect 360562 5624 360568 5636
rect 357860 5596 360568 5624
rect 357860 5584 357866 5596
rect 360562 5584 360568 5596
rect 360620 5584 360626 5636
rect 364702 5584 364708 5636
rect 364760 5624 364766 5636
rect 367462 5624 367468 5636
rect 364760 5596 367468 5624
rect 364760 5584 364766 5596
rect 367462 5584 367468 5596
rect 367520 5584 367526 5636
rect 377306 5584 377312 5636
rect 377364 5624 377370 5636
rect 380434 5624 380440 5636
rect 377364 5596 380440 5624
rect 377364 5584 377370 5596
rect 380434 5584 380440 5596
rect 380492 5584 380498 5636
rect 384114 5584 384120 5636
rect 384172 5624 384178 5636
rect 387334 5624 387340 5636
rect 384172 5596 387340 5624
rect 384172 5584 384178 5596
rect 387334 5584 387340 5596
rect 387392 5584 387398 5636
rect 389910 5584 389916 5636
rect 389968 5624 389974 5636
rect 391934 5624 391940 5636
rect 389968 5596 391940 5624
rect 389968 5584 389974 5596
rect 391934 5584 391940 5596
rect 391992 5584 391998 5636
rect 393314 5584 393320 5636
rect 393372 5624 393378 5636
rect 396534 5624 396540 5636
rect 393372 5596 396540 5624
rect 393372 5584 393378 5596
rect 396534 5584 396540 5596
rect 396592 5584 396598 5636
rect 397914 5584 397920 5636
rect 397972 5624 397978 5636
rect 400490 5624 400496 5636
rect 397972 5596 400496 5624
rect 397972 5584 397978 5596
rect 400490 5584 400496 5596
rect 400548 5584 400554 5636
rect 403618 5584 403624 5636
rect 403676 5624 403682 5636
rect 407022 5624 407028 5636
rect 403676 5596 407028 5624
rect 403676 5584 403682 5596
rect 407022 5584 407028 5596
rect 407080 5584 407086 5636
rect 409322 5584 409328 5636
rect 409380 5624 409386 5636
rect 411254 5624 411260 5636
rect 409380 5596 411260 5624
rect 409380 5584 409386 5596
rect 411254 5584 411260 5596
rect 411312 5584 411318 5636
rect 412726 5584 412732 5636
rect 412784 5624 412790 5636
rect 416498 5624 416504 5636
rect 412784 5596 416504 5624
rect 412784 5584 412790 5596
rect 416498 5584 416504 5596
rect 416556 5584 416562 5636
rect 423122 5584 423128 5636
rect 423180 5624 423186 5636
rect 426250 5624 426256 5636
rect 423180 5596 426256 5624
rect 423180 5584 423186 5596
rect 426250 5584 426256 5596
rect 426308 5584 426314 5636
rect 432230 5584 432236 5636
rect 432288 5624 432294 5636
rect 436002 5624 436008 5636
rect 432288 5596 436008 5624
rect 432288 5584 432294 5596
rect 436002 5584 436008 5596
rect 436060 5584 436066 5636
rect 451734 5584 451740 5636
rect 451792 5624 451798 5636
rect 455322 5624 455328 5636
rect 451792 5596 455328 5624
rect 451792 5584 451798 5596
rect 455322 5584 455328 5596
rect 455380 5584 455386 5636
rect 518158 5584 518164 5636
rect 518216 5624 518222 5636
rect 521562 5624 521568 5636
rect 518216 5596 521568 5624
rect 518216 5584 518222 5596
rect 521562 5584 521568 5596
rect 521620 5584 521626 5636
rect 547874 5584 547880 5636
rect 547932 5624 547938 5636
rect 551922 5624 551928 5636
rect 547932 5596 551928 5624
rect 547932 5584 547938 5596
rect 551922 5584 551928 5596
rect 551980 5584 551986 5636
rect 15194 5516 15200 5568
rect 15252 5556 15258 5568
rect 17678 5556 17684 5568
rect 15252 5528 17684 5556
rect 15252 5516 15258 5528
rect 17678 5516 17684 5528
rect 17736 5516 17742 5568
rect 18322 5516 18328 5568
rect 18380 5556 18386 5568
rect 19978 5556 19984 5568
rect 18380 5528 19984 5556
rect 18380 5516 18386 5528
rect 19978 5516 19984 5528
rect 20036 5516 20042 5568
rect 20806 5516 20812 5568
rect 20864 5556 20870 5568
rect 23382 5556 23388 5568
rect 20864 5528 23388 5556
rect 20864 5516 20870 5528
rect 23382 5516 23388 5528
rect 23440 5516 23446 5568
rect 23474 5516 23480 5568
rect 23532 5556 23538 5568
rect 25682 5556 25688 5568
rect 23532 5528 25688 5556
rect 23532 5516 23538 5528
rect 25682 5516 25688 5528
rect 25740 5516 25746 5568
rect 26602 5516 26608 5568
rect 26660 5556 26666 5568
rect 29178 5556 29184 5568
rect 26660 5528 29184 5556
rect 26660 5516 26666 5528
rect 29178 5516 29184 5528
rect 29236 5516 29242 5568
rect 30374 5516 30380 5568
rect 30432 5556 30438 5568
rect 32582 5556 32588 5568
rect 30432 5528 32588 5556
rect 30432 5516 30438 5528
rect 32582 5516 32588 5528
rect 32640 5516 32646 5568
rect 36722 5516 36728 5568
rect 36780 5556 36786 5568
rect 38286 5556 38292 5568
rect 36780 5528 38292 5556
rect 36780 5516 36786 5528
rect 38286 5516 38292 5528
rect 38344 5516 38350 5568
rect 40034 5516 40040 5568
rect 40092 5556 40098 5568
rect 41414 5556 41420 5568
rect 40092 5528 41420 5556
rect 40092 5516 40098 5528
rect 41414 5516 41420 5528
rect 41472 5516 41478 5568
rect 42794 5516 42800 5568
rect 42852 5556 42858 5568
rect 45186 5556 45192 5568
rect 42852 5528 45192 5556
rect 42852 5516 42858 5528
rect 45186 5516 45192 5528
rect 45244 5516 45250 5568
rect 53834 5516 53840 5568
rect 53892 5556 53898 5568
rect 55490 5556 55496 5568
rect 53892 5528 55496 5556
rect 53892 5516 53898 5528
rect 55490 5516 55496 5528
rect 55548 5516 55554 5568
rect 62114 5516 62120 5568
rect 62172 5556 62178 5568
rect 63494 5556 63500 5568
rect 62172 5528 63500 5556
rect 62172 5516 62178 5528
rect 63494 5516 63500 5528
rect 63552 5516 63558 5568
rect 71866 5516 71872 5568
rect 71924 5556 71930 5568
rect 77202 5556 77208 5568
rect 71924 5528 77208 5556
rect 71924 5516 71930 5528
rect 77202 5516 77208 5528
rect 77260 5516 77266 5568
rect 80238 5516 80244 5568
rect 80296 5556 80302 5568
rect 85206 5556 85212 5568
rect 80296 5528 85212 5556
rect 80296 5516 80302 5528
rect 85206 5516 85212 5528
rect 85264 5516 85270 5568
rect 89714 5516 89720 5568
rect 89772 5556 89778 5568
rect 94406 5556 94412 5568
rect 89772 5528 94412 5556
rect 89772 5516 89778 5528
rect 94406 5516 94412 5528
rect 94464 5516 94470 5568
rect 95694 5516 95700 5568
rect 95752 5556 95758 5568
rect 100110 5556 100116 5568
rect 95752 5528 100116 5556
rect 95752 5516 95758 5528
rect 100110 5516 100116 5528
rect 100168 5516 100174 5568
rect 100478 5516 100484 5568
rect 100536 5556 100542 5568
rect 104710 5556 104716 5568
rect 100536 5528 104716 5556
rect 100536 5516 100542 5528
rect 104710 5516 104716 5528
rect 104768 5516 104774 5568
rect 106366 5516 106372 5568
rect 106424 5556 106430 5568
rect 110414 5556 110420 5568
rect 106424 5528 110420 5556
rect 106424 5516 106430 5528
rect 110414 5516 110420 5528
rect 110472 5516 110478 5568
rect 111150 5516 111156 5568
rect 111208 5556 111214 5568
rect 115014 5556 115020 5568
rect 111208 5528 115020 5556
rect 111208 5516 111214 5528
rect 115014 5516 115020 5528
rect 115072 5516 115078 5568
rect 117130 5516 117136 5568
rect 117188 5556 117194 5568
rect 120718 5556 120724 5568
rect 117188 5528 120724 5556
rect 117188 5516 117194 5528
rect 120718 5516 120724 5528
rect 120776 5516 120782 5568
rect 121822 5516 121828 5568
rect 121880 5556 121886 5568
rect 125318 5556 125324 5568
rect 121880 5528 125324 5556
rect 121880 5516 121886 5528
rect 125318 5516 125324 5528
rect 125376 5516 125382 5568
rect 126606 5516 126612 5568
rect 126664 5556 126670 5568
rect 129918 5556 129924 5568
rect 126664 5528 129924 5556
rect 126664 5516 126670 5528
rect 129918 5516 129924 5528
rect 129976 5516 129982 5568
rect 130194 5516 130200 5568
rect 130252 5556 130258 5568
rect 133322 5556 133328 5568
rect 130252 5528 133328 5556
rect 130252 5516 130258 5528
rect 133322 5516 133328 5528
rect 133380 5516 133386 5568
rect 133782 5516 133788 5568
rect 133840 5556 133846 5568
rect 136818 5556 136824 5568
rect 133840 5528 136824 5556
rect 133840 5516 133846 5528
rect 136818 5516 136824 5528
rect 136876 5516 136882 5568
rect 137278 5516 137284 5568
rect 137336 5556 137342 5568
rect 140222 5556 140228 5568
rect 137336 5528 140228 5556
rect 137336 5516 137342 5528
rect 140222 5516 140228 5528
rect 140280 5516 140286 5568
rect 140866 5516 140872 5568
rect 140924 5556 140930 5568
rect 143626 5556 143632 5568
rect 140924 5528 143632 5556
rect 140924 5516 140930 5528
rect 143626 5516 143632 5528
rect 143684 5516 143690 5568
rect 145650 5516 145656 5568
rect 145708 5556 145714 5568
rect 148226 5556 148232 5568
rect 145708 5528 148232 5556
rect 145708 5516 145714 5528
rect 148226 5516 148232 5528
rect 148284 5516 148290 5568
rect 149238 5516 149244 5568
rect 149296 5556 149302 5568
rect 151630 5556 151636 5568
rect 149296 5528 151636 5556
rect 149296 5516 149302 5528
rect 151630 5516 151636 5528
rect 151688 5516 151694 5568
rect 153930 5516 153936 5568
rect 153988 5556 153994 5568
rect 156230 5556 156236 5568
rect 153988 5528 156236 5556
rect 153988 5516 153994 5528
rect 156230 5516 156236 5528
rect 156288 5516 156294 5568
rect 156322 5516 156328 5568
rect 156380 5556 156386 5568
rect 158530 5556 158536 5568
rect 156380 5528 158536 5556
rect 156380 5516 156386 5528
rect 158530 5516 158536 5528
rect 158588 5516 158594 5568
rect 159910 5516 159916 5568
rect 159968 5556 159974 5568
rect 161934 5556 161940 5568
rect 159968 5528 161940 5556
rect 159968 5516 159974 5528
rect 161934 5516 161940 5528
rect 161992 5516 161998 5568
rect 162302 5516 162308 5568
rect 162360 5556 162366 5568
rect 164234 5556 164240 5568
rect 162360 5528 164240 5556
rect 162360 5516 162366 5528
rect 164234 5516 164240 5528
rect 164292 5516 164298 5568
rect 164694 5516 164700 5568
rect 164752 5556 164758 5568
rect 166534 5556 166540 5568
rect 164752 5528 166540 5556
rect 164752 5516 164758 5528
rect 166534 5516 166540 5528
rect 166592 5516 166598 5568
rect 167086 5516 167092 5568
rect 167144 5556 167150 5568
rect 168834 5556 168840 5568
rect 167144 5528 168840 5556
rect 167144 5516 167150 5528
rect 168834 5516 168840 5528
rect 168892 5516 168898 5568
rect 169386 5516 169392 5568
rect 169444 5556 169450 5568
rect 171134 5556 171140 5568
rect 169444 5528 171140 5556
rect 169444 5516 169450 5528
rect 171134 5516 171140 5528
rect 171192 5516 171198 5568
rect 172974 5516 172980 5568
rect 173032 5556 173038 5568
rect 174538 5556 174544 5568
rect 173032 5528 174544 5556
rect 173032 5516 173038 5528
rect 174538 5516 174544 5528
rect 174596 5516 174602 5568
rect 175366 5516 175372 5568
rect 175424 5556 175430 5568
rect 176838 5556 176844 5568
rect 175424 5528 176844 5556
rect 175424 5516 175430 5528
rect 176838 5516 176844 5528
rect 176896 5516 176902 5568
rect 177758 5516 177764 5568
rect 177816 5556 177822 5568
rect 179138 5556 179144 5568
rect 177816 5528 179144 5556
rect 177816 5516 177822 5528
rect 179138 5516 179144 5528
rect 179196 5516 179202 5568
rect 180150 5516 180156 5568
rect 180208 5556 180214 5568
rect 181438 5556 181444 5568
rect 180208 5528 181444 5556
rect 180208 5516 180214 5528
rect 181438 5516 181444 5528
rect 181496 5516 181502 5568
rect 182542 5516 182548 5568
rect 182600 5556 182606 5568
rect 183738 5556 183744 5568
rect 182600 5528 183744 5556
rect 182600 5516 182606 5528
rect 183738 5516 183744 5528
rect 183796 5516 183802 5568
rect 186038 5516 186044 5568
rect 186096 5556 186102 5568
rect 187142 5556 187148 5568
rect 186096 5528 187148 5556
rect 186096 5516 186102 5528
rect 187142 5516 187148 5528
rect 187200 5516 187206 5568
rect 187234 5516 187240 5568
rect 187292 5556 187298 5568
rect 188338 5556 188344 5568
rect 187292 5528 188344 5556
rect 187292 5516 187298 5528
rect 188338 5516 188344 5528
rect 188396 5516 188402 5568
rect 188430 5516 188436 5568
rect 188488 5556 188494 5568
rect 189442 5556 189448 5568
rect 188488 5528 189448 5556
rect 188488 5516 188494 5528
rect 189442 5516 189448 5528
rect 189500 5516 189506 5568
rect 189626 5516 189632 5568
rect 189684 5556 189690 5568
rect 190638 5556 190644 5568
rect 189684 5528 190644 5556
rect 189684 5516 189690 5528
rect 190638 5516 190644 5528
rect 190696 5516 190702 5568
rect 194410 5516 194416 5568
rect 194468 5556 194474 5568
rect 195146 5556 195152 5568
rect 194468 5528 195152 5556
rect 194468 5516 194474 5528
rect 195146 5516 195152 5528
rect 195204 5516 195210 5568
rect 196802 5516 196808 5568
rect 196860 5556 196866 5568
rect 197446 5556 197452 5568
rect 196860 5528 197452 5556
rect 196860 5516 196866 5528
rect 197446 5516 197452 5528
rect 197504 5516 197510 5568
rect 202690 5516 202696 5568
rect 202748 5556 202754 5568
rect 203242 5556 203248 5568
rect 202748 5528 203248 5556
rect 202748 5516 202754 5528
rect 203242 5516 203248 5528
rect 203300 5516 203306 5568
rect 232958 5516 232964 5568
rect 233016 5556 233022 5568
rect 233694 5556 233700 5568
rect 233016 5528 233700 5556
rect 233016 5516 233022 5528
rect 233694 5516 233700 5528
rect 233752 5516 233758 5568
rect 238662 5516 238668 5568
rect 238720 5556 238726 5568
rect 239582 5556 239588 5568
rect 238720 5528 239588 5556
rect 238720 5516 238726 5528
rect 239582 5516 239588 5528
rect 239640 5516 239646 5568
rect 239858 5516 239864 5568
rect 239916 5556 239922 5568
rect 240778 5556 240784 5568
rect 239916 5528 240784 5556
rect 239916 5516 239922 5528
rect 240778 5516 240784 5528
rect 240836 5516 240842 5568
rect 240962 5516 240968 5568
rect 241020 5556 241026 5568
rect 241974 5556 241980 5568
rect 241020 5528 241980 5556
rect 241020 5516 241026 5528
rect 241974 5516 241980 5528
rect 242032 5516 242038 5568
rect 242158 5516 242164 5568
rect 242216 5556 242222 5568
rect 243170 5556 243176 5568
rect 242216 5528 243176 5556
rect 242216 5516 242222 5528
rect 243170 5516 243176 5528
rect 243228 5516 243234 5568
rect 243262 5516 243268 5568
rect 243320 5556 243326 5568
rect 244366 5556 244372 5568
rect 243320 5528 244372 5556
rect 243320 5516 243326 5528
rect 244366 5516 244372 5528
rect 244424 5516 244430 5568
rect 245562 5516 245568 5568
rect 245620 5556 245626 5568
rect 246666 5556 246672 5568
rect 245620 5528 246672 5556
rect 245620 5516 245626 5528
rect 246666 5516 246672 5528
rect 246724 5516 246730 5568
rect 246758 5516 246764 5568
rect 246816 5556 246822 5568
rect 247954 5556 247960 5568
rect 246816 5528 247960 5556
rect 246816 5516 246822 5528
rect 247954 5516 247960 5528
rect 248012 5516 248018 5568
rect 250162 5516 250168 5568
rect 250220 5556 250226 5568
rect 251450 5556 251456 5568
rect 250220 5528 251456 5556
rect 250220 5516 250226 5528
rect 251450 5516 251456 5528
rect 251508 5516 251514 5568
rect 252462 5516 252468 5568
rect 252520 5556 252526 5568
rect 253842 5556 253848 5568
rect 252520 5528 253848 5556
rect 252520 5516 252526 5528
rect 253842 5516 253848 5528
rect 253900 5516 253906 5568
rect 254762 5516 254768 5568
rect 254820 5556 254826 5568
rect 256234 5556 256240 5568
rect 254820 5528 256240 5556
rect 254820 5516 254826 5528
rect 256234 5516 256240 5528
rect 256292 5516 256298 5568
rect 257062 5516 257068 5568
rect 257120 5556 257126 5568
rect 258626 5556 258632 5568
rect 257120 5528 258632 5556
rect 257120 5516 257126 5528
rect 258626 5516 258632 5528
rect 258684 5516 258690 5568
rect 259362 5516 259368 5568
rect 259420 5556 259426 5568
rect 261018 5556 261024 5568
rect 259420 5528 261024 5556
rect 259420 5516 259426 5528
rect 261018 5516 261024 5528
rect 261076 5516 261082 5568
rect 261570 5516 261576 5568
rect 261628 5556 261634 5568
rect 263410 5556 263416 5568
rect 261628 5528 263416 5556
rect 261628 5516 261634 5528
rect 263410 5516 263416 5528
rect 263468 5516 263474 5568
rect 263870 5516 263876 5568
rect 263928 5556 263934 5568
rect 265802 5556 265808 5568
rect 263928 5528 265808 5556
rect 263928 5516 263934 5528
rect 265802 5516 265808 5528
rect 265860 5516 265866 5568
rect 267366 5516 267372 5568
rect 267424 5556 267430 5568
rect 269298 5556 269304 5568
rect 267424 5528 269304 5556
rect 267424 5516 267430 5528
rect 269298 5516 269304 5528
rect 269356 5516 269362 5568
rect 269666 5516 269672 5568
rect 269724 5556 269730 5568
rect 271690 5556 271696 5568
rect 269724 5528 271696 5556
rect 269724 5516 269730 5528
rect 271690 5516 271696 5528
rect 271748 5516 271754 5568
rect 271874 5516 271880 5568
rect 271932 5556 271938 5568
rect 274082 5556 274088 5568
rect 271932 5528 274088 5556
rect 271932 5516 271938 5528
rect 274082 5516 274088 5528
rect 274140 5516 274146 5568
rect 274174 5516 274180 5568
rect 274232 5556 274238 5568
rect 276474 5556 276480 5568
rect 274232 5528 276480 5556
rect 274232 5516 274238 5528
rect 276474 5516 276480 5528
rect 276532 5516 276538 5568
rect 278774 5516 278780 5568
rect 278832 5556 278838 5568
rect 281258 5556 281264 5568
rect 278832 5528 281264 5556
rect 278832 5516 278838 5528
rect 281258 5516 281264 5528
rect 281316 5516 281322 5568
rect 284478 5516 284484 5568
rect 284536 5556 284542 5568
rect 287146 5556 287152 5568
rect 284536 5528 287152 5556
rect 284536 5516 284542 5528
rect 287146 5516 287152 5528
rect 287204 5516 287210 5568
rect 287974 5516 287980 5568
rect 288032 5556 288038 5568
rect 290734 5556 290740 5568
rect 288032 5528 290740 5556
rect 288032 5516 288038 5528
rect 290734 5516 290740 5528
rect 290792 5516 290798 5568
rect 293678 5516 293684 5568
rect 293736 5556 293742 5568
rect 296622 5556 296628 5568
rect 293736 5528 296628 5556
rect 293736 5516 293742 5528
rect 296622 5516 296628 5528
rect 296680 5516 296686 5568
rect 298278 5516 298284 5568
rect 298336 5556 298342 5568
rect 301406 5556 301412 5568
rect 298336 5528 301412 5556
rect 298336 5516 298342 5528
rect 301406 5516 301412 5528
rect 301464 5516 301470 5568
rect 303982 5516 303988 5568
rect 304040 5556 304046 5568
rect 307478 5556 307484 5568
rect 304040 5528 307484 5556
rect 304040 5516 304046 5528
rect 307478 5516 307484 5528
rect 307536 5516 307542 5568
rect 309686 5516 309692 5568
rect 309744 5556 309750 5568
rect 313182 5556 313188 5568
rect 309744 5528 313188 5556
rect 309744 5516 309750 5528
rect 313182 5516 313188 5528
rect 313240 5516 313246 5568
rect 314286 5516 314292 5568
rect 314344 5556 314350 5568
rect 316494 5556 316500 5568
rect 314344 5528 316500 5556
rect 314344 5516 314350 5528
rect 316494 5516 316500 5528
rect 316552 5516 316558 5568
rect 316586 5516 316592 5568
rect 316644 5556 316650 5568
rect 320082 5556 320088 5568
rect 316644 5528 320088 5556
rect 316644 5516 316650 5528
rect 320082 5516 320088 5528
rect 320140 5516 320146 5568
rect 323486 5516 323492 5568
rect 323544 5556 323550 5568
rect 326522 5556 326528 5568
rect 323544 5528 326528 5556
rect 323544 5516 323550 5528
rect 326522 5516 326528 5528
rect 326580 5516 326586 5568
rect 326890 5516 326896 5568
rect 326948 5556 326954 5568
rect 329006 5556 329012 5568
rect 326948 5528 329012 5556
rect 326948 5516 326954 5528
rect 329006 5516 329012 5528
rect 329064 5516 329070 5568
rect 329190 5516 329196 5568
rect 329248 5556 329254 5568
rect 331306 5556 331312 5568
rect 329248 5528 331312 5556
rect 329248 5516 329254 5528
rect 331306 5516 331312 5528
rect 331364 5516 331370 5568
rect 336090 5516 336096 5568
rect 336148 5556 336154 5568
rect 338298 5556 338304 5568
rect 336148 5528 338304 5556
rect 336148 5516 336154 5528
rect 338298 5516 338304 5528
rect 338356 5516 338362 5568
rect 344094 5516 344100 5568
rect 344152 5556 344158 5568
rect 346854 5556 346860 5568
rect 344152 5528 346860 5556
rect 344152 5516 344158 5528
rect 346854 5516 346860 5528
rect 346912 5516 346918 5568
rect 347498 5516 347504 5568
rect 347556 5556 347562 5568
rect 349982 5556 349988 5568
rect 347556 5528 349988 5556
rect 347556 5516 347562 5528
rect 349982 5516 349988 5528
rect 350040 5516 350046 5568
rect 356698 5516 356704 5568
rect 356756 5556 356762 5568
rect 359366 5556 359372 5568
rect 356756 5528 359372 5556
rect 356756 5516 356762 5528
rect 359366 5516 359372 5528
rect 359424 5516 359430 5568
rect 362402 5516 362408 5568
rect 362460 5556 362466 5568
rect 365622 5556 365628 5568
rect 362460 5528 365628 5556
rect 362460 5516 362466 5528
rect 365622 5516 365628 5528
rect 365680 5516 365686 5568
rect 367002 5516 367008 5568
rect 367060 5556 367066 5568
rect 369762 5556 369768 5568
rect 367060 5528 369768 5556
rect 367060 5516 367066 5528
rect 369762 5516 369768 5528
rect 369820 5516 369826 5568
rect 371510 5516 371516 5568
rect 371568 5556 371574 5568
rect 374730 5556 374736 5568
rect 371568 5528 374736 5556
rect 371568 5516 371574 5528
rect 374730 5516 374736 5528
rect 374788 5516 374794 5568
rect 375006 5516 375012 5568
rect 375064 5556 375070 5568
rect 378042 5556 378048 5568
rect 375064 5528 378048 5556
rect 375064 5516 375070 5528
rect 378042 5516 378048 5528
rect 378100 5516 378106 5568
rect 378410 5516 378416 5568
rect 378468 5556 378474 5568
rect 380894 5556 380900 5568
rect 378468 5528 380900 5556
rect 378468 5516 378474 5528
rect 380894 5516 380900 5528
rect 380952 5516 380958 5568
rect 381814 5516 381820 5568
rect 381872 5556 381878 5568
rect 384942 5556 384948 5568
rect 381872 5528 384948 5556
rect 381872 5516 381878 5528
rect 384942 5516 384948 5528
rect 385000 5516 385006 5568
rect 385310 5516 385316 5568
rect 385368 5556 385374 5568
rect 388530 5556 388536 5568
rect 385368 5528 388536 5556
rect 385368 5516 385374 5528
rect 388530 5516 388536 5528
rect 388588 5516 388594 5568
rect 391014 5516 391020 5568
rect 391072 5556 391078 5568
rect 393590 5556 393596 5568
rect 391072 5528 393596 5556
rect 391072 5516 391078 5528
rect 393590 5516 393596 5528
rect 393648 5516 393654 5568
rect 394418 5516 394424 5568
rect 394476 5556 394482 5568
rect 396718 5556 396724 5568
rect 394476 5528 396724 5556
rect 394476 5516 394482 5528
rect 396718 5516 396724 5528
rect 396776 5516 396782 5568
rect 400214 5516 400220 5568
rect 400272 5556 400278 5568
rect 404078 5556 404084 5568
rect 400272 5528 404084 5556
rect 400272 5516 400278 5528
rect 404078 5516 404084 5528
rect 404136 5516 404142 5568
rect 404722 5516 404728 5568
rect 404780 5556 404786 5568
rect 408402 5556 408408 5568
rect 404780 5528 408408 5556
rect 404780 5516 404786 5528
rect 408402 5516 408408 5528
rect 408460 5516 408466 5568
rect 411622 5516 411628 5568
rect 411680 5556 411686 5568
rect 414658 5556 414664 5568
rect 411680 5528 414664 5556
rect 411680 5516 411686 5528
rect 414658 5516 414664 5528
rect 414716 5516 414722 5568
rect 417326 5516 417332 5568
rect 417384 5556 417390 5568
rect 419810 5556 419816 5568
rect 417384 5528 419816 5556
rect 417384 5516 417390 5528
rect 419810 5516 419816 5528
rect 419868 5516 419874 5568
rect 424226 5516 424232 5568
rect 424284 5556 424290 5568
rect 426434 5556 426440 5568
rect 424284 5528 426440 5556
rect 424284 5516 424290 5528
rect 426434 5516 426440 5528
rect 426492 5516 426498 5568
rect 426526 5516 426532 5568
rect 426584 5556 426590 5568
rect 429194 5556 429200 5568
rect 426584 5528 429200 5556
rect 426584 5516 426590 5528
rect 429194 5516 429200 5528
rect 429252 5516 429258 5568
rect 429930 5516 429936 5568
rect 429988 5556 429994 5568
rect 432690 5556 432696 5568
rect 429988 5528 432696 5556
rect 429988 5516 429994 5528
rect 432690 5516 432696 5528
rect 432748 5516 432754 5568
rect 435634 5516 435640 5568
rect 435692 5556 435698 5568
rect 438578 5556 438584 5568
rect 435692 5528 438584 5556
rect 435692 5516 435698 5528
rect 438578 5516 438584 5528
rect 438636 5516 438642 5568
rect 439130 5516 439136 5568
rect 439188 5556 439194 5568
rect 442074 5556 442080 5568
rect 439188 5528 442080 5556
rect 439188 5516 439194 5528
rect 442074 5516 442080 5528
rect 442132 5516 442138 5568
rect 452838 5516 452844 5568
rect 452896 5556 452902 5568
rect 455414 5556 455420 5568
rect 452896 5528 455420 5556
rect 452896 5516 452902 5528
rect 455414 5516 455420 5528
rect 455472 5516 455478 5568
rect 459738 5516 459744 5568
rect 459796 5556 459802 5568
rect 463602 5556 463608 5568
rect 459796 5528 463608 5556
rect 459796 5516 459802 5528
rect 463602 5516 463608 5528
rect 463660 5516 463666 5568
rect 472342 5516 472348 5568
rect 472400 5556 472406 5568
rect 474734 5556 474740 5568
rect 472400 5528 474740 5556
rect 472400 5516 472406 5528
rect 474734 5516 474740 5528
rect 474792 5516 474798 5568
rect 503254 5516 503260 5568
rect 503312 5556 503318 5568
rect 506290 5556 506296 5568
rect 503312 5528 506296 5556
rect 503312 5516 503318 5528
rect 506290 5516 506296 5528
rect 506348 5516 506354 5568
rect 532970 5516 532976 5568
rect 533028 5556 533034 5568
rect 535454 5556 535460 5568
rect 533028 5528 535460 5556
rect 533028 5516 533034 5528
rect 535454 5516 535460 5528
rect 535512 5516 535518 5568
rect 549070 5516 549076 5568
rect 549128 5556 549134 5568
rect 550726 5556 550732 5568
rect 549128 5528 550732 5556
rect 549128 5516 549134 5528
rect 550726 5516 550732 5528
rect 550784 5516 550790 5568
rect 1104 5466 582820 5488
rect 1104 5414 36822 5466
rect 36874 5414 36886 5466
rect 36938 5414 36950 5466
rect 37002 5414 37014 5466
rect 37066 5414 37078 5466
rect 37130 5414 37142 5466
rect 37194 5414 37206 5466
rect 37258 5414 37270 5466
rect 37322 5414 37334 5466
rect 37386 5414 72822 5466
rect 72874 5414 72886 5466
rect 72938 5414 72950 5466
rect 73002 5414 73014 5466
rect 73066 5414 73078 5466
rect 73130 5414 73142 5466
rect 73194 5414 73206 5466
rect 73258 5414 73270 5466
rect 73322 5414 73334 5466
rect 73386 5414 108822 5466
rect 108874 5414 108886 5466
rect 108938 5414 108950 5466
rect 109002 5414 109014 5466
rect 109066 5414 109078 5466
rect 109130 5414 109142 5466
rect 109194 5414 109206 5466
rect 109258 5414 109270 5466
rect 109322 5414 109334 5466
rect 109386 5414 144822 5466
rect 144874 5414 144886 5466
rect 144938 5414 144950 5466
rect 145002 5414 145014 5466
rect 145066 5414 145078 5466
rect 145130 5414 145142 5466
rect 145194 5414 145206 5466
rect 145258 5414 145270 5466
rect 145322 5414 145334 5466
rect 145386 5414 180822 5466
rect 180874 5414 180886 5466
rect 180938 5414 180950 5466
rect 181002 5414 181014 5466
rect 181066 5414 181078 5466
rect 181130 5414 181142 5466
rect 181194 5414 181206 5466
rect 181258 5414 181270 5466
rect 181322 5414 181334 5466
rect 181386 5414 216822 5466
rect 216874 5414 216886 5466
rect 216938 5414 216950 5466
rect 217002 5414 217014 5466
rect 217066 5414 217078 5466
rect 217130 5414 217142 5466
rect 217194 5414 217206 5466
rect 217258 5414 217270 5466
rect 217322 5414 217334 5466
rect 217386 5414 252822 5466
rect 252874 5414 252886 5466
rect 252938 5414 252950 5466
rect 253002 5414 253014 5466
rect 253066 5414 253078 5466
rect 253130 5414 253142 5466
rect 253194 5414 253206 5466
rect 253258 5414 253270 5466
rect 253322 5414 253334 5466
rect 253386 5414 288822 5466
rect 288874 5414 288886 5466
rect 288938 5414 288950 5466
rect 289002 5414 289014 5466
rect 289066 5414 289078 5466
rect 289130 5414 289142 5466
rect 289194 5414 289206 5466
rect 289258 5414 289270 5466
rect 289322 5414 289334 5466
rect 289386 5414 324822 5466
rect 324874 5414 324886 5466
rect 324938 5414 324950 5466
rect 325002 5414 325014 5466
rect 325066 5414 325078 5466
rect 325130 5414 325142 5466
rect 325194 5414 325206 5466
rect 325258 5414 325270 5466
rect 325322 5414 325334 5466
rect 325386 5414 360822 5466
rect 360874 5414 360886 5466
rect 360938 5414 360950 5466
rect 361002 5414 361014 5466
rect 361066 5414 361078 5466
rect 361130 5414 361142 5466
rect 361194 5414 361206 5466
rect 361258 5414 361270 5466
rect 361322 5414 361334 5466
rect 361386 5414 396822 5466
rect 396874 5414 396886 5466
rect 396938 5414 396950 5466
rect 397002 5414 397014 5466
rect 397066 5414 397078 5466
rect 397130 5414 397142 5466
rect 397194 5414 397206 5466
rect 397258 5414 397270 5466
rect 397322 5414 397334 5466
rect 397386 5414 432822 5466
rect 432874 5414 432886 5466
rect 432938 5414 432950 5466
rect 433002 5414 433014 5466
rect 433066 5414 433078 5466
rect 433130 5414 433142 5466
rect 433194 5414 433206 5466
rect 433258 5414 433270 5466
rect 433322 5414 433334 5466
rect 433386 5414 468822 5466
rect 468874 5414 468886 5466
rect 468938 5414 468950 5466
rect 469002 5414 469014 5466
rect 469066 5414 469078 5466
rect 469130 5414 469142 5466
rect 469194 5414 469206 5466
rect 469258 5414 469270 5466
rect 469322 5414 469334 5466
rect 469386 5414 504822 5466
rect 504874 5414 504886 5466
rect 504938 5414 504950 5466
rect 505002 5414 505014 5466
rect 505066 5414 505078 5466
rect 505130 5414 505142 5466
rect 505194 5414 505206 5466
rect 505258 5414 505270 5466
rect 505322 5414 505334 5466
rect 505386 5414 540822 5466
rect 540874 5414 540886 5466
rect 540938 5414 540950 5466
rect 541002 5414 541014 5466
rect 541066 5414 541078 5466
rect 541130 5414 541142 5466
rect 541194 5414 541206 5466
rect 541258 5414 541270 5466
rect 541322 5414 541334 5466
rect 541386 5414 576822 5466
rect 576874 5414 576886 5466
rect 576938 5414 576950 5466
rect 577002 5414 577014 5466
rect 577066 5414 577078 5466
rect 577130 5414 577142 5466
rect 577194 5414 577206 5466
rect 577258 5414 577270 5466
rect 577322 5414 577334 5466
rect 577386 5414 582820 5466
rect 1104 5392 582820 5414
rect 1104 4922 582820 4944
rect 1104 4870 18822 4922
rect 18874 4870 18886 4922
rect 18938 4870 18950 4922
rect 19002 4870 19014 4922
rect 19066 4870 19078 4922
rect 19130 4870 19142 4922
rect 19194 4870 19206 4922
rect 19258 4870 19270 4922
rect 19322 4870 19334 4922
rect 19386 4870 54822 4922
rect 54874 4870 54886 4922
rect 54938 4870 54950 4922
rect 55002 4870 55014 4922
rect 55066 4870 55078 4922
rect 55130 4870 55142 4922
rect 55194 4870 55206 4922
rect 55258 4870 55270 4922
rect 55322 4870 55334 4922
rect 55386 4870 90822 4922
rect 90874 4870 90886 4922
rect 90938 4870 90950 4922
rect 91002 4870 91014 4922
rect 91066 4870 91078 4922
rect 91130 4870 91142 4922
rect 91194 4870 91206 4922
rect 91258 4870 91270 4922
rect 91322 4870 91334 4922
rect 91386 4870 126822 4922
rect 126874 4870 126886 4922
rect 126938 4870 126950 4922
rect 127002 4870 127014 4922
rect 127066 4870 127078 4922
rect 127130 4870 127142 4922
rect 127194 4870 127206 4922
rect 127258 4870 127270 4922
rect 127322 4870 127334 4922
rect 127386 4870 162822 4922
rect 162874 4870 162886 4922
rect 162938 4870 162950 4922
rect 163002 4870 163014 4922
rect 163066 4870 163078 4922
rect 163130 4870 163142 4922
rect 163194 4870 163206 4922
rect 163258 4870 163270 4922
rect 163322 4870 163334 4922
rect 163386 4870 198822 4922
rect 198874 4870 198886 4922
rect 198938 4870 198950 4922
rect 199002 4870 199014 4922
rect 199066 4870 199078 4922
rect 199130 4870 199142 4922
rect 199194 4870 199206 4922
rect 199258 4870 199270 4922
rect 199322 4870 199334 4922
rect 199386 4870 234822 4922
rect 234874 4870 234886 4922
rect 234938 4870 234950 4922
rect 235002 4870 235014 4922
rect 235066 4870 235078 4922
rect 235130 4870 235142 4922
rect 235194 4870 235206 4922
rect 235258 4870 235270 4922
rect 235322 4870 235334 4922
rect 235386 4870 270822 4922
rect 270874 4870 270886 4922
rect 270938 4870 270950 4922
rect 271002 4870 271014 4922
rect 271066 4870 271078 4922
rect 271130 4870 271142 4922
rect 271194 4870 271206 4922
rect 271258 4870 271270 4922
rect 271322 4870 271334 4922
rect 271386 4870 306822 4922
rect 306874 4870 306886 4922
rect 306938 4870 306950 4922
rect 307002 4870 307014 4922
rect 307066 4870 307078 4922
rect 307130 4870 307142 4922
rect 307194 4870 307206 4922
rect 307258 4870 307270 4922
rect 307322 4870 307334 4922
rect 307386 4870 342822 4922
rect 342874 4870 342886 4922
rect 342938 4870 342950 4922
rect 343002 4870 343014 4922
rect 343066 4870 343078 4922
rect 343130 4870 343142 4922
rect 343194 4870 343206 4922
rect 343258 4870 343270 4922
rect 343322 4870 343334 4922
rect 343386 4870 378822 4922
rect 378874 4870 378886 4922
rect 378938 4870 378950 4922
rect 379002 4870 379014 4922
rect 379066 4870 379078 4922
rect 379130 4870 379142 4922
rect 379194 4870 379206 4922
rect 379258 4870 379270 4922
rect 379322 4870 379334 4922
rect 379386 4870 414822 4922
rect 414874 4870 414886 4922
rect 414938 4870 414950 4922
rect 415002 4870 415014 4922
rect 415066 4870 415078 4922
rect 415130 4870 415142 4922
rect 415194 4870 415206 4922
rect 415258 4870 415270 4922
rect 415322 4870 415334 4922
rect 415386 4870 450822 4922
rect 450874 4870 450886 4922
rect 450938 4870 450950 4922
rect 451002 4870 451014 4922
rect 451066 4870 451078 4922
rect 451130 4870 451142 4922
rect 451194 4870 451206 4922
rect 451258 4870 451270 4922
rect 451322 4870 451334 4922
rect 451386 4870 486822 4922
rect 486874 4870 486886 4922
rect 486938 4870 486950 4922
rect 487002 4870 487014 4922
rect 487066 4870 487078 4922
rect 487130 4870 487142 4922
rect 487194 4870 487206 4922
rect 487258 4870 487270 4922
rect 487322 4870 487334 4922
rect 487386 4870 522822 4922
rect 522874 4870 522886 4922
rect 522938 4870 522950 4922
rect 523002 4870 523014 4922
rect 523066 4870 523078 4922
rect 523130 4870 523142 4922
rect 523194 4870 523206 4922
rect 523258 4870 523270 4922
rect 523322 4870 523334 4922
rect 523386 4870 558822 4922
rect 558874 4870 558886 4922
rect 558938 4870 558950 4922
rect 559002 4870 559014 4922
rect 559066 4870 559078 4922
rect 559130 4870 559142 4922
rect 559194 4870 559206 4922
rect 559258 4870 559270 4922
rect 559322 4870 559334 4922
rect 559386 4870 582820 4922
rect 1104 4848 582820 4870
rect 1104 4378 582820 4400
rect 1104 4326 36822 4378
rect 36874 4326 36886 4378
rect 36938 4326 36950 4378
rect 37002 4326 37014 4378
rect 37066 4326 37078 4378
rect 37130 4326 37142 4378
rect 37194 4326 37206 4378
rect 37258 4326 37270 4378
rect 37322 4326 37334 4378
rect 37386 4326 72822 4378
rect 72874 4326 72886 4378
rect 72938 4326 72950 4378
rect 73002 4326 73014 4378
rect 73066 4326 73078 4378
rect 73130 4326 73142 4378
rect 73194 4326 73206 4378
rect 73258 4326 73270 4378
rect 73322 4326 73334 4378
rect 73386 4326 108822 4378
rect 108874 4326 108886 4378
rect 108938 4326 108950 4378
rect 109002 4326 109014 4378
rect 109066 4326 109078 4378
rect 109130 4326 109142 4378
rect 109194 4326 109206 4378
rect 109258 4326 109270 4378
rect 109322 4326 109334 4378
rect 109386 4326 144822 4378
rect 144874 4326 144886 4378
rect 144938 4326 144950 4378
rect 145002 4326 145014 4378
rect 145066 4326 145078 4378
rect 145130 4326 145142 4378
rect 145194 4326 145206 4378
rect 145258 4326 145270 4378
rect 145322 4326 145334 4378
rect 145386 4326 180822 4378
rect 180874 4326 180886 4378
rect 180938 4326 180950 4378
rect 181002 4326 181014 4378
rect 181066 4326 181078 4378
rect 181130 4326 181142 4378
rect 181194 4326 181206 4378
rect 181258 4326 181270 4378
rect 181322 4326 181334 4378
rect 181386 4326 216822 4378
rect 216874 4326 216886 4378
rect 216938 4326 216950 4378
rect 217002 4326 217014 4378
rect 217066 4326 217078 4378
rect 217130 4326 217142 4378
rect 217194 4326 217206 4378
rect 217258 4326 217270 4378
rect 217322 4326 217334 4378
rect 217386 4326 252822 4378
rect 252874 4326 252886 4378
rect 252938 4326 252950 4378
rect 253002 4326 253014 4378
rect 253066 4326 253078 4378
rect 253130 4326 253142 4378
rect 253194 4326 253206 4378
rect 253258 4326 253270 4378
rect 253322 4326 253334 4378
rect 253386 4326 288822 4378
rect 288874 4326 288886 4378
rect 288938 4326 288950 4378
rect 289002 4326 289014 4378
rect 289066 4326 289078 4378
rect 289130 4326 289142 4378
rect 289194 4326 289206 4378
rect 289258 4326 289270 4378
rect 289322 4326 289334 4378
rect 289386 4326 324822 4378
rect 324874 4326 324886 4378
rect 324938 4326 324950 4378
rect 325002 4326 325014 4378
rect 325066 4326 325078 4378
rect 325130 4326 325142 4378
rect 325194 4326 325206 4378
rect 325258 4326 325270 4378
rect 325322 4326 325334 4378
rect 325386 4326 360822 4378
rect 360874 4326 360886 4378
rect 360938 4326 360950 4378
rect 361002 4326 361014 4378
rect 361066 4326 361078 4378
rect 361130 4326 361142 4378
rect 361194 4326 361206 4378
rect 361258 4326 361270 4378
rect 361322 4326 361334 4378
rect 361386 4326 396822 4378
rect 396874 4326 396886 4378
rect 396938 4326 396950 4378
rect 397002 4326 397014 4378
rect 397066 4326 397078 4378
rect 397130 4326 397142 4378
rect 397194 4326 397206 4378
rect 397258 4326 397270 4378
rect 397322 4326 397334 4378
rect 397386 4326 432822 4378
rect 432874 4326 432886 4378
rect 432938 4326 432950 4378
rect 433002 4326 433014 4378
rect 433066 4326 433078 4378
rect 433130 4326 433142 4378
rect 433194 4326 433206 4378
rect 433258 4326 433270 4378
rect 433322 4326 433334 4378
rect 433386 4326 468822 4378
rect 468874 4326 468886 4378
rect 468938 4326 468950 4378
rect 469002 4326 469014 4378
rect 469066 4326 469078 4378
rect 469130 4326 469142 4378
rect 469194 4326 469206 4378
rect 469258 4326 469270 4378
rect 469322 4326 469334 4378
rect 469386 4326 504822 4378
rect 504874 4326 504886 4378
rect 504938 4326 504950 4378
rect 505002 4326 505014 4378
rect 505066 4326 505078 4378
rect 505130 4326 505142 4378
rect 505194 4326 505206 4378
rect 505258 4326 505270 4378
rect 505322 4326 505334 4378
rect 505386 4326 540822 4378
rect 540874 4326 540886 4378
rect 540938 4326 540950 4378
rect 541002 4326 541014 4378
rect 541066 4326 541078 4378
rect 541130 4326 541142 4378
rect 541194 4326 541206 4378
rect 541258 4326 541270 4378
rect 541322 4326 541334 4378
rect 541386 4326 576822 4378
rect 576874 4326 576886 4378
rect 576938 4326 576950 4378
rect 577002 4326 577014 4378
rect 577066 4326 577078 4378
rect 577130 4326 577142 4378
rect 577194 4326 577206 4378
rect 577258 4326 577270 4378
rect 577322 4326 577334 4378
rect 577386 4326 582820 4378
rect 1104 4304 582820 4326
rect 51626 4088 51632 4140
rect 51684 4128 51690 4140
rect 57790 4128 57796 4140
rect 51684 4100 57796 4128
rect 51684 4088 51690 4100
rect 57790 4088 57796 4100
rect 57848 4088 57854 4140
rect 70670 4088 70676 4140
rect 70728 4128 70734 4140
rect 76098 4128 76104 4140
rect 70728 4100 76104 4128
rect 70728 4088 70734 4100
rect 76098 4088 76104 4100
rect 76156 4088 76162 4140
rect 355502 4088 355508 4140
rect 355560 4128 355566 4140
rect 358538 4128 358544 4140
rect 355560 4100 358544 4128
rect 355560 4088 355566 4100
rect 358538 4088 358544 4100
rect 358596 4088 358602 4140
rect 366542 4088 366548 4140
rect 366600 4128 366606 4140
rect 369210 4128 369216 4140
rect 366600 4100 369216 4128
rect 366600 4088 366606 4100
rect 369210 4088 369216 4100
rect 369268 4088 369274 4140
rect 371602 4088 371608 4140
rect 371660 4128 371666 4140
rect 375190 4128 375196 4140
rect 371660 4100 375196 4128
rect 371660 4088 371666 4100
rect 375190 4088 375196 4100
rect 375248 4088 375254 4140
rect 375834 4088 375840 4140
rect 375892 4128 375898 4140
rect 378686 4128 378692 4140
rect 375892 4100 378692 4128
rect 375892 4088 375898 4100
rect 378686 4088 378692 4100
rect 378744 4088 378750 4140
rect 380894 4088 380900 4140
rect 380952 4128 380958 4140
rect 384666 4128 384672 4140
rect 380952 4100 384672 4128
rect 380952 4088 380958 4100
rect 384666 4088 384672 4100
rect 384724 4088 384730 4140
rect 391106 4088 391112 4140
rect 391164 4128 391170 4140
rect 395430 4128 395436 4140
rect 391164 4100 395436 4128
rect 391164 4088 391170 4100
rect 395430 4088 395436 4100
rect 395488 4088 395494 4140
rect 404078 4088 404084 4140
rect 404136 4128 404142 4140
rect 407298 4128 407304 4140
rect 404136 4100 407304 4128
rect 404136 4088 404142 4100
rect 407298 4088 407304 4100
rect 407356 4088 407362 4140
rect 408494 4088 408500 4140
rect 408552 4128 408558 4140
rect 414474 4128 414480 4140
rect 408552 4100 414480 4128
rect 408552 4088 408558 4100
rect 414474 4088 414480 4100
rect 414532 4088 414538 4140
rect 448054 4088 448060 4140
rect 448112 4128 448118 4140
rect 453666 4128 453672 4140
rect 448112 4100 453672 4128
rect 448112 4088 448118 4100
rect 453666 4088 453672 4100
rect 453724 4088 453730 4140
rect 539410 4088 539416 4140
rect 539468 4128 539474 4140
rect 540514 4128 540520 4140
rect 539468 4100 540520 4128
rect 539468 4088 539474 4100
rect 540514 4088 540520 4100
rect 540572 4088 540578 4140
rect 546494 4088 546500 4140
rect 546552 4128 546558 4140
rect 548886 4128 548892 4140
rect 546552 4100 548892 4128
rect 546552 4088 546558 4100
rect 548886 4088 548892 4100
rect 548944 4088 548950 4140
rect 568206 4088 568212 4140
rect 568264 4128 568270 4140
rect 571426 4128 571432 4140
rect 568264 4100 571432 4128
rect 568264 4088 568270 4100
rect 571426 4088 571432 4100
rect 571484 4088 571490 4140
rect 566 4020 572 4072
rect 624 4060 630 4072
rect 8570 4060 8576 4072
rect 624 4032 8576 4060
rect 624 4020 630 4032
rect 8570 4020 8576 4032
rect 8628 4020 8634 4072
rect 20714 4020 20720 4072
rect 20772 4060 20778 4072
rect 27522 4060 27528 4072
rect 20772 4032 27528 4060
rect 20772 4020 20778 4032
rect 27522 4020 27528 4032
rect 27580 4020 27586 4072
rect 31478 4020 31484 4072
rect 31536 4060 31542 4072
rect 36722 4060 36728 4072
rect 31536 4032 36728 4060
rect 31536 4020 31542 4032
rect 36722 4020 36728 4032
rect 36780 4020 36786 4072
rect 40954 4020 40960 4072
rect 41012 4060 41018 4072
rect 46842 4060 46848 4072
rect 41012 4032 46848 4060
rect 41012 4020 41018 4032
rect 46842 4020 46848 4032
rect 46900 4020 46906 4072
rect 50522 4020 50528 4072
rect 50580 4060 50586 4072
rect 56502 4060 56508 4072
rect 50580 4032 56508 4060
rect 50580 4020 50586 4032
rect 56502 4020 56508 4032
rect 56560 4020 56566 4072
rect 59998 4020 60004 4072
rect 60056 4060 60062 4072
rect 65794 4060 65800 4072
rect 60056 4032 65800 4060
rect 60056 4020 60062 4032
rect 65794 4020 65800 4032
rect 65852 4020 65858 4072
rect 69474 4020 69480 4072
rect 69532 4060 69538 4072
rect 74902 4060 74908 4072
rect 69532 4032 74908 4060
rect 69532 4020 69538 4032
rect 74902 4020 74908 4032
rect 74960 4020 74966 4072
rect 90726 4020 90732 4072
rect 90784 4060 90790 4072
rect 95602 4060 95608 4072
rect 90784 4032 95608 4060
rect 90784 4020 90790 4032
rect 95602 4020 95608 4032
rect 95660 4020 95666 4072
rect 99282 4020 99288 4072
rect 99340 4060 99346 4072
rect 103606 4060 103612 4072
rect 99340 4032 103612 4060
rect 99340 4020 99346 4032
rect 103606 4020 103612 4032
rect 103664 4020 103670 4072
rect 307938 4020 307944 4072
rect 307996 4060 308002 4072
rect 309778 4060 309784 4072
rect 307996 4032 309784 4060
rect 307996 4020 308002 4032
rect 309778 4020 309784 4032
rect 309836 4020 309842 4072
rect 324314 4020 324320 4072
rect 324372 4060 324378 4072
rect 326430 4060 326436 4072
rect 324372 4032 326436 4060
rect 324372 4020 324378 4032
rect 326430 4020 326436 4032
rect 326488 4020 326494 4072
rect 343634 4020 343640 4072
rect 343692 4060 343698 4072
rect 346670 4060 346676 4072
rect 343692 4032 346676 4060
rect 343692 4020 343698 4032
rect 346670 4020 346676 4032
rect 346728 4020 346734 4072
rect 352282 4020 352288 4072
rect 352340 4060 352346 4072
rect 354950 4060 354956 4072
rect 352340 4032 354956 4060
rect 352340 4020 352346 4032
rect 354950 4020 354956 4032
rect 355008 4020 355014 4072
rect 362954 4020 362960 4072
rect 363012 4060 363018 4072
rect 366910 4060 366916 4072
rect 363012 4032 366916 4060
rect 363012 4020 363018 4032
rect 366910 4020 366916 4032
rect 366968 4020 366974 4072
rect 371050 4020 371056 4072
rect 371108 4060 371114 4072
rect 373994 4060 374000 4072
rect 371108 4032 374000 4060
rect 371108 4020 371114 4032
rect 373994 4020 374000 4032
rect 374052 4020 374058 4072
rect 382366 4020 382372 4072
rect 382424 4060 382430 4072
rect 385862 4060 385868 4072
rect 382424 4032 385868 4060
rect 382424 4020 382430 4032
rect 385862 4020 385868 4032
rect 385920 4020 385926 4072
rect 393590 4020 393596 4072
rect 393648 4060 393654 4072
rect 397822 4060 397828 4072
rect 393648 4032 397828 4060
rect 393648 4020 393654 4032
rect 397822 4020 397828 4032
rect 397880 4020 397886 4072
rect 400490 4020 400496 4072
rect 400548 4060 400554 4072
rect 404906 4060 404912 4072
rect 400548 4032 404912 4060
rect 400548 4020 400554 4032
rect 404906 4020 404912 4032
rect 404964 4020 404970 4072
rect 409414 4020 409420 4072
rect 409472 4060 409478 4072
rect 413278 4060 413284 4072
rect 409472 4032 413284 4060
rect 409472 4020 409478 4032
rect 413278 4020 413284 4032
rect 413336 4020 413342 4072
rect 418154 4020 418160 4072
rect 418212 4060 418218 4072
rect 423950 4060 423956 4072
rect 418212 4032 423956 4060
rect 418212 4020 418218 4032
rect 423950 4020 423956 4032
rect 424008 4020 424014 4072
rect 429194 4020 429200 4072
rect 429252 4060 429258 4072
rect 434622 4060 434628 4072
rect 429252 4032 434628 4060
rect 429252 4020 429258 4032
rect 434622 4020 434628 4032
rect 434680 4020 434686 4072
rect 438578 4020 438584 4072
rect 438636 4060 438642 4072
rect 444190 4060 444196 4072
rect 438636 4032 444196 4060
rect 438636 4020 438642 4032
rect 444190 4020 444196 4032
rect 444248 4020 444254 4072
rect 457530 4020 457536 4072
rect 457588 4060 457594 4072
rect 463234 4060 463240 4072
rect 457588 4032 463240 4060
rect 457588 4020 457594 4032
rect 463234 4020 463240 4032
rect 463292 4020 463298 4072
rect 564434 4020 564440 4072
rect 564492 4060 564498 4072
rect 567838 4060 567844 4072
rect 564492 4032 567844 4060
rect 564492 4020 564498 4032
rect 567838 4020 567844 4032
rect 567896 4020 567902 4072
rect 570138 4020 570144 4072
rect 570196 4060 570202 4072
rect 573818 4060 573824 4072
rect 570196 4032 573824 4060
rect 570196 4020 570202 4032
rect 573818 4020 573824 4032
rect 573876 4020 573882 4072
rect 11238 3952 11244 4004
rect 11296 3992 11302 4004
rect 17586 3992 17592 4004
rect 11296 3964 17592 3992
rect 11296 3952 11302 3964
rect 17586 3952 17592 3964
rect 17644 3952 17650 4004
rect 55398 3952 55404 4004
rect 55456 3992 55462 4004
rect 61194 3992 61200 4004
rect 55456 3964 61200 3992
rect 55456 3952 55462 3964
rect 61194 3952 61200 3964
rect 61252 3952 61258 4004
rect 74258 3952 74264 4004
rect 74316 3992 74322 4004
rect 79502 3992 79508 4004
rect 74316 3964 79508 3992
rect 74316 3952 74322 3964
rect 79502 3952 79508 3964
rect 79560 3952 79566 4004
rect 314654 3952 314660 4004
rect 314712 3992 314718 4004
rect 316954 3992 316960 4004
rect 314712 3964 316960 3992
rect 314712 3952 314718 3964
rect 316954 3952 316960 3964
rect 317012 3952 317018 4004
rect 399846 3952 399852 4004
rect 399904 3992 399910 4004
rect 403710 3992 403716 4004
rect 399904 3964 403716 3992
rect 399904 3952 399910 3964
rect 403710 3952 403716 3964
rect 403768 3952 403774 4004
rect 571334 3952 571340 4004
rect 571392 3992 571398 4004
rect 575014 3992 575020 4004
rect 571392 3964 575020 3992
rect 571392 3952 571398 3964
rect 575014 3952 575020 3964
rect 575072 3952 575078 4004
rect 14826 3884 14832 3936
rect 14884 3924 14890 3936
rect 19426 3924 19432 3936
rect 14884 3896 19432 3924
rect 14884 3884 14890 3896
rect 19426 3884 19432 3896
rect 19484 3884 19490 3936
rect 25498 3884 25504 3936
rect 25556 3924 25562 3936
rect 30374 3924 30380 3936
rect 25556 3896 30380 3924
rect 25556 3884 25562 3896
rect 30374 3884 30380 3896
rect 30432 3884 30438 3936
rect 52822 3884 52828 3936
rect 52880 3924 52886 3936
rect 58894 3924 58900 3936
rect 52880 3896 58900 3924
rect 52880 3884 52886 3896
rect 58894 3884 58900 3896
rect 58952 3884 58958 3936
rect 63586 3884 63592 3936
rect 63644 3924 63650 3936
rect 69198 3924 69204 3936
rect 63644 3896 69204 3924
rect 63644 3884 63650 3896
rect 69198 3884 69204 3896
rect 69256 3884 69262 3936
rect 316494 3884 316500 3936
rect 316552 3924 316558 3936
rect 318058 3924 318064 3936
rect 316552 3896 318064 3924
rect 316552 3884 316558 3896
rect 318058 3884 318064 3896
rect 318116 3884 318122 3936
rect 335814 3884 335820 3936
rect 335872 3924 335878 3936
rect 337102 3924 337108 3936
rect 335872 3896 337108 3924
rect 335872 3884 335878 3896
rect 337102 3884 337108 3896
rect 337160 3884 337166 3936
rect 361574 3884 361580 3936
rect 361632 3924 361638 3936
rect 364518 3924 364524 3936
rect 361632 3896 364524 3924
rect 361632 3884 361638 3896
rect 364518 3884 364524 3896
rect 364576 3884 364582 3936
rect 442074 3884 442080 3936
rect 442132 3924 442138 3936
rect 447778 3924 447784 3936
rect 442132 3896 447784 3924
rect 442132 3884 442138 3896
rect 447778 3884 447784 3896
rect 447836 3884 447842 3936
rect 448606 3884 448612 3936
rect 448664 3924 448670 3936
rect 454862 3924 454868 3936
rect 448664 3896 454868 3924
rect 448664 3884 448670 3896
rect 454862 3884 454868 3896
rect 454920 3884 454926 3936
rect 490374 3884 490380 3936
rect 490432 3924 490438 3936
rect 498930 3924 498936 3936
rect 490432 3896 498936 3924
rect 490432 3884 490438 3896
rect 498930 3884 498936 3896
rect 498988 3884 498994 3936
rect 1104 3834 582820 3856
rect 1104 3782 18822 3834
rect 18874 3782 18886 3834
rect 18938 3782 18950 3834
rect 19002 3782 19014 3834
rect 19066 3782 19078 3834
rect 19130 3782 19142 3834
rect 19194 3782 19206 3834
rect 19258 3782 19270 3834
rect 19322 3782 19334 3834
rect 19386 3782 54822 3834
rect 54874 3782 54886 3834
rect 54938 3782 54950 3834
rect 55002 3782 55014 3834
rect 55066 3782 55078 3834
rect 55130 3782 55142 3834
rect 55194 3782 55206 3834
rect 55258 3782 55270 3834
rect 55322 3782 55334 3834
rect 55386 3782 90822 3834
rect 90874 3782 90886 3834
rect 90938 3782 90950 3834
rect 91002 3782 91014 3834
rect 91066 3782 91078 3834
rect 91130 3782 91142 3834
rect 91194 3782 91206 3834
rect 91258 3782 91270 3834
rect 91322 3782 91334 3834
rect 91386 3782 126822 3834
rect 126874 3782 126886 3834
rect 126938 3782 126950 3834
rect 127002 3782 127014 3834
rect 127066 3782 127078 3834
rect 127130 3782 127142 3834
rect 127194 3782 127206 3834
rect 127258 3782 127270 3834
rect 127322 3782 127334 3834
rect 127386 3782 162822 3834
rect 162874 3782 162886 3834
rect 162938 3782 162950 3834
rect 163002 3782 163014 3834
rect 163066 3782 163078 3834
rect 163130 3782 163142 3834
rect 163194 3782 163206 3834
rect 163258 3782 163270 3834
rect 163322 3782 163334 3834
rect 163386 3782 198822 3834
rect 198874 3782 198886 3834
rect 198938 3782 198950 3834
rect 199002 3782 199014 3834
rect 199066 3782 199078 3834
rect 199130 3782 199142 3834
rect 199194 3782 199206 3834
rect 199258 3782 199270 3834
rect 199322 3782 199334 3834
rect 199386 3782 234822 3834
rect 234874 3782 234886 3834
rect 234938 3782 234950 3834
rect 235002 3782 235014 3834
rect 235066 3782 235078 3834
rect 235130 3782 235142 3834
rect 235194 3782 235206 3834
rect 235258 3782 235270 3834
rect 235322 3782 235334 3834
rect 235386 3782 270822 3834
rect 270874 3782 270886 3834
rect 270938 3782 270950 3834
rect 271002 3782 271014 3834
rect 271066 3782 271078 3834
rect 271130 3782 271142 3834
rect 271194 3782 271206 3834
rect 271258 3782 271270 3834
rect 271322 3782 271334 3834
rect 271386 3782 306822 3834
rect 306874 3782 306886 3834
rect 306938 3782 306950 3834
rect 307002 3782 307014 3834
rect 307066 3782 307078 3834
rect 307130 3782 307142 3834
rect 307194 3782 307206 3834
rect 307258 3782 307270 3834
rect 307322 3782 307334 3834
rect 307386 3782 342822 3834
rect 342874 3782 342886 3834
rect 342938 3782 342950 3834
rect 343002 3782 343014 3834
rect 343066 3782 343078 3834
rect 343130 3782 343142 3834
rect 343194 3782 343206 3834
rect 343258 3782 343270 3834
rect 343322 3782 343334 3834
rect 343386 3782 378822 3834
rect 378874 3782 378886 3834
rect 378938 3782 378950 3834
rect 379002 3782 379014 3834
rect 379066 3782 379078 3834
rect 379130 3782 379142 3834
rect 379194 3782 379206 3834
rect 379258 3782 379270 3834
rect 379322 3782 379334 3834
rect 379386 3782 414822 3834
rect 414874 3782 414886 3834
rect 414938 3782 414950 3834
rect 415002 3782 415014 3834
rect 415066 3782 415078 3834
rect 415130 3782 415142 3834
rect 415194 3782 415206 3834
rect 415258 3782 415270 3834
rect 415322 3782 415334 3834
rect 415386 3782 450822 3834
rect 450874 3782 450886 3834
rect 450938 3782 450950 3834
rect 451002 3782 451014 3834
rect 451066 3782 451078 3834
rect 451130 3782 451142 3834
rect 451194 3782 451206 3834
rect 451258 3782 451270 3834
rect 451322 3782 451334 3834
rect 451386 3782 486822 3834
rect 486874 3782 486886 3834
rect 486938 3782 486950 3834
rect 487002 3782 487014 3834
rect 487066 3782 487078 3834
rect 487130 3782 487142 3834
rect 487194 3782 487206 3834
rect 487258 3782 487270 3834
rect 487322 3782 487334 3834
rect 487386 3782 522822 3834
rect 522874 3782 522886 3834
rect 522938 3782 522950 3834
rect 523002 3782 523014 3834
rect 523066 3782 523078 3834
rect 523130 3782 523142 3834
rect 523194 3782 523206 3834
rect 523258 3782 523270 3834
rect 523322 3782 523334 3834
rect 523386 3782 558822 3834
rect 558874 3782 558886 3834
rect 558938 3782 558950 3834
rect 559002 3782 559014 3834
rect 559066 3782 559078 3834
rect 559130 3782 559142 3834
rect 559194 3782 559206 3834
rect 559258 3782 559270 3834
rect 559322 3782 559334 3834
rect 559386 3782 582820 3834
rect 1104 3760 582820 3782
rect 5258 3680 5264 3732
rect 5316 3720 5322 3732
rect 12342 3720 12348 3732
rect 5316 3692 12348 3720
rect 5316 3680 5322 3692
rect 12342 3680 12348 3692
rect 12400 3680 12406 3732
rect 44542 3680 44548 3732
rect 44600 3720 44606 3732
rect 50890 3720 50896 3732
rect 44600 3692 50896 3720
rect 44600 3680 44606 3692
rect 50890 3680 50896 3692
rect 50948 3680 50954 3732
rect 61194 3680 61200 3732
rect 61252 3720 61258 3732
rect 66898 3720 66904 3732
rect 61252 3692 66904 3720
rect 61252 3680 61258 3692
rect 66898 3680 66904 3692
rect 66956 3680 66962 3732
rect 353294 3680 353300 3732
rect 353352 3720 353358 3732
rect 356146 3720 356152 3732
rect 353352 3692 356152 3720
rect 353352 3680 353358 3692
rect 356146 3680 356152 3692
rect 356204 3680 356210 3732
rect 374730 3680 374736 3732
rect 374788 3720 374794 3732
rect 377582 3720 377588 3732
rect 374788 3692 377588 3720
rect 374788 3680 374794 3692
rect 377582 3680 377588 3692
rect 377640 3680 377646 3732
rect 384942 3680 384948 3732
rect 385000 3720 385006 3732
rect 388254 3720 388260 3732
rect 385000 3692 388260 3720
rect 385000 3680 385006 3692
rect 388254 3680 388260 3692
rect 388312 3680 388318 3732
rect 403894 3680 403900 3732
rect 403952 3720 403958 3732
rect 408494 3720 408500 3732
rect 403952 3692 408500 3720
rect 403952 3680 403958 3692
rect 408494 3680 408500 3692
rect 408552 3680 408558 3732
rect 420914 3680 420920 3732
rect 420972 3720 420978 3732
rect 426342 3720 426348 3732
rect 420972 3692 426348 3720
rect 420972 3680 420978 3692
rect 426342 3680 426348 3692
rect 426400 3680 426406 3732
rect 449894 3680 449900 3732
rect 449952 3720 449958 3732
rect 456058 3720 456064 3732
rect 449952 3692 456064 3720
rect 449952 3680 449958 3692
rect 456058 3680 456064 3692
rect 456116 3680 456122 3732
rect 553394 3680 553400 3732
rect 553452 3720 553458 3732
rect 555970 3720 555976 3732
rect 553452 3692 555976 3720
rect 553452 3680 553458 3692
rect 555970 3680 555976 3692
rect 556028 3680 556034 3732
rect 6454 3612 6460 3664
rect 6512 3652 6518 3664
rect 12526 3652 12532 3664
rect 6512 3624 12532 3652
rect 6512 3612 6518 3624
rect 12526 3612 12532 3624
rect 12584 3612 12590 3664
rect 16022 3612 16028 3664
rect 16080 3652 16086 3664
rect 20806 3652 20812 3664
rect 16080 3624 20812 3652
rect 16080 3612 16086 3624
rect 20806 3612 20812 3624
rect 20864 3612 20870 3664
rect 36170 3612 36176 3664
rect 36228 3652 36234 3664
rect 42610 3652 42616 3664
rect 36228 3624 42616 3652
rect 36228 3612 36234 3624
rect 42610 3612 42616 3624
rect 42668 3612 42674 3664
rect 43346 3612 43352 3664
rect 43404 3652 43410 3664
rect 49602 3652 49608 3664
rect 43404 3624 49608 3652
rect 43404 3612 43410 3624
rect 49602 3612 49608 3624
rect 49660 3612 49666 3664
rect 54018 3612 54024 3664
rect 54076 3652 54082 3664
rect 60090 3652 60096 3664
rect 54076 3624 60096 3652
rect 54076 3612 54082 3624
rect 60090 3612 60096 3624
rect 60148 3612 60154 3664
rect 401594 3612 401600 3664
rect 401652 3652 401658 3664
rect 406102 3652 406108 3664
rect 401652 3624 406108 3652
rect 401652 3612 401658 3624
rect 406102 3612 406108 3624
rect 406160 3612 406166 3664
rect 429838 3612 429844 3664
rect 429896 3652 429902 3664
rect 435818 3652 435824 3664
rect 429896 3624 435824 3652
rect 429896 3612 429902 3624
rect 435818 3612 435824 3624
rect 435876 3612 435882 3664
rect 440326 3612 440332 3664
rect 440384 3652 440390 3664
rect 446582 3652 446588 3664
rect 440384 3624 446588 3652
rect 440384 3612 440390 3624
rect 446582 3612 446588 3624
rect 446640 3612 446646 3664
rect 27890 3544 27896 3596
rect 27948 3584 27954 3596
rect 34330 3584 34336 3596
rect 27948 3556 34336 3584
rect 27948 3544 27954 3556
rect 34330 3544 34336 3556
rect 34388 3544 34394 3596
rect 34974 3544 34980 3596
rect 35032 3584 35038 3596
rect 40034 3584 40040 3596
rect 35032 3556 40040 3584
rect 35032 3544 35038 3556
rect 40034 3544 40040 3556
rect 40092 3544 40098 3596
rect 57606 3544 57612 3596
rect 57664 3584 57670 3596
rect 62114 3584 62120 3596
rect 57664 3556 62120 3584
rect 57664 3544 57670 3556
rect 62114 3544 62120 3556
rect 62172 3544 62178 3596
rect 67174 3544 67180 3596
rect 67232 3584 67238 3596
rect 72326 3584 72332 3596
rect 67232 3556 72332 3584
rect 67232 3544 67238 3556
rect 72326 3544 72332 3556
rect 72384 3544 72390 3596
rect 72694 3544 72700 3596
rect 72752 3584 72758 3596
rect 78398 3584 78404 3596
rect 72752 3556 78404 3584
rect 72752 3544 72758 3556
rect 78398 3544 78404 3556
rect 78456 3544 78462 3596
rect 82630 3544 82636 3596
rect 82688 3584 82694 3596
rect 87506 3584 87512 3596
rect 82688 3556 87512 3584
rect 82688 3544 82694 3556
rect 87506 3544 87512 3556
rect 87564 3544 87570 3596
rect 342714 3544 342720 3596
rect 342772 3584 342778 3596
rect 345474 3584 345480 3596
rect 342772 3556 345480 3584
rect 342772 3544 342778 3556
rect 345474 3544 345480 3556
rect 345532 3544 345538 3596
rect 347774 3544 347780 3596
rect 347832 3584 347838 3596
rect 350258 3584 350264 3596
rect 347832 3556 350264 3584
rect 347832 3544 347838 3556
rect 350258 3544 350264 3556
rect 350316 3544 350322 3596
rect 358170 3544 358176 3596
rect 358228 3584 358234 3596
rect 360746 3584 360752 3596
rect 358228 3556 360752 3584
rect 358228 3544 358234 3556
rect 360746 3544 360752 3556
rect 360804 3544 360810 3596
rect 362218 3544 362224 3596
rect 362276 3584 362282 3596
rect 365714 3584 365720 3596
rect 362276 3556 365720 3584
rect 362276 3544 362282 3556
rect 365714 3544 365720 3556
rect 365772 3544 365778 3596
rect 369762 3544 369768 3596
rect 369820 3584 369826 3596
rect 372798 3584 372804 3596
rect 369820 3556 372804 3584
rect 369820 3544 369826 3556
rect 372798 3544 372804 3556
rect 372856 3544 372862 3596
rect 379422 3544 379428 3596
rect 379480 3584 379486 3596
rect 382366 3584 382372 3596
rect 379480 3556 382372 3584
rect 379480 3544 379486 3556
rect 382366 3544 382372 3556
rect 382424 3544 382430 3596
rect 389174 3544 389180 3596
rect 389232 3584 389238 3596
rect 394234 3584 394240 3596
rect 389232 3556 394240 3584
rect 389232 3544 389238 3556
rect 394234 3544 394240 3556
rect 394292 3544 394298 3596
rect 396534 3544 396540 3596
rect 396592 3584 396598 3596
rect 400214 3584 400220 3596
rect 396592 3556 400220 3584
rect 396592 3544 396598 3556
rect 400214 3544 400220 3556
rect 400272 3544 400278 3596
rect 408402 3544 408408 3596
rect 408460 3584 408466 3596
rect 412082 3584 412088 3596
rect 408460 3556 412088 3584
rect 408460 3544 408466 3556
rect 412082 3544 412088 3556
rect 412140 3544 412146 3596
rect 416498 3544 416504 3596
rect 416556 3584 416562 3596
rect 420362 3584 420368 3596
rect 416556 3556 420368 3584
rect 416556 3544 416562 3556
rect 420362 3544 420368 3556
rect 420420 3544 420426 3596
rect 430574 3544 430580 3596
rect 430632 3584 430638 3596
rect 437014 3584 437020 3596
rect 430632 3556 437020 3584
rect 430632 3544 430638 3556
rect 437014 3544 437020 3556
rect 437072 3544 437078 3596
rect 516134 3544 516140 3596
rect 516192 3584 516198 3596
rect 517882 3584 517888 3596
rect 516192 3556 517888 3584
rect 516192 3544 516198 3556
rect 517882 3544 517888 3556
rect 517940 3544 517946 3596
rect 531314 3544 531320 3596
rect 531372 3584 531378 3596
rect 533430 3584 533436 3596
rect 531372 3556 533436 3584
rect 531372 3544 531378 3556
rect 533430 3544 533436 3556
rect 533488 3544 533494 3596
rect 545114 3544 545120 3596
rect 545172 3584 545178 3596
rect 547690 3584 547696 3596
rect 545172 3556 547696 3584
rect 545172 3544 545178 3556
rect 547690 3544 547696 3556
rect 547748 3544 547754 3596
rect 556154 3544 556160 3596
rect 556212 3584 556218 3596
rect 559558 3584 559564 3596
rect 556212 3556 559564 3584
rect 556212 3544 556218 3556
rect 559558 3544 559564 3556
rect 559616 3544 559622 3596
rect 4062 3476 4068 3528
rect 4120 3516 4126 3528
rect 11974 3516 11980 3528
rect 4120 3488 11980 3516
rect 4120 3476 4126 3488
rect 11974 3476 11980 3488
rect 12032 3476 12038 3528
rect 17218 3476 17224 3528
rect 17276 3516 17282 3528
rect 22094 3516 22100 3528
rect 17276 3488 22100 3516
rect 17276 3476 17282 3488
rect 22094 3476 22100 3488
rect 22152 3476 22158 3528
rect 24302 3476 24308 3528
rect 24360 3516 24366 3528
rect 28994 3516 29000 3528
rect 24360 3488 29000 3516
rect 24360 3476 24366 3488
rect 28994 3476 29000 3488
rect 29052 3476 29058 3528
rect 37458 3476 37464 3528
rect 37516 3516 37522 3528
rect 43990 3516 43996 3528
rect 37516 3488 43996 3516
rect 37516 3476 37522 3488
rect 43990 3476 43996 3488
rect 44048 3476 44054 3528
rect 46934 3476 46940 3528
rect 46992 3516 46998 3528
rect 53190 3516 53196 3528
rect 46992 3488 53196 3516
rect 46992 3476 46998 3488
rect 53190 3476 53196 3488
rect 53248 3476 53254 3528
rect 56410 3476 56416 3528
rect 56468 3516 56474 3528
rect 61930 3516 61936 3528
rect 56468 3488 61936 3516
rect 56468 3476 56474 3488
rect 61930 3476 61936 3488
rect 61988 3476 61994 3528
rect 62390 3476 62396 3528
rect 62448 3516 62454 3528
rect 68094 3516 68100 3528
rect 62448 3488 68100 3516
rect 62448 3476 62454 3488
rect 68094 3476 68100 3488
rect 68152 3476 68158 3528
rect 68278 3476 68284 3528
rect 68336 3516 68342 3528
rect 73798 3516 73804 3528
rect 68336 3488 73804 3516
rect 68336 3476 68342 3488
rect 73798 3476 73804 3488
rect 73856 3476 73862 3528
rect 76650 3476 76656 3528
rect 76708 3516 76714 3528
rect 81802 3516 81808 3528
rect 76708 3488 81808 3516
rect 76708 3476 76714 3488
rect 81802 3476 81808 3488
rect 81860 3476 81866 3528
rect 83826 3476 83832 3528
rect 83884 3516 83890 3528
rect 88702 3516 88708 3528
rect 83884 3488 88708 3516
rect 83884 3476 83890 3488
rect 88702 3476 88708 3488
rect 88760 3476 88766 3528
rect 92106 3476 92112 3528
rect 92164 3516 92170 3528
rect 96706 3516 96712 3528
rect 92164 3488 96712 3516
rect 92164 3476 92170 3488
rect 96706 3476 96712 3488
rect 96764 3476 96770 3528
rect 183738 3476 183744 3528
rect 183796 3516 183802 3528
rect 184842 3516 184848 3528
rect 183796 3488 184848 3516
rect 183796 3476 183802 3488
rect 184842 3476 184848 3488
rect 184900 3476 184906 3528
rect 190822 3476 190828 3528
rect 190880 3516 190886 3528
rect 191742 3516 191748 3528
rect 190880 3488 191748 3516
rect 190880 3476 190886 3488
rect 191742 3476 191748 3488
rect 191800 3476 191806 3528
rect 192018 3476 192024 3528
rect 192076 3516 192082 3528
rect 192938 3516 192944 3528
rect 192076 3488 192944 3516
rect 192076 3476 192082 3488
rect 192938 3476 192944 3488
rect 192996 3476 193002 3528
rect 193214 3476 193220 3528
rect 193272 3516 193278 3528
rect 194042 3516 194048 3528
rect 193272 3488 194048 3516
rect 193272 3476 193278 3488
rect 194042 3476 194048 3488
rect 194100 3476 194106 3528
rect 236454 3476 236460 3528
rect 236512 3516 236518 3528
rect 237190 3516 237196 3528
rect 236512 3488 237196 3516
rect 236512 3476 236518 3488
rect 237190 3476 237196 3488
rect 237248 3476 237254 3528
rect 237558 3476 237564 3528
rect 237616 3516 237622 3528
rect 238386 3516 238392 3528
rect 237616 3488 238392 3516
rect 237616 3476 237622 3488
rect 238386 3476 238392 3488
rect 238444 3476 238450 3528
rect 244458 3476 244464 3528
rect 244516 3516 244522 3528
rect 245562 3516 245568 3528
rect 244516 3488 245568 3516
rect 244516 3476 244522 3488
rect 245562 3476 245568 3488
rect 245620 3476 245626 3528
rect 301038 3476 301044 3528
rect 301096 3516 301102 3528
rect 302602 3516 302608 3528
rect 301096 3488 302608 3516
rect 301096 3476 301102 3488
rect 302602 3476 302608 3488
rect 302660 3476 302666 3528
rect 322014 3476 322020 3528
rect 322072 3516 322078 3528
rect 324038 3516 324044 3528
rect 322072 3488 324044 3516
rect 322072 3476 322078 3488
rect 324038 3476 324044 3488
rect 324096 3476 324102 3528
rect 324130 3476 324136 3528
rect 324188 3516 324194 3528
rect 325418 3516 325424 3528
rect 324188 3488 325424 3516
rect 324188 3476 324194 3488
rect 325418 3476 325424 3488
rect 325476 3476 325482 3528
rect 331306 3476 331312 3528
rect 331364 3516 331370 3528
rect 333606 3516 333612 3528
rect 331364 3488 333612 3516
rect 331364 3476 331370 3488
rect 333606 3476 333612 3488
rect 333664 3476 333670 3528
rect 338298 3476 338304 3528
rect 338356 3516 338362 3528
rect 340690 3516 340696 3528
rect 338356 3488 340696 3516
rect 338356 3476 338362 3488
rect 340690 3476 340696 3488
rect 340748 3476 340754 3528
rect 342254 3476 342260 3528
rect 342312 3516 342318 3528
rect 344278 3516 344284 3528
rect 342312 3488 344284 3516
rect 342312 3476 342318 3488
rect 344278 3476 344284 3488
rect 344336 3476 344342 3528
rect 349154 3476 349160 3528
rect 349212 3516 349218 3528
rect 351362 3516 351368 3528
rect 349212 3488 351368 3516
rect 349212 3476 349218 3488
rect 351362 3476 351368 3488
rect 351420 3476 351426 3528
rect 359366 3476 359372 3528
rect 359424 3516 359430 3528
rect 362126 3516 362132 3528
rect 359424 3488 362132 3516
rect 359424 3476 359430 3488
rect 362126 3476 362132 3488
rect 362184 3476 362190 3528
rect 367462 3476 367468 3528
rect 367520 3516 367526 3528
rect 370406 3516 370412 3528
rect 367520 3488 370412 3516
rect 367520 3476 367526 3488
rect 370406 3476 370412 3488
rect 370464 3476 370470 3528
rect 378042 3476 378048 3528
rect 378100 3516 378106 3528
rect 381170 3516 381176 3528
rect 378100 3488 381176 3516
rect 378100 3476 378106 3488
rect 381170 3476 381176 3488
rect 381228 3476 381234 3528
rect 382274 3476 382280 3528
rect 382332 3516 382338 3528
rect 387058 3516 387064 3528
rect 382332 3488 387064 3516
rect 382332 3476 382338 3488
rect 387058 3476 387064 3488
rect 387116 3476 387122 3528
rect 387334 3476 387340 3528
rect 387392 3516 387398 3528
rect 390646 3516 390652 3528
rect 387392 3488 390652 3516
rect 387392 3476 387398 3488
rect 390646 3476 390652 3488
rect 390704 3476 390710 3528
rect 391934 3476 391940 3528
rect 391992 3516 391998 3528
rect 396626 3516 396632 3528
rect 391992 3488 396632 3516
rect 391992 3476 391998 3488
rect 396626 3476 396632 3488
rect 396684 3476 396690 3528
rect 398742 3476 398748 3528
rect 398800 3516 398806 3528
rect 402514 3516 402520 3528
rect 398800 3488 402520 3516
rect 398800 3476 398806 3488
rect 402514 3476 402520 3488
rect 402572 3476 402578 3528
rect 410426 3476 410432 3528
rect 410484 3516 410490 3528
rect 415670 3516 415676 3528
rect 410484 3488 415676 3516
rect 410484 3476 410490 3488
rect 415670 3476 415676 3488
rect 415728 3476 415734 3528
rect 419810 3476 419816 3528
rect 419868 3516 419874 3528
rect 425146 3516 425152 3528
rect 419868 3488 425152 3516
rect 419868 3476 419874 3488
rect 425146 3476 425152 3488
rect 425204 3476 425210 3528
rect 426250 3476 426256 3528
rect 426308 3516 426314 3528
rect 431126 3516 431132 3528
rect 426308 3488 431132 3516
rect 426308 3476 426314 3488
rect 431126 3476 431132 3488
rect 431184 3476 431190 3528
rect 436002 3476 436008 3528
rect 436060 3516 436066 3528
rect 440602 3516 440608 3528
rect 436060 3488 440608 3516
rect 436060 3476 436066 3488
rect 440602 3476 440608 3488
rect 440660 3476 440666 3528
rect 459554 3476 459560 3528
rect 459612 3516 459618 3528
rect 466822 3516 466828 3528
rect 459612 3488 466828 3516
rect 459612 3476 459618 3488
rect 466822 3476 466828 3488
rect 466880 3476 466886 3528
rect 551922 3476 551928 3528
rect 551980 3516 551986 3528
rect 560754 3516 560760 3528
rect 551980 3488 560760 3516
rect 551980 3476 551986 3488
rect 560754 3476 560760 3488
rect 560812 3476 560818 3528
rect 7650 3408 7656 3460
rect 7708 3448 7714 3460
rect 12434 3448 12440 3460
rect 7708 3420 12440 3448
rect 7708 3408 7714 3420
rect 12434 3408 12440 3420
rect 12492 3408 12498 3460
rect 26694 3408 26700 3460
rect 26752 3448 26758 3460
rect 31754 3448 31760 3460
rect 26752 3420 31760 3448
rect 26752 3408 26758 3420
rect 31754 3408 31760 3420
rect 31812 3408 31818 3460
rect 33870 3408 33876 3460
rect 33928 3448 33934 3460
rect 39850 3448 39856 3460
rect 33928 3420 39856 3448
rect 33928 3408 33934 3420
rect 39850 3408 39856 3420
rect 39908 3408 39914 3460
rect 48130 3408 48136 3460
rect 48188 3448 48194 3460
rect 53742 3448 53748 3460
rect 48188 3420 53748 3448
rect 48188 3408 48194 3420
rect 53742 3408 53748 3420
rect 53800 3408 53806 3460
rect 58802 3408 58808 3460
rect 58860 3448 58866 3460
rect 64598 3448 64604 3460
rect 58860 3420 64604 3448
rect 58860 3408 58866 3420
rect 64598 3408 64604 3420
rect 64656 3408 64662 3460
rect 64782 3408 64788 3460
rect 64840 3448 64846 3460
rect 70210 3448 70216 3460
rect 64840 3420 70216 3448
rect 64840 3408 64846 3420
rect 70210 3408 70216 3420
rect 70268 3408 70274 3460
rect 77846 3408 77852 3460
rect 77904 3448 77910 3460
rect 82998 3448 83004 3460
rect 77904 3420 83004 3448
rect 77904 3408 77910 3420
rect 82998 3408 83004 3420
rect 83056 3408 83062 3460
rect 329006 3408 329012 3460
rect 329064 3448 329070 3460
rect 331214 3448 331220 3460
rect 329064 3420 331220 3448
rect 329064 3408 329070 3420
rect 331214 3408 331220 3420
rect 331272 3408 331278 3460
rect 333974 3408 333980 3460
rect 334032 3448 334038 3460
rect 335906 3448 335912 3460
rect 334032 3420 335912 3448
rect 334032 3408 334038 3420
rect 335906 3408 335912 3420
rect 335964 3408 335970 3460
rect 340874 3408 340880 3460
rect 340932 3448 340938 3460
rect 342714 3448 342720 3460
rect 340932 3420 342720 3448
rect 340932 3408 340938 3420
rect 342714 3408 342720 3420
rect 342772 3408 342778 3460
rect 360562 3408 360568 3460
rect 360620 3448 360626 3460
rect 363322 3448 363328 3460
rect 360620 3420 363328 3448
rect 360620 3408 360626 3420
rect 363322 3408 363328 3420
rect 363380 3408 363386 3460
rect 372614 3408 372620 3460
rect 372672 3448 372678 3460
rect 376386 3448 376392 3460
rect 372672 3420 376392 3448
rect 372672 3408 372678 3420
rect 376386 3408 376392 3420
rect 376444 3408 376450 3460
rect 380434 3408 380440 3460
rect 380492 3448 380498 3460
rect 383562 3448 383568 3460
rect 380492 3420 383568 3448
rect 380492 3408 380498 3420
rect 383562 3408 383568 3420
rect 383620 3408 383626 3460
rect 388530 3408 388536 3460
rect 388588 3448 388594 3460
rect 391842 3448 391848 3460
rect 388588 3420 391848 3448
rect 388588 3408 388594 3420
rect 391842 3408 391848 3420
rect 391900 3408 391906 3460
rect 396718 3408 396724 3460
rect 396776 3448 396782 3460
rect 401318 3448 401324 3460
rect 396776 3420 401324 3448
rect 396776 3408 396782 3420
rect 401318 3408 401324 3420
rect 401376 3408 401382 3460
rect 407022 3408 407028 3460
rect 407080 3448 407086 3460
rect 410886 3448 410892 3460
rect 407080 3420 410892 3448
rect 407080 3408 407086 3420
rect 410886 3408 410892 3420
rect 410944 3408 410950 3460
rect 411254 3408 411260 3460
rect 411312 3448 411318 3460
rect 416866 3448 416872 3460
rect 411312 3420 416872 3448
rect 411312 3408 411318 3420
rect 416866 3408 416872 3420
rect 416924 3408 416930 3460
rect 416958 3408 416964 3460
rect 417016 3448 417022 3460
rect 422754 3448 422760 3460
rect 417016 3420 422760 3448
rect 417016 3408 417022 3420
rect 422754 3408 422760 3420
rect 422812 3408 422818 3460
rect 427814 3408 427820 3460
rect 427872 3448 427878 3460
rect 433518 3448 433524 3460
rect 427872 3420 433524 3448
rect 427872 3408 427878 3420
rect 433518 3408 433524 3420
rect 433576 3408 433582 3460
rect 439222 3408 439228 3460
rect 439280 3448 439286 3460
rect 445386 3448 445392 3460
rect 439280 3420 445392 3448
rect 439280 3408 439286 3420
rect 445386 3408 445392 3420
rect 445444 3408 445450 3460
rect 445478 3408 445484 3460
rect 445536 3448 445542 3460
rect 451458 3448 451464 3460
rect 445536 3420 451464 3448
rect 445536 3408 445542 3420
rect 451458 3408 451464 3420
rect 451516 3408 451522 3460
rect 458634 3408 458640 3460
rect 458692 3448 458698 3460
rect 465626 3448 465632 3460
rect 458692 3420 465632 3448
rect 458692 3408 458698 3420
rect 465626 3408 465632 3420
rect 465684 3408 465690 3460
rect 473354 3408 473360 3460
rect 473412 3448 473418 3460
rect 481082 3448 481088 3460
rect 473412 3420 481088 3448
rect 473412 3408 473418 3420
rect 481082 3408 481088 3420
rect 481140 3408 481146 3460
rect 506290 3408 506296 3460
rect 506348 3448 506354 3460
rect 514386 3448 514392 3460
rect 506348 3420 514392 3448
rect 506348 3408 506354 3420
rect 514386 3408 514392 3420
rect 514444 3408 514450 3460
rect 521562 3408 521568 3460
rect 521620 3448 521626 3460
rect 529842 3448 529848 3460
rect 521620 3420 529848 3448
rect 521620 3408 521626 3420
rect 529842 3408 529848 3420
rect 529900 3408 529906 3460
rect 535454 3408 535460 3460
rect 535512 3448 535518 3460
rect 545298 3448 545304 3460
rect 535512 3420 545304 3448
rect 535512 3408 535518 3420
rect 545298 3408 545304 3420
rect 545356 3408 545362 3460
rect 546586 3408 546592 3460
rect 546644 3448 546650 3460
rect 550082 3448 550088 3460
rect 546644 3420 550088 3448
rect 546644 3408 546650 3420
rect 550082 3408 550088 3420
rect 550140 3408 550146 3460
rect 550726 3408 550732 3460
rect 550784 3448 550790 3460
rect 561950 3448 561956 3460
rect 550784 3420 561956 3448
rect 550784 3408 550790 3420
rect 561950 3408 561956 3420
rect 562008 3408 562014 3460
rect 568390 3408 568396 3460
rect 568448 3448 568454 3460
rect 570230 3448 570236 3460
rect 568448 3420 570236 3448
rect 568448 3408 568454 3420
rect 570230 3408 570236 3420
rect 570288 3408 570294 3460
rect 38562 3340 38568 3392
rect 38620 3380 38626 3392
rect 42794 3380 42800 3392
rect 38620 3352 42800 3380
rect 38620 3340 38626 3352
rect 42794 3340 42800 3352
rect 42852 3340 42858 3392
rect 332594 3340 332600 3392
rect 332652 3380 332658 3392
rect 334710 3380 334716 3392
rect 332652 3352 334716 3380
rect 332652 3340 332658 3352
rect 334710 3340 334716 3352
rect 334768 3340 334774 3392
rect 339494 3340 339500 3392
rect 339552 3380 339558 3392
rect 341886 3380 341892 3392
rect 339552 3352 341892 3380
rect 339552 3340 339558 3352
rect 341886 3340 341892 3352
rect 341944 3340 341950 3392
rect 389634 3340 389640 3392
rect 389692 3380 389698 3392
rect 393038 3380 393044 3392
rect 389692 3352 393044 3380
rect 389692 3340 389698 3352
rect 393038 3340 393044 3352
rect 393096 3340 393102 3392
rect 416682 3340 416688 3392
rect 416740 3380 416746 3392
rect 421558 3380 421564 3392
rect 416740 3352 421564 3380
rect 416740 3340 416746 3352
rect 421558 3340 421564 3352
rect 421616 3340 421622 3392
rect 436094 3340 436100 3392
rect 436152 3380 436158 3392
rect 441798 3380 441804 3392
rect 436152 3352 441804 3380
rect 436152 3340 436158 3352
rect 441798 3340 441804 3352
rect 441856 3340 441862 3392
rect 474734 3340 474740 3392
rect 474792 3380 474798 3392
rect 482278 3380 482284 3392
rect 474792 3352 482284 3380
rect 474792 3340 474798 3352
rect 482278 3340 482284 3352
rect 482336 3340 482342 3392
rect 541526 3340 541532 3392
rect 541584 3380 541590 3392
rect 542906 3380 542912 3392
rect 541584 3352 542912 3380
rect 541584 3340 541590 3352
rect 542906 3340 542912 3352
rect 542964 3340 542970 3392
rect 549530 3340 549536 3392
rect 549588 3380 549594 3392
rect 551186 3380 551192 3392
rect 549588 3352 551192 3380
rect 549588 3340 549594 3352
rect 551186 3340 551192 3352
rect 551244 3340 551250 3392
rect 556246 3340 556252 3392
rect 556304 3380 556310 3392
rect 558362 3380 558368 3392
rect 556304 3352 558368 3380
rect 556304 3340 556310 3352
rect 558362 3340 558368 3352
rect 558420 3340 558426 3392
rect 560386 3340 560392 3392
rect 560444 3380 560450 3392
rect 563146 3380 563152 3392
rect 560444 3352 563152 3380
rect 560444 3340 560450 3352
rect 563146 3340 563152 3352
rect 563204 3340 563210 3392
rect 1104 3290 582820 3312
rect 1104 3238 36822 3290
rect 36874 3238 36886 3290
rect 36938 3238 36950 3290
rect 37002 3238 37014 3290
rect 37066 3238 37078 3290
rect 37130 3238 37142 3290
rect 37194 3238 37206 3290
rect 37258 3238 37270 3290
rect 37322 3238 37334 3290
rect 37386 3238 72822 3290
rect 72874 3238 72886 3290
rect 72938 3238 72950 3290
rect 73002 3238 73014 3290
rect 73066 3238 73078 3290
rect 73130 3238 73142 3290
rect 73194 3238 73206 3290
rect 73258 3238 73270 3290
rect 73322 3238 73334 3290
rect 73386 3238 108822 3290
rect 108874 3238 108886 3290
rect 108938 3238 108950 3290
rect 109002 3238 109014 3290
rect 109066 3238 109078 3290
rect 109130 3238 109142 3290
rect 109194 3238 109206 3290
rect 109258 3238 109270 3290
rect 109322 3238 109334 3290
rect 109386 3238 144822 3290
rect 144874 3238 144886 3290
rect 144938 3238 144950 3290
rect 145002 3238 145014 3290
rect 145066 3238 145078 3290
rect 145130 3238 145142 3290
rect 145194 3238 145206 3290
rect 145258 3238 145270 3290
rect 145322 3238 145334 3290
rect 145386 3238 180822 3290
rect 180874 3238 180886 3290
rect 180938 3238 180950 3290
rect 181002 3238 181014 3290
rect 181066 3238 181078 3290
rect 181130 3238 181142 3290
rect 181194 3238 181206 3290
rect 181258 3238 181270 3290
rect 181322 3238 181334 3290
rect 181386 3238 216822 3290
rect 216874 3238 216886 3290
rect 216938 3238 216950 3290
rect 217002 3238 217014 3290
rect 217066 3238 217078 3290
rect 217130 3238 217142 3290
rect 217194 3238 217206 3290
rect 217258 3238 217270 3290
rect 217322 3238 217334 3290
rect 217386 3238 252822 3290
rect 252874 3238 252886 3290
rect 252938 3238 252950 3290
rect 253002 3238 253014 3290
rect 253066 3238 253078 3290
rect 253130 3238 253142 3290
rect 253194 3238 253206 3290
rect 253258 3238 253270 3290
rect 253322 3238 253334 3290
rect 253386 3238 288822 3290
rect 288874 3238 288886 3290
rect 288938 3238 288950 3290
rect 289002 3238 289014 3290
rect 289066 3238 289078 3290
rect 289130 3238 289142 3290
rect 289194 3238 289206 3290
rect 289258 3238 289270 3290
rect 289322 3238 289334 3290
rect 289386 3238 324822 3290
rect 324874 3238 324886 3290
rect 324938 3238 324950 3290
rect 325002 3238 325014 3290
rect 325066 3238 325078 3290
rect 325130 3238 325142 3290
rect 325194 3238 325206 3290
rect 325258 3238 325270 3290
rect 325322 3238 325334 3290
rect 325386 3238 360822 3290
rect 360874 3238 360886 3290
rect 360938 3238 360950 3290
rect 361002 3238 361014 3290
rect 361066 3238 361078 3290
rect 361130 3238 361142 3290
rect 361194 3238 361206 3290
rect 361258 3238 361270 3290
rect 361322 3238 361334 3290
rect 361386 3238 396822 3290
rect 396874 3238 396886 3290
rect 396938 3238 396950 3290
rect 397002 3238 397014 3290
rect 397066 3238 397078 3290
rect 397130 3238 397142 3290
rect 397194 3238 397206 3290
rect 397258 3238 397270 3290
rect 397322 3238 397334 3290
rect 397386 3238 432822 3290
rect 432874 3238 432886 3290
rect 432938 3238 432950 3290
rect 433002 3238 433014 3290
rect 433066 3238 433078 3290
rect 433130 3238 433142 3290
rect 433194 3238 433206 3290
rect 433258 3238 433270 3290
rect 433322 3238 433334 3290
rect 433386 3238 468822 3290
rect 468874 3238 468886 3290
rect 468938 3238 468950 3290
rect 469002 3238 469014 3290
rect 469066 3238 469078 3290
rect 469130 3238 469142 3290
rect 469194 3238 469206 3290
rect 469258 3238 469270 3290
rect 469322 3238 469334 3290
rect 469386 3238 504822 3290
rect 504874 3238 504886 3290
rect 504938 3238 504950 3290
rect 505002 3238 505014 3290
rect 505066 3238 505078 3290
rect 505130 3238 505142 3290
rect 505194 3238 505206 3290
rect 505258 3238 505270 3290
rect 505322 3238 505334 3290
rect 505386 3238 540822 3290
rect 540874 3238 540886 3290
rect 540938 3238 540950 3290
rect 541002 3238 541014 3290
rect 541066 3238 541078 3290
rect 541130 3238 541142 3290
rect 541194 3238 541206 3290
rect 541258 3238 541270 3290
rect 541322 3238 541334 3290
rect 541386 3238 576822 3290
rect 576874 3238 576886 3290
rect 576938 3238 576950 3290
rect 577002 3238 577014 3290
rect 577066 3238 577078 3290
rect 577130 3238 577142 3290
rect 577194 3238 577206 3290
rect 577258 3238 577270 3290
rect 577322 3238 577334 3290
rect 577386 3238 582820 3290
rect 1104 3216 582820 3238
rect 23106 3136 23112 3188
rect 23164 3176 23170 3188
rect 28258 3176 28264 3188
rect 23164 3148 28264 3176
rect 23164 3136 23170 3148
rect 28258 3136 28264 3148
rect 28316 3136 28322 3188
rect 45738 3136 45744 3188
rect 45796 3176 45802 3188
rect 52086 3176 52092 3188
rect 45796 3148 52092 3176
rect 45796 3136 45802 3148
rect 52086 3136 52092 3148
rect 52144 3136 52150 3188
rect 65978 3136 65984 3188
rect 66036 3176 66042 3188
rect 71498 3176 71504 3188
rect 66036 3148 71504 3176
rect 66036 3136 66042 3148
rect 71498 3136 71504 3148
rect 71556 3136 71562 3188
rect 75454 3136 75460 3188
rect 75512 3176 75518 3188
rect 80698 3176 80704 3188
rect 75512 3148 80704 3176
rect 75512 3136 75518 3148
rect 80698 3136 80704 3148
rect 80756 3136 80762 3188
rect 309134 3136 309140 3188
rect 309192 3176 309198 3188
rect 310974 3176 310980 3188
rect 309192 3148 310980 3176
rect 309192 3136 309198 3148
rect 310974 3136 310980 3148
rect 311032 3136 311038 3188
rect 330110 3136 330116 3188
rect 330168 3176 330174 3188
rect 332410 3176 332416 3188
rect 330168 3148 332416 3176
rect 330168 3136 330174 3148
rect 332410 3136 332416 3148
rect 332468 3136 332474 3188
rect 349982 3136 349988 3188
rect 350040 3176 350046 3188
rect 352558 3176 352564 3188
rect 350040 3148 352564 3176
rect 350040 3136 350046 3148
rect 352558 3136 352564 3148
rect 352616 3136 352622 3188
rect 368658 3136 368664 3188
rect 368716 3176 368722 3188
rect 371602 3176 371608 3188
rect 368716 3148 371608 3176
rect 368716 3136 368722 3148
rect 371602 3136 371608 3148
rect 371660 3136 371666 3188
rect 376662 3136 376668 3188
rect 376720 3176 376726 3188
rect 379974 3176 379980 3188
rect 376720 3148 379980 3176
rect 376720 3136 376726 3148
rect 379974 3136 379980 3148
rect 380032 3136 380038 3188
rect 405642 3136 405648 3188
rect 405700 3176 405706 3188
rect 409690 3176 409696 3188
rect 405700 3148 409696 3176
rect 405700 3136 405706 3148
rect 409690 3136 409696 3148
rect 409748 3136 409754 3188
rect 423582 3136 423588 3188
rect 423640 3176 423646 3188
rect 427538 3176 427544 3188
rect 423640 3148 427544 3176
rect 423640 3136 423646 3148
rect 427538 3136 427544 3148
rect 427596 3136 427602 3188
rect 445846 3136 445852 3188
rect 445904 3176 445910 3188
rect 452470 3176 452476 3188
rect 445904 3148 452476 3176
rect 445904 3136 445910 3148
rect 452470 3136 452476 3148
rect 452528 3136 452534 3188
rect 463602 3136 463608 3188
rect 463660 3176 463666 3188
rect 468662 3176 468668 3188
rect 463660 3148 468668 3176
rect 463660 3136 463666 3148
rect 468662 3136 468668 3148
rect 468720 3136 468726 3188
rect 510982 3136 510988 3188
rect 511040 3176 511046 3188
rect 513190 3176 513196 3188
rect 511040 3148 513196 3176
rect 511040 3136 511046 3148
rect 513190 3136 513196 3148
rect 513248 3136 513254 3188
rect 524414 3136 524420 3188
rect 524472 3176 524478 3188
rect 526254 3176 526260 3188
rect 524472 3148 526260 3176
rect 524472 3136 524478 3148
rect 526254 3136 526260 3148
rect 526312 3136 526318 3188
rect 541434 3136 541440 3188
rect 541492 3176 541498 3188
rect 544102 3176 544108 3188
rect 541492 3148 544108 3176
rect 541492 3136 541498 3148
rect 544102 3136 544108 3148
rect 544160 3136 544166 3188
rect 550634 3136 550640 3188
rect 550692 3176 550698 3188
rect 552382 3176 552388 3188
rect 550692 3148 552388 3176
rect 550692 3136 550698 3148
rect 552382 3136 552388 3148
rect 552440 3136 552446 3188
rect 554866 3136 554872 3188
rect 554924 3176 554930 3188
rect 557166 3176 557172 3188
rect 554924 3148 557172 3176
rect 554924 3136 554930 3148
rect 557166 3136 557172 3148
rect 557224 3136 557230 3188
rect 561674 3136 561680 3188
rect 561732 3176 561738 3188
rect 565538 3176 565544 3188
rect 561732 3148 565544 3176
rect 561732 3136 561738 3148
rect 565538 3136 565544 3148
rect 565596 3136 565602 3188
rect 575474 3136 575480 3188
rect 575532 3176 575538 3188
rect 577406 3176 577412 3188
rect 575532 3148 577412 3176
rect 575532 3136 575538 3148
rect 577406 3136 577412 3148
rect 577464 3136 577470 3188
rect 577682 3136 577688 3188
rect 577740 3176 577746 3188
rect 578602 3176 578608 3188
rect 577740 3148 578608 3176
rect 577740 3136 577746 3148
rect 578602 3136 578608 3148
rect 578660 3136 578666 3188
rect 12434 3068 12440 3120
rect 12492 3108 12498 3120
rect 18322 3108 18328 3120
rect 12492 3080 18328 3108
rect 12492 3068 12498 3080
rect 18322 3068 18328 3080
rect 18380 3068 18386 3120
rect 32674 3068 32680 3120
rect 32732 3108 32738 3120
rect 37642 3108 37648 3120
rect 32732 3080 37648 3108
rect 32732 3068 32738 3080
rect 37642 3068 37648 3080
rect 37700 3068 37706 3120
rect 42150 3068 42156 3120
rect 42208 3108 42214 3120
rect 48222 3108 48228 3120
rect 42208 3080 48228 3108
rect 42208 3068 42214 3080
rect 48222 3068 48228 3080
rect 48280 3068 48286 3120
rect 346118 3068 346124 3120
rect 346176 3108 346182 3120
rect 347866 3108 347872 3120
rect 346176 3080 347872 3108
rect 346176 3068 346182 3080
rect 347866 3068 347872 3080
rect 347924 3068 347930 3120
rect 351086 3068 351092 3120
rect 351144 3108 351150 3120
rect 353754 3108 353760 3120
rect 351144 3080 353760 3108
rect 351144 3068 351150 3080
rect 353754 3068 353760 3080
rect 353812 3068 353818 3120
rect 426434 3068 426440 3120
rect 426492 3108 426498 3120
rect 432322 3108 432328 3120
rect 426492 3080 432328 3108
rect 426492 3068 426498 3080
rect 432322 3068 432328 3080
rect 432380 3068 432386 3120
rect 455414 3068 455420 3120
rect 455472 3108 455478 3120
rect 462038 3108 462044 3120
rect 455472 3080 462044 3108
rect 455472 3068 455478 3080
rect 462038 3068 462044 3080
rect 462096 3068 462102 3120
rect 490742 3068 490748 3120
rect 490800 3108 490806 3120
rect 497734 3108 497740 3120
rect 490800 3080 497740 3108
rect 490800 3068 490806 3080
rect 497734 3068 497740 3080
rect 497792 3068 497798 3120
rect 539962 3068 539968 3120
rect 540020 3108 540026 3120
rect 541710 3108 541716 3120
rect 540020 3080 541716 3108
rect 540020 3068 540026 3080
rect 541710 3068 541716 3080
rect 541768 3068 541774 3120
rect 552014 3068 552020 3120
rect 552072 3108 552078 3120
rect 554774 3108 554780 3120
rect 552072 3080 554780 3108
rect 552072 3068 552078 3080
rect 554774 3068 554780 3080
rect 554832 3068 554838 3120
rect 561766 3068 561772 3120
rect 561824 3108 561830 3120
rect 564342 3108 564348 3120
rect 561824 3080 564348 3108
rect 561824 3068 561830 3080
rect 564342 3068 564348 3080
rect 564400 3068 564406 3120
rect 564618 3068 564624 3120
rect 564676 3108 564682 3120
rect 566734 3108 566740 3120
rect 564676 3080 566740 3108
rect 564676 3068 564682 3080
rect 566734 3068 566740 3080
rect 566792 3068 566798 3120
rect 1670 3000 1676 3052
rect 1728 3040 1734 3052
rect 9582 3040 9588 3052
rect 1728 3012 9588 3040
rect 1728 3000 1734 3012
rect 9582 3000 9588 3012
rect 9640 3000 9646 3052
rect 19518 3000 19524 3052
rect 19576 3040 19582 3052
rect 26142 3040 26148 3052
rect 19576 3012 26148 3040
rect 19576 3000 19582 3012
rect 26142 3000 26148 3012
rect 26200 3000 26206 3052
rect 326522 3000 326528 3052
rect 326580 3040 326586 3052
rect 327626 3040 327632 3052
rect 326580 3012 327632 3040
rect 326580 3000 326586 3012
rect 327626 3000 327632 3012
rect 327684 3000 327690 3052
rect 365622 3000 365628 3052
rect 365680 3040 365686 3052
rect 368014 3040 368020 3052
rect 365680 3012 368020 3040
rect 365680 3000 365686 3012
rect 368014 3000 368020 3012
rect 368072 3000 368078 3052
rect 386138 3000 386144 3052
rect 386196 3040 386202 3052
rect 389450 3040 389456 3052
rect 386196 3012 389456 3040
rect 386196 3000 386202 3012
rect 389450 3000 389456 3012
rect 389508 3000 389514 3052
rect 413738 3000 413744 3052
rect 413796 3040 413802 3052
rect 417970 3040 417976 3052
rect 413796 3012 417976 3040
rect 413796 3000 413802 3012
rect 417970 3000 417976 3012
rect 418028 3000 418034 3052
rect 434162 3000 434168 3052
rect 434220 3040 434226 3052
rect 439406 3040 439412 3052
rect 434220 3012 439412 3040
rect 434220 3000 434226 3012
rect 439406 3000 439412 3012
rect 439464 3000 439470 3052
rect 455322 3000 455328 3052
rect 455380 3040 455386 3052
rect 460842 3040 460848 3052
rect 455380 3012 460848 3040
rect 455380 3000 455386 3012
rect 460842 3000 460848 3012
rect 460900 3000 460906 3052
rect 525794 3000 525800 3052
rect 525852 3040 525858 3052
rect 528646 3040 528652 3052
rect 525852 3012 528652 3040
rect 525852 3000 525858 3012
rect 528646 3000 528652 3012
rect 528704 3000 528710 3052
rect 531498 3000 531504 3052
rect 531556 3040 531562 3052
rect 534534 3040 534540 3052
rect 531556 3012 534540 3040
rect 531556 3000 531562 3012
rect 534534 3000 534540 3012
rect 534592 3000 534598 3052
rect 564526 3000 564532 3052
rect 564584 3040 564590 3052
rect 569034 3040 569040 3052
rect 564584 3012 569040 3040
rect 564584 3000 564590 3012
rect 569034 3000 569040 3012
rect 569092 3000 569098 3052
rect 8846 2932 8852 2984
rect 8904 2972 8910 2984
rect 13814 2972 13820 2984
rect 8904 2944 13820 2972
rect 8904 2932 8910 2944
rect 13814 2932 13820 2944
rect 13872 2932 13878 2984
rect 18322 2932 18328 2984
rect 18380 2972 18386 2984
rect 23474 2972 23480 2984
rect 18380 2944 23480 2972
rect 18380 2932 18386 2944
rect 23474 2932 23480 2944
rect 23532 2932 23538 2984
rect 84930 2932 84936 2984
rect 84988 2972 84994 2984
rect 89806 2972 89812 2984
rect 84988 2944 89812 2972
rect 84988 2932 84994 2944
rect 89806 2932 89812 2944
rect 89864 2932 89870 2984
rect 336642 2932 336648 2984
rect 336700 2972 336706 2984
rect 338298 2972 338304 2984
rect 336700 2944 338304 2972
rect 336700 2932 336706 2944
rect 338298 2932 338304 2944
rect 338356 2932 338362 2984
rect 424502 2932 424508 2984
rect 424560 2972 424566 2984
rect 429930 2972 429936 2984
rect 424560 2944 429936 2972
rect 424560 2932 424566 2944
rect 429930 2932 429936 2944
rect 429988 2932 429994 2984
rect 443822 2932 443828 2984
rect 443880 2972 443886 2984
rect 448974 2972 448980 2984
rect 443880 2944 448980 2972
rect 443880 2932 443886 2944
rect 448974 2932 448980 2944
rect 449032 2932 449038 2984
rect 2866 2864 2872 2916
rect 2924 2904 2930 2916
rect 5534 2904 5540 2916
rect 2924 2876 5540 2904
rect 2924 2864 2930 2876
rect 5534 2864 5540 2876
rect 5592 2864 5598 2916
rect 10042 2864 10048 2916
rect 10100 2904 10106 2916
rect 15194 2904 15200 2916
rect 10100 2876 15200 2904
rect 10100 2864 10106 2876
rect 15194 2864 15200 2876
rect 15252 2864 15258 2916
rect 21910 2864 21916 2916
rect 21968 2904 21974 2916
rect 26602 2904 26608 2916
rect 21968 2876 26608 2904
rect 21968 2864 21974 2876
rect 26602 2864 26608 2876
rect 26660 2864 26666 2916
rect 29086 2864 29092 2916
rect 29144 2904 29150 2916
rect 35802 2904 35808 2916
rect 29144 2876 35808 2904
rect 29144 2864 29150 2876
rect 35802 2864 35808 2876
rect 35860 2864 35866 2916
rect 327166 2864 327172 2916
rect 327224 2904 327230 2916
rect 328822 2904 328828 2916
rect 327224 2876 328828 2904
rect 327224 2864 327230 2876
rect 328822 2864 328828 2876
rect 328880 2864 328886 2916
rect 337286 2864 337292 2916
rect 337344 2904 337350 2916
rect 339494 2904 339500 2916
rect 337344 2876 339500 2904
rect 337344 2864 337350 2876
rect 339494 2864 339500 2876
rect 339552 2864 339558 2916
rect 357250 2864 357256 2916
rect 357308 2904 357314 2916
rect 359734 2904 359740 2916
rect 357308 2876 359740 2904
rect 357308 2864 357314 2876
rect 359734 2864 359740 2876
rect 359792 2864 359798 2916
rect 395338 2864 395344 2916
rect 395396 2904 395402 2916
rect 399018 2904 399024 2916
rect 395396 2876 399024 2904
rect 395396 2864 395402 2876
rect 399018 2864 399024 2876
rect 399076 2864 399082 2916
rect 423306 2864 423312 2916
rect 423364 2904 423370 2916
rect 428734 2904 428740 2916
rect 423364 2876 428740 2904
rect 423364 2864 423370 2876
rect 428734 2864 428740 2876
rect 428792 2864 428798 2916
rect 432690 2864 432696 2916
rect 432748 2904 432754 2916
rect 438210 2904 438216 2916
rect 432748 2876 438216 2904
rect 432748 2864 432754 2876
rect 438210 2864 438216 2876
rect 438268 2864 438274 2916
rect 443454 2864 443460 2916
rect 443512 2904 443518 2916
rect 450170 2904 450176 2916
rect 443512 2876 450176 2904
rect 443512 2864 443518 2876
rect 450170 2864 450176 2876
rect 450228 2864 450234 2916
rect 13630 2796 13636 2848
rect 13688 2836 13694 2848
rect 18690 2836 18696 2848
rect 13688 2808 18696 2836
rect 13688 2796 13694 2808
rect 18690 2796 18696 2808
rect 18748 2796 18754 2848
rect 30282 2796 30288 2848
rect 30340 2836 30346 2848
rect 34514 2836 34520 2848
rect 30340 2808 34520 2836
rect 30340 2796 30346 2808
rect 34514 2796 34520 2808
rect 34572 2796 34578 2848
rect 39758 2796 39764 2848
rect 39816 2836 39822 2848
rect 44174 2836 44180 2848
rect 39816 2808 44180 2836
rect 39816 2796 39822 2808
rect 44174 2796 44180 2808
rect 44232 2796 44238 2848
rect 49326 2796 49332 2848
rect 49384 2836 49390 2848
rect 53834 2836 53840 2848
rect 49384 2808 53840 2836
rect 49384 2796 49390 2808
rect 53834 2796 53840 2808
rect 53892 2796 53898 2848
rect 317690 2796 317696 2848
rect 317748 2836 317754 2848
rect 319254 2836 319260 2848
rect 317748 2808 319260 2836
rect 317748 2796 317754 2808
rect 319254 2796 319260 2808
rect 319312 2796 319318 2848
rect 346854 2796 346860 2848
rect 346912 2836 346918 2848
rect 349062 2836 349068 2848
rect 346912 2808 349068 2836
rect 346912 2796 346918 2808
rect 349062 2796 349068 2808
rect 349120 2796 349126 2848
rect 355594 2796 355600 2848
rect 355652 2836 355658 2848
rect 357342 2836 357348 2848
rect 355652 2808 357348 2836
rect 355652 2796 355658 2808
rect 357342 2796 357348 2808
rect 357400 2796 357406 2848
rect 414658 2796 414664 2848
rect 414716 2836 414722 2848
rect 419166 2836 419172 2848
rect 414716 2808 419172 2836
rect 414716 2796 414722 2808
rect 419166 2796 419172 2808
rect 419224 2796 419230 2848
rect 1104 2746 582820 2768
rect 1104 2694 18822 2746
rect 18874 2694 18886 2746
rect 18938 2694 18950 2746
rect 19002 2694 19014 2746
rect 19066 2694 19078 2746
rect 19130 2694 19142 2746
rect 19194 2694 19206 2746
rect 19258 2694 19270 2746
rect 19322 2694 19334 2746
rect 19386 2694 54822 2746
rect 54874 2694 54886 2746
rect 54938 2694 54950 2746
rect 55002 2694 55014 2746
rect 55066 2694 55078 2746
rect 55130 2694 55142 2746
rect 55194 2694 55206 2746
rect 55258 2694 55270 2746
rect 55322 2694 55334 2746
rect 55386 2694 90822 2746
rect 90874 2694 90886 2746
rect 90938 2694 90950 2746
rect 91002 2694 91014 2746
rect 91066 2694 91078 2746
rect 91130 2694 91142 2746
rect 91194 2694 91206 2746
rect 91258 2694 91270 2746
rect 91322 2694 91334 2746
rect 91386 2694 126822 2746
rect 126874 2694 126886 2746
rect 126938 2694 126950 2746
rect 127002 2694 127014 2746
rect 127066 2694 127078 2746
rect 127130 2694 127142 2746
rect 127194 2694 127206 2746
rect 127258 2694 127270 2746
rect 127322 2694 127334 2746
rect 127386 2694 162822 2746
rect 162874 2694 162886 2746
rect 162938 2694 162950 2746
rect 163002 2694 163014 2746
rect 163066 2694 163078 2746
rect 163130 2694 163142 2746
rect 163194 2694 163206 2746
rect 163258 2694 163270 2746
rect 163322 2694 163334 2746
rect 163386 2694 198822 2746
rect 198874 2694 198886 2746
rect 198938 2694 198950 2746
rect 199002 2694 199014 2746
rect 199066 2694 199078 2746
rect 199130 2694 199142 2746
rect 199194 2694 199206 2746
rect 199258 2694 199270 2746
rect 199322 2694 199334 2746
rect 199386 2694 234822 2746
rect 234874 2694 234886 2746
rect 234938 2694 234950 2746
rect 235002 2694 235014 2746
rect 235066 2694 235078 2746
rect 235130 2694 235142 2746
rect 235194 2694 235206 2746
rect 235258 2694 235270 2746
rect 235322 2694 235334 2746
rect 235386 2694 270822 2746
rect 270874 2694 270886 2746
rect 270938 2694 270950 2746
rect 271002 2694 271014 2746
rect 271066 2694 271078 2746
rect 271130 2694 271142 2746
rect 271194 2694 271206 2746
rect 271258 2694 271270 2746
rect 271322 2694 271334 2746
rect 271386 2694 306822 2746
rect 306874 2694 306886 2746
rect 306938 2694 306950 2746
rect 307002 2694 307014 2746
rect 307066 2694 307078 2746
rect 307130 2694 307142 2746
rect 307194 2694 307206 2746
rect 307258 2694 307270 2746
rect 307322 2694 307334 2746
rect 307386 2694 342822 2746
rect 342874 2694 342886 2746
rect 342938 2694 342950 2746
rect 343002 2694 343014 2746
rect 343066 2694 343078 2746
rect 343130 2694 343142 2746
rect 343194 2694 343206 2746
rect 343258 2694 343270 2746
rect 343322 2694 343334 2746
rect 343386 2694 378822 2746
rect 378874 2694 378886 2746
rect 378938 2694 378950 2746
rect 379002 2694 379014 2746
rect 379066 2694 379078 2746
rect 379130 2694 379142 2746
rect 379194 2694 379206 2746
rect 379258 2694 379270 2746
rect 379322 2694 379334 2746
rect 379386 2694 414822 2746
rect 414874 2694 414886 2746
rect 414938 2694 414950 2746
rect 415002 2694 415014 2746
rect 415066 2694 415078 2746
rect 415130 2694 415142 2746
rect 415194 2694 415206 2746
rect 415258 2694 415270 2746
rect 415322 2694 415334 2746
rect 415386 2694 450822 2746
rect 450874 2694 450886 2746
rect 450938 2694 450950 2746
rect 451002 2694 451014 2746
rect 451066 2694 451078 2746
rect 451130 2694 451142 2746
rect 451194 2694 451206 2746
rect 451258 2694 451270 2746
rect 451322 2694 451334 2746
rect 451386 2694 486822 2746
rect 486874 2694 486886 2746
rect 486938 2694 486950 2746
rect 487002 2694 487014 2746
rect 487066 2694 487078 2746
rect 487130 2694 487142 2746
rect 487194 2694 487206 2746
rect 487258 2694 487270 2746
rect 487322 2694 487334 2746
rect 487386 2694 522822 2746
rect 522874 2694 522886 2746
rect 522938 2694 522950 2746
rect 523002 2694 523014 2746
rect 523066 2694 523078 2746
rect 523130 2694 523142 2746
rect 523194 2694 523206 2746
rect 523258 2694 523270 2746
rect 523322 2694 523334 2746
rect 523386 2694 558822 2746
rect 558874 2694 558886 2746
rect 558938 2694 558950 2746
rect 559002 2694 559014 2746
rect 559066 2694 559078 2746
rect 559130 2694 559142 2746
rect 559194 2694 559206 2746
rect 559258 2694 559270 2746
rect 559322 2694 559334 2746
rect 559386 2694 582820 2746
rect 1104 2672 582820 2694
rect 1104 2202 582820 2224
rect 1104 2150 36822 2202
rect 36874 2150 36886 2202
rect 36938 2150 36950 2202
rect 37002 2150 37014 2202
rect 37066 2150 37078 2202
rect 37130 2150 37142 2202
rect 37194 2150 37206 2202
rect 37258 2150 37270 2202
rect 37322 2150 37334 2202
rect 37386 2150 72822 2202
rect 72874 2150 72886 2202
rect 72938 2150 72950 2202
rect 73002 2150 73014 2202
rect 73066 2150 73078 2202
rect 73130 2150 73142 2202
rect 73194 2150 73206 2202
rect 73258 2150 73270 2202
rect 73322 2150 73334 2202
rect 73386 2150 108822 2202
rect 108874 2150 108886 2202
rect 108938 2150 108950 2202
rect 109002 2150 109014 2202
rect 109066 2150 109078 2202
rect 109130 2150 109142 2202
rect 109194 2150 109206 2202
rect 109258 2150 109270 2202
rect 109322 2150 109334 2202
rect 109386 2150 144822 2202
rect 144874 2150 144886 2202
rect 144938 2150 144950 2202
rect 145002 2150 145014 2202
rect 145066 2150 145078 2202
rect 145130 2150 145142 2202
rect 145194 2150 145206 2202
rect 145258 2150 145270 2202
rect 145322 2150 145334 2202
rect 145386 2150 180822 2202
rect 180874 2150 180886 2202
rect 180938 2150 180950 2202
rect 181002 2150 181014 2202
rect 181066 2150 181078 2202
rect 181130 2150 181142 2202
rect 181194 2150 181206 2202
rect 181258 2150 181270 2202
rect 181322 2150 181334 2202
rect 181386 2150 216822 2202
rect 216874 2150 216886 2202
rect 216938 2150 216950 2202
rect 217002 2150 217014 2202
rect 217066 2150 217078 2202
rect 217130 2150 217142 2202
rect 217194 2150 217206 2202
rect 217258 2150 217270 2202
rect 217322 2150 217334 2202
rect 217386 2150 252822 2202
rect 252874 2150 252886 2202
rect 252938 2150 252950 2202
rect 253002 2150 253014 2202
rect 253066 2150 253078 2202
rect 253130 2150 253142 2202
rect 253194 2150 253206 2202
rect 253258 2150 253270 2202
rect 253322 2150 253334 2202
rect 253386 2150 288822 2202
rect 288874 2150 288886 2202
rect 288938 2150 288950 2202
rect 289002 2150 289014 2202
rect 289066 2150 289078 2202
rect 289130 2150 289142 2202
rect 289194 2150 289206 2202
rect 289258 2150 289270 2202
rect 289322 2150 289334 2202
rect 289386 2150 324822 2202
rect 324874 2150 324886 2202
rect 324938 2150 324950 2202
rect 325002 2150 325014 2202
rect 325066 2150 325078 2202
rect 325130 2150 325142 2202
rect 325194 2150 325206 2202
rect 325258 2150 325270 2202
rect 325322 2150 325334 2202
rect 325386 2150 360822 2202
rect 360874 2150 360886 2202
rect 360938 2150 360950 2202
rect 361002 2150 361014 2202
rect 361066 2150 361078 2202
rect 361130 2150 361142 2202
rect 361194 2150 361206 2202
rect 361258 2150 361270 2202
rect 361322 2150 361334 2202
rect 361386 2150 396822 2202
rect 396874 2150 396886 2202
rect 396938 2150 396950 2202
rect 397002 2150 397014 2202
rect 397066 2150 397078 2202
rect 397130 2150 397142 2202
rect 397194 2150 397206 2202
rect 397258 2150 397270 2202
rect 397322 2150 397334 2202
rect 397386 2150 432822 2202
rect 432874 2150 432886 2202
rect 432938 2150 432950 2202
rect 433002 2150 433014 2202
rect 433066 2150 433078 2202
rect 433130 2150 433142 2202
rect 433194 2150 433206 2202
rect 433258 2150 433270 2202
rect 433322 2150 433334 2202
rect 433386 2150 468822 2202
rect 468874 2150 468886 2202
rect 468938 2150 468950 2202
rect 469002 2150 469014 2202
rect 469066 2150 469078 2202
rect 469130 2150 469142 2202
rect 469194 2150 469206 2202
rect 469258 2150 469270 2202
rect 469322 2150 469334 2202
rect 469386 2150 504822 2202
rect 504874 2150 504886 2202
rect 504938 2150 504950 2202
rect 505002 2150 505014 2202
rect 505066 2150 505078 2202
rect 505130 2150 505142 2202
rect 505194 2150 505206 2202
rect 505258 2150 505270 2202
rect 505322 2150 505334 2202
rect 505386 2150 540822 2202
rect 540874 2150 540886 2202
rect 540938 2150 540950 2202
rect 541002 2150 541014 2202
rect 541066 2150 541078 2202
rect 541130 2150 541142 2202
rect 541194 2150 541206 2202
rect 541258 2150 541270 2202
rect 541322 2150 541334 2202
rect 541386 2150 576822 2202
rect 576874 2150 576886 2202
rect 576938 2150 576950 2202
rect 577002 2150 577014 2202
rect 577066 2150 577078 2202
rect 577130 2150 577142 2202
rect 577194 2150 577206 2202
rect 577258 2150 577270 2202
rect 577322 2150 577334 2202
rect 577386 2150 582820 2202
rect 1104 2128 582820 2150
rect 226334 552 226340 604
rect 226392 592 226398 604
rect 226518 592 226524 604
rect 226392 564 226524 592
rect 226392 552 226398 564
rect 226518 552 226524 564
rect 226576 552 226582 604
<< via1 >>
rect 251640 701972 251692 702024
rect 429844 701972 429896 702024
rect 237472 701904 237524 701956
rect 494796 701904 494848 701956
rect 223304 701836 223356 701888
rect 559656 701836 559708 701888
rect 36822 701734 36874 701786
rect 36886 701734 36938 701786
rect 36950 701734 37002 701786
rect 37014 701734 37066 701786
rect 37078 701734 37130 701786
rect 37142 701734 37194 701786
rect 37206 701734 37258 701786
rect 37270 701734 37322 701786
rect 37334 701734 37386 701786
rect 72822 701734 72874 701786
rect 72886 701734 72938 701786
rect 72950 701734 73002 701786
rect 73014 701734 73066 701786
rect 73078 701734 73130 701786
rect 73142 701734 73194 701786
rect 73206 701734 73258 701786
rect 73270 701734 73322 701786
rect 73334 701734 73386 701786
rect 108822 701734 108874 701786
rect 108886 701734 108938 701786
rect 108950 701734 109002 701786
rect 109014 701734 109066 701786
rect 109078 701734 109130 701786
rect 109142 701734 109194 701786
rect 109206 701734 109258 701786
rect 109270 701734 109322 701786
rect 109334 701734 109386 701786
rect 144822 701734 144874 701786
rect 144886 701734 144938 701786
rect 144950 701734 145002 701786
rect 145014 701734 145066 701786
rect 145078 701734 145130 701786
rect 145142 701734 145194 701786
rect 145206 701734 145258 701786
rect 145270 701734 145322 701786
rect 145334 701734 145386 701786
rect 180822 701734 180874 701786
rect 180886 701734 180938 701786
rect 180950 701734 181002 701786
rect 181014 701734 181066 701786
rect 181078 701734 181130 701786
rect 181142 701734 181194 701786
rect 181206 701734 181258 701786
rect 181270 701734 181322 701786
rect 181334 701734 181386 701786
rect 216822 701734 216874 701786
rect 216886 701734 216938 701786
rect 216950 701734 217002 701786
rect 217014 701734 217066 701786
rect 217078 701734 217130 701786
rect 217142 701734 217194 701786
rect 217206 701734 217258 701786
rect 217270 701734 217322 701786
rect 217334 701734 217386 701786
rect 252822 701734 252874 701786
rect 252886 701734 252938 701786
rect 252950 701734 253002 701786
rect 253014 701734 253066 701786
rect 253078 701734 253130 701786
rect 253142 701734 253194 701786
rect 253206 701734 253258 701786
rect 253270 701734 253322 701786
rect 253334 701734 253386 701786
rect 288822 701734 288874 701786
rect 288886 701734 288938 701786
rect 288950 701734 289002 701786
rect 289014 701734 289066 701786
rect 289078 701734 289130 701786
rect 289142 701734 289194 701786
rect 289206 701734 289258 701786
rect 289270 701734 289322 701786
rect 289334 701734 289386 701786
rect 324822 701734 324874 701786
rect 324886 701734 324938 701786
rect 324950 701734 325002 701786
rect 325014 701734 325066 701786
rect 325078 701734 325130 701786
rect 325142 701734 325194 701786
rect 325206 701734 325258 701786
rect 325270 701734 325322 701786
rect 325334 701734 325386 701786
rect 360822 701734 360874 701786
rect 360886 701734 360938 701786
rect 360950 701734 361002 701786
rect 361014 701734 361066 701786
rect 361078 701734 361130 701786
rect 361142 701734 361194 701786
rect 361206 701734 361258 701786
rect 361270 701734 361322 701786
rect 361334 701734 361386 701786
rect 396822 701734 396874 701786
rect 396886 701734 396938 701786
rect 396950 701734 397002 701786
rect 397014 701734 397066 701786
rect 397078 701734 397130 701786
rect 397142 701734 397194 701786
rect 397206 701734 397258 701786
rect 397270 701734 397322 701786
rect 397334 701734 397386 701786
rect 432822 701734 432874 701786
rect 432886 701734 432938 701786
rect 432950 701734 433002 701786
rect 433014 701734 433066 701786
rect 433078 701734 433130 701786
rect 433142 701734 433194 701786
rect 433206 701734 433258 701786
rect 433270 701734 433322 701786
rect 433334 701734 433386 701786
rect 468822 701734 468874 701786
rect 468886 701734 468938 701786
rect 468950 701734 469002 701786
rect 469014 701734 469066 701786
rect 469078 701734 469130 701786
rect 469142 701734 469194 701786
rect 469206 701734 469258 701786
rect 469270 701734 469322 701786
rect 469334 701734 469386 701786
rect 504822 701734 504874 701786
rect 504886 701734 504938 701786
rect 504950 701734 505002 701786
rect 505014 701734 505066 701786
rect 505078 701734 505130 701786
rect 505142 701734 505194 701786
rect 505206 701734 505258 701786
rect 505270 701734 505322 701786
rect 505334 701734 505386 701786
rect 540822 701734 540874 701786
rect 540886 701734 540938 701786
rect 540950 701734 541002 701786
rect 541014 701734 541066 701786
rect 541078 701734 541130 701786
rect 541142 701734 541194 701786
rect 541206 701734 541258 701786
rect 541270 701734 541322 701786
rect 541334 701734 541386 701786
rect 576822 701734 576874 701786
rect 576886 701734 576938 701786
rect 576950 701734 577002 701786
rect 577014 701734 577066 701786
rect 577078 701734 577130 701786
rect 577142 701734 577194 701786
rect 577206 701734 577258 701786
rect 577270 701734 577322 701786
rect 577334 701734 577386 701786
rect 235172 701632 235224 701684
rect 18822 701190 18874 701242
rect 18886 701190 18938 701242
rect 18950 701190 19002 701242
rect 19014 701190 19066 701242
rect 19078 701190 19130 701242
rect 19142 701190 19194 701242
rect 19206 701190 19258 701242
rect 19270 701190 19322 701242
rect 19334 701190 19386 701242
rect 54822 701190 54874 701242
rect 54886 701190 54938 701242
rect 54950 701190 55002 701242
rect 55014 701190 55066 701242
rect 55078 701190 55130 701242
rect 55142 701190 55194 701242
rect 55206 701190 55258 701242
rect 55270 701190 55322 701242
rect 55334 701190 55386 701242
rect 90822 701190 90874 701242
rect 90886 701190 90938 701242
rect 90950 701190 91002 701242
rect 91014 701190 91066 701242
rect 91078 701190 91130 701242
rect 91142 701190 91194 701242
rect 91206 701190 91258 701242
rect 91270 701190 91322 701242
rect 91334 701190 91386 701242
rect 126822 701190 126874 701242
rect 126886 701190 126938 701242
rect 126950 701190 127002 701242
rect 127014 701190 127066 701242
rect 127078 701190 127130 701242
rect 127142 701190 127194 701242
rect 127206 701190 127258 701242
rect 127270 701190 127322 701242
rect 127334 701190 127386 701242
rect 162822 701190 162874 701242
rect 162886 701190 162938 701242
rect 162950 701190 163002 701242
rect 163014 701190 163066 701242
rect 163078 701190 163130 701242
rect 163142 701190 163194 701242
rect 163206 701190 163258 701242
rect 163270 701190 163322 701242
rect 163334 701190 163386 701242
rect 198822 701190 198874 701242
rect 198886 701190 198938 701242
rect 198950 701190 199002 701242
rect 199014 701190 199066 701242
rect 199078 701190 199130 701242
rect 199142 701190 199194 701242
rect 199206 701190 199258 701242
rect 199270 701190 199322 701242
rect 199334 701190 199386 701242
rect 234822 701190 234874 701242
rect 234886 701190 234938 701242
rect 234950 701190 235002 701242
rect 235014 701190 235066 701242
rect 235078 701190 235130 701242
rect 235142 701190 235194 701242
rect 235206 701190 235258 701242
rect 235270 701190 235322 701242
rect 235334 701190 235386 701242
rect 270822 701190 270874 701242
rect 270886 701190 270938 701242
rect 270950 701190 271002 701242
rect 271014 701190 271066 701242
rect 271078 701190 271130 701242
rect 271142 701190 271194 701242
rect 271206 701190 271258 701242
rect 271270 701190 271322 701242
rect 271334 701190 271386 701242
rect 306822 701190 306874 701242
rect 306886 701190 306938 701242
rect 306950 701190 307002 701242
rect 307014 701190 307066 701242
rect 307078 701190 307130 701242
rect 307142 701190 307194 701242
rect 307206 701190 307258 701242
rect 307270 701190 307322 701242
rect 307334 701190 307386 701242
rect 342822 701190 342874 701242
rect 342886 701190 342938 701242
rect 342950 701190 343002 701242
rect 343014 701190 343066 701242
rect 343078 701190 343130 701242
rect 343142 701190 343194 701242
rect 343206 701190 343258 701242
rect 343270 701190 343322 701242
rect 343334 701190 343386 701242
rect 378822 701190 378874 701242
rect 378886 701190 378938 701242
rect 378950 701190 379002 701242
rect 379014 701190 379066 701242
rect 379078 701190 379130 701242
rect 379142 701190 379194 701242
rect 379206 701190 379258 701242
rect 379270 701190 379322 701242
rect 379334 701190 379386 701242
rect 414822 701190 414874 701242
rect 414886 701190 414938 701242
rect 414950 701190 415002 701242
rect 415014 701190 415066 701242
rect 415078 701190 415130 701242
rect 415142 701190 415194 701242
rect 415206 701190 415258 701242
rect 415270 701190 415322 701242
rect 415334 701190 415386 701242
rect 450822 701190 450874 701242
rect 450886 701190 450938 701242
rect 450950 701190 451002 701242
rect 451014 701190 451066 701242
rect 451078 701190 451130 701242
rect 451142 701190 451194 701242
rect 451206 701190 451258 701242
rect 451270 701190 451322 701242
rect 451334 701190 451386 701242
rect 486822 701190 486874 701242
rect 486886 701190 486938 701242
rect 486950 701190 487002 701242
rect 487014 701190 487066 701242
rect 487078 701190 487130 701242
rect 487142 701190 487194 701242
rect 487206 701190 487258 701242
rect 487270 701190 487322 701242
rect 487334 701190 487386 701242
rect 522822 701190 522874 701242
rect 522886 701190 522938 701242
rect 522950 701190 523002 701242
rect 523014 701190 523066 701242
rect 523078 701190 523130 701242
rect 523142 701190 523194 701242
rect 523206 701190 523258 701242
rect 523270 701190 523322 701242
rect 523334 701190 523386 701242
rect 558822 701190 558874 701242
rect 558886 701190 558938 701242
rect 558950 701190 559002 701242
rect 559014 701190 559066 701242
rect 559078 701190 559130 701242
rect 559142 701190 559194 701242
rect 559206 701190 559258 701242
rect 559270 701190 559322 701242
rect 559334 701190 559386 701242
rect 256424 700952 256476 701004
rect 397460 700952 397512 701004
rect 154120 700884 154172 700936
rect 317972 700884 318024 700936
rect 137836 700816 137888 700868
rect 313188 700816 313240 700868
rect 105452 700748 105504 700800
rect 322664 700748 322716 700800
rect 36822 700646 36874 700698
rect 36886 700646 36938 700698
rect 36950 700646 37002 700698
rect 37014 700646 37066 700698
rect 37078 700646 37130 700698
rect 37142 700646 37194 700698
rect 37206 700646 37258 700698
rect 37270 700646 37322 700698
rect 37334 700646 37386 700698
rect 72822 700646 72874 700698
rect 72886 700646 72938 700698
rect 72950 700646 73002 700698
rect 73014 700646 73066 700698
rect 73078 700646 73130 700698
rect 73142 700646 73194 700698
rect 73206 700646 73258 700698
rect 73270 700646 73322 700698
rect 73334 700646 73386 700698
rect 108822 700646 108874 700698
rect 108886 700646 108938 700698
rect 108950 700646 109002 700698
rect 109014 700646 109066 700698
rect 109078 700646 109130 700698
rect 109142 700646 109194 700698
rect 109206 700646 109258 700698
rect 109270 700646 109322 700698
rect 109334 700646 109386 700698
rect 144822 700646 144874 700698
rect 144886 700646 144938 700698
rect 144950 700646 145002 700698
rect 145014 700646 145066 700698
rect 145078 700646 145130 700698
rect 145142 700646 145194 700698
rect 145206 700646 145258 700698
rect 145270 700646 145322 700698
rect 145334 700646 145386 700698
rect 180822 700646 180874 700698
rect 180886 700646 180938 700698
rect 180950 700646 181002 700698
rect 181014 700646 181066 700698
rect 181078 700646 181130 700698
rect 181142 700646 181194 700698
rect 181206 700646 181258 700698
rect 181270 700646 181322 700698
rect 181334 700646 181386 700698
rect 216822 700646 216874 700698
rect 216886 700646 216938 700698
rect 216950 700646 217002 700698
rect 217014 700646 217066 700698
rect 217078 700646 217130 700698
rect 217142 700646 217194 700698
rect 217206 700646 217258 700698
rect 217270 700646 217322 700698
rect 217334 700646 217386 700698
rect 252822 700646 252874 700698
rect 252886 700646 252938 700698
rect 252950 700646 253002 700698
rect 253014 700646 253066 700698
rect 253078 700646 253130 700698
rect 253142 700646 253194 700698
rect 253206 700646 253258 700698
rect 253270 700646 253322 700698
rect 253334 700646 253386 700698
rect 288822 700646 288874 700698
rect 288886 700646 288938 700698
rect 288950 700646 289002 700698
rect 289014 700646 289066 700698
rect 289078 700646 289130 700698
rect 289142 700646 289194 700698
rect 289206 700646 289258 700698
rect 289270 700646 289322 700698
rect 289334 700646 289386 700698
rect 324822 700646 324874 700698
rect 324886 700646 324938 700698
rect 324950 700646 325002 700698
rect 325014 700646 325066 700698
rect 325078 700646 325130 700698
rect 325142 700646 325194 700698
rect 325206 700646 325258 700698
rect 325270 700646 325322 700698
rect 325334 700646 325386 700698
rect 360822 700646 360874 700698
rect 360886 700646 360938 700698
rect 360950 700646 361002 700698
rect 361014 700646 361066 700698
rect 361078 700646 361130 700698
rect 361142 700646 361194 700698
rect 361206 700646 361258 700698
rect 361270 700646 361322 700698
rect 361334 700646 361386 700698
rect 396822 700646 396874 700698
rect 396886 700646 396938 700698
rect 396950 700646 397002 700698
rect 397014 700646 397066 700698
rect 397078 700646 397130 700698
rect 397142 700646 397194 700698
rect 397206 700646 397258 700698
rect 397270 700646 397322 700698
rect 397334 700646 397386 700698
rect 432822 700646 432874 700698
rect 432886 700646 432938 700698
rect 432950 700646 433002 700698
rect 433014 700646 433066 700698
rect 433078 700646 433130 700698
rect 433142 700646 433194 700698
rect 433206 700646 433258 700698
rect 433270 700646 433322 700698
rect 433334 700646 433386 700698
rect 468822 700646 468874 700698
rect 468886 700646 468938 700698
rect 468950 700646 469002 700698
rect 469014 700646 469066 700698
rect 469078 700646 469130 700698
rect 469142 700646 469194 700698
rect 469206 700646 469258 700698
rect 469270 700646 469322 700698
rect 469334 700646 469386 700698
rect 504822 700646 504874 700698
rect 504886 700646 504938 700698
rect 504950 700646 505002 700698
rect 505014 700646 505066 700698
rect 505078 700646 505130 700698
rect 505142 700646 505194 700698
rect 505206 700646 505258 700698
rect 505270 700646 505322 700698
rect 505334 700646 505386 700698
rect 540822 700646 540874 700698
rect 540886 700646 540938 700698
rect 540950 700646 541002 700698
rect 541014 700646 541066 700698
rect 541078 700646 541130 700698
rect 541142 700646 541194 700698
rect 541206 700646 541258 700698
rect 541270 700646 541322 700698
rect 541334 700646 541386 700698
rect 576822 700646 576874 700698
rect 576886 700646 576938 700698
rect 576950 700646 577002 700698
rect 577014 700646 577066 700698
rect 577078 700646 577130 700698
rect 577142 700646 577194 700698
rect 577206 700646 577258 700698
rect 577270 700646 577322 700698
rect 577334 700646 577386 700698
rect 242256 700544 242308 700596
rect 462320 700544 462372 700596
rect 246948 700476 247000 700528
rect 478512 700476 478564 700528
rect 89168 700408 89220 700460
rect 332140 700408 332192 700460
rect 202788 700340 202840 700392
rect 292580 700340 292632 700392
rect 292672 700340 292724 700392
rect 300124 700340 300176 700392
rect 300216 700340 300268 700392
rect 543464 700340 543516 700392
rect 72700 700272 72752 700324
rect 327448 700272 327500 700324
rect 170312 700204 170364 700256
rect 308496 700204 308548 700256
rect 18822 700102 18874 700154
rect 18886 700102 18938 700154
rect 18950 700102 19002 700154
rect 19014 700102 19066 700154
rect 19078 700102 19130 700154
rect 19142 700102 19194 700154
rect 19206 700102 19258 700154
rect 19270 700102 19322 700154
rect 19334 700102 19386 700154
rect 54822 700102 54874 700154
rect 54886 700102 54938 700154
rect 54950 700102 55002 700154
rect 55014 700102 55066 700154
rect 55078 700102 55130 700154
rect 55142 700102 55194 700154
rect 55206 700102 55258 700154
rect 55270 700102 55322 700154
rect 55334 700102 55386 700154
rect 90822 700102 90874 700154
rect 90886 700102 90938 700154
rect 90950 700102 91002 700154
rect 91014 700102 91066 700154
rect 91078 700102 91130 700154
rect 91142 700102 91194 700154
rect 91206 700102 91258 700154
rect 91270 700102 91322 700154
rect 91334 700102 91386 700154
rect 126822 700102 126874 700154
rect 126886 700102 126938 700154
rect 126950 700102 127002 700154
rect 127014 700102 127066 700154
rect 127078 700102 127130 700154
rect 127142 700102 127194 700154
rect 127206 700102 127258 700154
rect 127270 700102 127322 700154
rect 127334 700102 127386 700154
rect 162822 700102 162874 700154
rect 162886 700102 162938 700154
rect 162950 700102 163002 700154
rect 163014 700102 163066 700154
rect 163078 700102 163130 700154
rect 163142 700102 163194 700154
rect 163206 700102 163258 700154
rect 163270 700102 163322 700154
rect 163334 700102 163386 700154
rect 198822 700102 198874 700154
rect 198886 700102 198938 700154
rect 198950 700102 199002 700154
rect 199014 700102 199066 700154
rect 199078 700102 199130 700154
rect 199142 700102 199194 700154
rect 199206 700102 199258 700154
rect 199270 700102 199322 700154
rect 199334 700102 199386 700154
rect 234822 700102 234874 700154
rect 234886 700102 234938 700154
rect 234950 700102 235002 700154
rect 235014 700102 235066 700154
rect 235078 700102 235130 700154
rect 235142 700102 235194 700154
rect 235206 700102 235258 700154
rect 235270 700102 235322 700154
rect 235334 700102 235386 700154
rect 270822 700102 270874 700154
rect 270886 700102 270938 700154
rect 270950 700102 271002 700154
rect 271014 700102 271066 700154
rect 271078 700102 271130 700154
rect 271142 700102 271194 700154
rect 271206 700102 271258 700154
rect 271270 700102 271322 700154
rect 271334 700102 271386 700154
rect 306822 700102 306874 700154
rect 306886 700102 306938 700154
rect 306950 700102 307002 700154
rect 307014 700102 307066 700154
rect 307078 700102 307130 700154
rect 307142 700102 307194 700154
rect 307206 700102 307258 700154
rect 307270 700102 307322 700154
rect 307334 700102 307386 700154
rect 342822 700102 342874 700154
rect 342886 700102 342938 700154
rect 342950 700102 343002 700154
rect 343014 700102 343066 700154
rect 343078 700102 343130 700154
rect 343142 700102 343194 700154
rect 343206 700102 343258 700154
rect 343270 700102 343322 700154
rect 343334 700102 343386 700154
rect 378822 700102 378874 700154
rect 378886 700102 378938 700154
rect 378950 700102 379002 700154
rect 379014 700102 379066 700154
rect 379078 700102 379130 700154
rect 379142 700102 379194 700154
rect 379206 700102 379258 700154
rect 379270 700102 379322 700154
rect 379334 700102 379386 700154
rect 414822 700102 414874 700154
rect 414886 700102 414938 700154
rect 414950 700102 415002 700154
rect 415014 700102 415066 700154
rect 415078 700102 415130 700154
rect 415142 700102 415194 700154
rect 415206 700102 415258 700154
rect 415270 700102 415322 700154
rect 415334 700102 415386 700154
rect 450822 700102 450874 700154
rect 450886 700102 450938 700154
rect 450950 700102 451002 700154
rect 451014 700102 451066 700154
rect 451078 700102 451130 700154
rect 451142 700102 451194 700154
rect 451206 700102 451258 700154
rect 451270 700102 451322 700154
rect 451334 700102 451386 700154
rect 486822 700102 486874 700154
rect 486886 700102 486938 700154
rect 486950 700102 487002 700154
rect 487014 700102 487066 700154
rect 487078 700102 487130 700154
rect 487142 700102 487194 700154
rect 487206 700102 487258 700154
rect 487270 700102 487322 700154
rect 487334 700102 487386 700154
rect 522822 700102 522874 700154
rect 522886 700102 522938 700154
rect 522950 700102 523002 700154
rect 523014 700102 523066 700154
rect 523078 700102 523130 700154
rect 523142 700102 523194 700154
rect 523206 700102 523258 700154
rect 523270 700102 523322 700154
rect 523334 700102 523386 700154
rect 558822 700102 558874 700154
rect 558886 700102 558938 700154
rect 558950 700102 559002 700154
rect 559014 700102 559066 700154
rect 559078 700102 559130 700154
rect 559142 700102 559194 700154
rect 559206 700102 559258 700154
rect 559270 700102 559322 700154
rect 559334 700102 559386 700154
rect 267648 700000 267700 700052
rect 283748 700000 283800 700052
rect 283840 700000 283892 700052
rect 289452 700000 289504 700052
rect 289544 700000 289596 700052
rect 413652 700000 413704 700052
rect 244188 699932 244240 699984
rect 251088 699932 251140 699984
rect 253848 699932 253900 699984
rect 265900 699932 265952 699984
rect 364984 699932 365036 699984
rect 218980 699864 219032 699916
rect 302056 699864 302108 699916
rect 241520 699728 241572 699780
rect 251088 699728 251140 699780
rect 270500 699796 270552 699848
rect 270592 699796 270644 699848
rect 263876 699728 263928 699780
rect 273536 699728 273588 699780
rect 275744 699728 275796 699780
rect 292488 699796 292540 699848
rect 301964 699796 302016 699848
rect 292304 699728 292356 699780
rect 292672 699728 292724 699780
rect 340788 699864 340840 699916
rect 348792 699796 348844 699848
rect 179328 699660 179380 699712
rect 273168 699660 273220 699712
rect 282920 699660 282972 699712
rect 288440 699660 288492 699712
rect 292580 699660 292632 699712
rect 311900 699660 311952 699712
rect 332508 699728 332560 699780
rect 331220 699660 331272 699712
rect 343548 699660 343600 699712
rect 374000 699660 374052 699712
rect 36822 699558 36874 699610
rect 36886 699558 36938 699610
rect 36950 699558 37002 699610
rect 37014 699558 37066 699610
rect 37078 699558 37130 699610
rect 37142 699558 37194 699610
rect 37206 699558 37258 699610
rect 37270 699558 37322 699610
rect 37334 699558 37386 699610
rect 72822 699558 72874 699610
rect 72886 699558 72938 699610
rect 72950 699558 73002 699610
rect 73014 699558 73066 699610
rect 73078 699558 73130 699610
rect 73142 699558 73194 699610
rect 73206 699558 73258 699610
rect 73270 699558 73322 699610
rect 73334 699558 73386 699610
rect 108822 699558 108874 699610
rect 108886 699558 108938 699610
rect 108950 699558 109002 699610
rect 109014 699558 109066 699610
rect 109078 699558 109130 699610
rect 109142 699558 109194 699610
rect 109206 699558 109258 699610
rect 109270 699558 109322 699610
rect 109334 699558 109386 699610
rect 144822 699558 144874 699610
rect 144886 699558 144938 699610
rect 144950 699558 145002 699610
rect 145014 699558 145066 699610
rect 145078 699558 145130 699610
rect 145142 699558 145194 699610
rect 145206 699558 145258 699610
rect 145270 699558 145322 699610
rect 145334 699558 145386 699610
rect 180822 699558 180874 699610
rect 180886 699558 180938 699610
rect 180950 699558 181002 699610
rect 181014 699558 181066 699610
rect 181078 699558 181130 699610
rect 181142 699558 181194 699610
rect 181206 699558 181258 699610
rect 181270 699558 181322 699610
rect 181334 699558 181386 699610
rect 216822 699558 216874 699610
rect 216886 699558 216938 699610
rect 216950 699558 217002 699610
rect 217014 699558 217066 699610
rect 217078 699558 217130 699610
rect 217142 699558 217194 699610
rect 217206 699558 217258 699610
rect 217270 699558 217322 699610
rect 217334 699558 217386 699610
rect 252822 699558 252874 699610
rect 252886 699558 252938 699610
rect 252950 699558 253002 699610
rect 253014 699558 253066 699610
rect 253078 699558 253130 699610
rect 253142 699558 253194 699610
rect 253206 699558 253258 699610
rect 253270 699558 253322 699610
rect 253334 699558 253386 699610
rect 288822 699558 288874 699610
rect 288886 699558 288938 699610
rect 288950 699558 289002 699610
rect 289014 699558 289066 699610
rect 289078 699558 289130 699610
rect 289142 699558 289194 699610
rect 289206 699558 289258 699610
rect 289270 699558 289322 699610
rect 289334 699558 289386 699610
rect 324822 699558 324874 699610
rect 324886 699558 324938 699610
rect 324950 699558 325002 699610
rect 325014 699558 325066 699610
rect 325078 699558 325130 699610
rect 325142 699558 325194 699610
rect 325206 699558 325258 699610
rect 325270 699558 325322 699610
rect 325334 699558 325386 699610
rect 360822 699558 360874 699610
rect 360886 699558 360938 699610
rect 360950 699558 361002 699610
rect 361014 699558 361066 699610
rect 361078 699558 361130 699610
rect 361142 699558 361194 699610
rect 361206 699558 361258 699610
rect 361270 699558 361322 699610
rect 361334 699558 361386 699610
rect 396822 699558 396874 699610
rect 396886 699558 396938 699610
rect 396950 699558 397002 699610
rect 397014 699558 397066 699610
rect 397078 699558 397130 699610
rect 397142 699558 397194 699610
rect 397206 699558 397258 699610
rect 397270 699558 397322 699610
rect 397334 699558 397386 699610
rect 432822 699558 432874 699610
rect 432886 699558 432938 699610
rect 432950 699558 433002 699610
rect 433014 699558 433066 699610
rect 433078 699558 433130 699610
rect 433142 699558 433194 699610
rect 433206 699558 433258 699610
rect 433270 699558 433322 699610
rect 433334 699558 433386 699610
rect 468822 699558 468874 699610
rect 468886 699558 468938 699610
rect 468950 699558 469002 699610
rect 469014 699558 469066 699610
rect 469078 699558 469130 699610
rect 469142 699558 469194 699610
rect 469206 699558 469258 699610
rect 469270 699558 469322 699610
rect 469334 699558 469386 699610
rect 504822 699558 504874 699610
rect 504886 699558 504938 699610
rect 504950 699558 505002 699610
rect 505014 699558 505066 699610
rect 505078 699558 505130 699610
rect 505142 699558 505194 699610
rect 505206 699558 505258 699610
rect 505270 699558 505322 699610
rect 505334 699558 505386 699610
rect 540822 699558 540874 699610
rect 540886 699558 540938 699610
rect 540950 699558 541002 699610
rect 541014 699558 541066 699610
rect 541078 699558 541130 699610
rect 541142 699558 541194 699610
rect 541206 699558 541258 699610
rect 541270 699558 541322 699610
rect 541334 699558 541386 699610
rect 576822 699558 576874 699610
rect 576886 699558 576938 699610
rect 576950 699558 577002 699610
rect 577014 699558 577066 699610
rect 577078 699558 577130 699610
rect 577142 699558 577194 699610
rect 577206 699558 577258 699610
rect 577270 699558 577322 699610
rect 577334 699558 577386 699610
rect 86040 699456 86092 699508
rect 403164 699456 403216 699508
rect 404268 699456 404320 699508
rect 417332 699456 417384 699508
rect 71780 699388 71832 699440
rect 273260 699388 273312 699440
rect 273352 699388 273404 699440
rect 282920 699388 282972 699440
rect 283012 699388 283064 699440
rect 292672 699388 292724 699440
rect 302148 699388 302200 699440
rect 431592 699388 431644 699440
rect 114376 699320 114428 699372
rect 407948 699320 408000 699372
rect 161756 699252 161808 699304
rect 577872 699252 577924 699304
rect 5172 699184 5224 699236
rect 133328 699116 133380 699168
rect 180800 699116 180852 699168
rect 190368 699116 190420 699168
rect 190460 699116 190512 699168
rect 200028 699116 200080 699168
rect 209780 699116 209832 699168
rect 219348 699116 219400 699168
rect 229100 699116 229152 699168
rect 234712 699184 234764 699236
rect 244096 699116 244148 699168
rect 244188 699116 244240 699168
rect 253664 699116 253716 699168
rect 253848 699184 253900 699236
rect 282736 699116 282788 699168
rect 282828 699116 282880 699168
rect 282920 699116 282972 699168
rect 283012 699116 283064 699168
rect 292396 699116 292448 699168
rect 292488 699116 292540 699168
rect 325516 699116 325568 699168
rect 325700 699116 325752 699168
rect 445760 699184 445812 699236
rect 340788 699116 340840 699168
rect 354496 699116 354548 699168
rect 579160 699116 579212 699168
rect 18822 699014 18874 699066
rect 18886 699014 18938 699066
rect 18950 699014 19002 699066
rect 19014 699014 19066 699066
rect 19078 699014 19130 699066
rect 19142 699014 19194 699066
rect 19206 699014 19258 699066
rect 19270 699014 19322 699066
rect 19334 699014 19386 699066
rect 54822 699014 54874 699066
rect 54886 699014 54938 699066
rect 54950 699014 55002 699066
rect 55014 699014 55066 699066
rect 55078 699014 55130 699066
rect 55142 699014 55194 699066
rect 55206 699014 55258 699066
rect 55270 699014 55322 699066
rect 55334 699014 55386 699066
rect 90822 699014 90874 699066
rect 90886 699014 90938 699066
rect 90950 699014 91002 699066
rect 91014 699014 91066 699066
rect 91078 699014 91130 699066
rect 91142 699014 91194 699066
rect 91206 699014 91258 699066
rect 91270 699014 91322 699066
rect 91334 699014 91386 699066
rect 126822 699014 126874 699066
rect 126886 699014 126938 699066
rect 126950 699014 127002 699066
rect 127014 699014 127066 699066
rect 127078 699014 127130 699066
rect 127142 699014 127194 699066
rect 127206 699014 127258 699066
rect 127270 699014 127322 699066
rect 127334 699014 127386 699066
rect 162822 699014 162874 699066
rect 162886 699014 162938 699066
rect 162950 699014 163002 699066
rect 163014 699014 163066 699066
rect 163078 699014 163130 699066
rect 163142 699014 163194 699066
rect 163206 699014 163258 699066
rect 163270 699014 163322 699066
rect 163334 699014 163386 699066
rect 198822 699014 198874 699066
rect 198886 699014 198938 699066
rect 198950 699014 199002 699066
rect 199014 699014 199066 699066
rect 199078 699014 199130 699066
rect 199142 699014 199194 699066
rect 199206 699014 199258 699066
rect 199270 699014 199322 699066
rect 199334 699014 199386 699066
rect 234822 699014 234874 699066
rect 234886 699014 234938 699066
rect 234950 699014 235002 699066
rect 235014 699014 235066 699066
rect 235078 699014 235130 699066
rect 235142 699014 235194 699066
rect 235206 699014 235258 699066
rect 235270 699014 235322 699066
rect 235334 699014 235386 699066
rect 270822 699014 270874 699066
rect 270886 699014 270938 699066
rect 270950 699014 271002 699066
rect 271014 699014 271066 699066
rect 271078 699014 271130 699066
rect 271142 699014 271194 699066
rect 271206 699014 271258 699066
rect 271270 699014 271322 699066
rect 271334 699014 271386 699066
rect 306822 699014 306874 699066
rect 306886 699014 306938 699066
rect 306950 699014 307002 699066
rect 307014 699014 307066 699066
rect 307078 699014 307130 699066
rect 307142 699014 307194 699066
rect 307206 699014 307258 699066
rect 307270 699014 307322 699066
rect 307334 699014 307386 699066
rect 342822 699014 342874 699066
rect 342886 699014 342938 699066
rect 342950 699014 343002 699066
rect 343014 699014 343066 699066
rect 343078 699014 343130 699066
rect 343142 699014 343194 699066
rect 343206 699014 343258 699066
rect 343270 699014 343322 699066
rect 343334 699014 343386 699066
rect 378822 699014 378874 699066
rect 378886 699014 378938 699066
rect 378950 699014 379002 699066
rect 379014 699014 379066 699066
rect 379078 699014 379130 699066
rect 379142 699014 379194 699066
rect 379206 699014 379258 699066
rect 379270 699014 379322 699066
rect 379334 699014 379386 699066
rect 414822 699014 414874 699066
rect 414886 699014 414938 699066
rect 414950 699014 415002 699066
rect 415014 699014 415066 699066
rect 415078 699014 415130 699066
rect 415142 699014 415194 699066
rect 415206 699014 415258 699066
rect 415270 699014 415322 699066
rect 415334 699014 415386 699066
rect 450822 699014 450874 699066
rect 450886 699014 450938 699066
rect 450950 699014 451002 699066
rect 451014 699014 451066 699066
rect 451078 699014 451130 699066
rect 451142 699014 451194 699066
rect 451206 699014 451258 699066
rect 451270 699014 451322 699066
rect 451334 699014 451386 699066
rect 486822 699014 486874 699066
rect 486886 699014 486938 699066
rect 486950 699014 487002 699066
rect 487014 699014 487066 699066
rect 487078 699014 487130 699066
rect 487142 699014 487194 699066
rect 487206 699014 487258 699066
rect 487270 699014 487322 699066
rect 487334 699014 487386 699066
rect 522822 699014 522874 699066
rect 522886 699014 522938 699066
rect 522950 699014 523002 699066
rect 523014 699014 523066 699066
rect 523078 699014 523130 699066
rect 523142 699014 523194 699066
rect 523206 699014 523258 699066
rect 523270 699014 523322 699066
rect 523334 699014 523386 699066
rect 558822 699014 558874 699066
rect 558886 699014 558938 699066
rect 558950 699014 559002 699066
rect 559014 699014 559066 699066
rect 559078 699014 559130 699066
rect 559142 699014 559194 699066
rect 559206 699014 559258 699066
rect 559270 699014 559322 699066
rect 559334 699014 559386 699066
rect 48136 698912 48188 698964
rect 119712 698912 119764 698964
rect 128636 698912 128688 698964
rect 576584 698912 576636 698964
rect 119160 698844 119212 698896
rect 253756 698844 253808 698896
rect 253848 698844 253900 698896
rect 263600 698844 263652 698896
rect 263692 698844 263744 698896
rect 306380 698844 306432 698896
rect 325608 698844 325660 698896
rect 340696 698844 340748 698896
rect 354588 698844 354640 698896
rect 577688 698844 577740 698896
rect 5264 698776 5316 698828
rect 474188 698776 474240 698828
rect 33968 698708 34020 698760
rect 89720 698708 89772 698760
rect 104992 698708 105044 698760
rect 577596 698708 577648 698760
rect 4988 698640 5040 698692
rect 488356 698640 488408 698692
rect 90732 698572 90784 698624
rect 576400 698572 576452 698624
rect 36822 698470 36874 698522
rect 36886 698470 36938 698522
rect 36950 698470 37002 698522
rect 37014 698470 37066 698522
rect 37078 698470 37130 698522
rect 37142 698470 37194 698522
rect 37206 698470 37258 698522
rect 37270 698470 37322 698522
rect 37334 698470 37386 698522
rect 72822 698470 72874 698522
rect 72886 698470 72938 698522
rect 72950 698470 73002 698522
rect 73014 698470 73066 698522
rect 73078 698470 73130 698522
rect 73142 698470 73194 698522
rect 73206 698470 73258 698522
rect 73270 698470 73322 698522
rect 73334 698470 73386 698522
rect 108822 698470 108874 698522
rect 108886 698470 108938 698522
rect 108950 698470 109002 698522
rect 109014 698470 109066 698522
rect 109078 698470 109130 698522
rect 109142 698470 109194 698522
rect 109206 698470 109258 698522
rect 109270 698470 109322 698522
rect 109334 698470 109386 698522
rect 144822 698470 144874 698522
rect 144886 698470 144938 698522
rect 144950 698470 145002 698522
rect 145014 698470 145066 698522
rect 145078 698470 145130 698522
rect 145142 698470 145194 698522
rect 145206 698470 145258 698522
rect 145270 698470 145322 698522
rect 145334 698470 145386 698522
rect 180822 698470 180874 698522
rect 180886 698470 180938 698522
rect 180950 698470 181002 698522
rect 181014 698470 181066 698522
rect 181078 698470 181130 698522
rect 181142 698470 181194 698522
rect 181206 698470 181258 698522
rect 181270 698470 181322 698522
rect 181334 698470 181386 698522
rect 216822 698470 216874 698522
rect 216886 698470 216938 698522
rect 216950 698470 217002 698522
rect 217014 698470 217066 698522
rect 217078 698470 217130 698522
rect 217142 698470 217194 698522
rect 217206 698470 217258 698522
rect 217270 698470 217322 698522
rect 217334 698470 217386 698522
rect 252822 698470 252874 698522
rect 252886 698470 252938 698522
rect 252950 698470 253002 698522
rect 253014 698470 253066 698522
rect 253078 698470 253130 698522
rect 253142 698470 253194 698522
rect 253206 698470 253258 698522
rect 253270 698470 253322 698522
rect 253334 698470 253386 698522
rect 288822 698470 288874 698522
rect 288886 698470 288938 698522
rect 288950 698470 289002 698522
rect 289014 698470 289066 698522
rect 289078 698470 289130 698522
rect 289142 698470 289194 698522
rect 289206 698470 289258 698522
rect 289270 698470 289322 698522
rect 289334 698470 289386 698522
rect 324822 698470 324874 698522
rect 324886 698470 324938 698522
rect 324950 698470 325002 698522
rect 325014 698470 325066 698522
rect 325078 698470 325130 698522
rect 325142 698470 325194 698522
rect 325206 698470 325258 698522
rect 325270 698470 325322 698522
rect 325334 698470 325386 698522
rect 360822 698470 360874 698522
rect 360886 698470 360938 698522
rect 360950 698470 361002 698522
rect 361014 698470 361066 698522
rect 361078 698470 361130 698522
rect 361142 698470 361194 698522
rect 361206 698470 361258 698522
rect 361270 698470 361322 698522
rect 361334 698470 361386 698522
rect 396822 698470 396874 698522
rect 396886 698470 396938 698522
rect 396950 698470 397002 698522
rect 397014 698470 397066 698522
rect 397078 698470 397130 698522
rect 397142 698470 397194 698522
rect 397206 698470 397258 698522
rect 397270 698470 397322 698522
rect 397334 698470 397386 698522
rect 432822 698470 432874 698522
rect 432886 698470 432938 698522
rect 432950 698470 433002 698522
rect 433014 698470 433066 698522
rect 433078 698470 433130 698522
rect 433142 698470 433194 698522
rect 433206 698470 433258 698522
rect 433270 698470 433322 698522
rect 433334 698470 433386 698522
rect 468822 698470 468874 698522
rect 468886 698470 468938 698522
rect 468950 698470 469002 698522
rect 469014 698470 469066 698522
rect 469078 698470 469130 698522
rect 469142 698470 469194 698522
rect 469206 698470 469258 698522
rect 469270 698470 469322 698522
rect 469334 698470 469386 698522
rect 504822 698470 504874 698522
rect 504886 698470 504938 698522
rect 504950 698470 505002 698522
rect 505014 698470 505066 698522
rect 505078 698470 505130 698522
rect 505142 698470 505194 698522
rect 505206 698470 505258 698522
rect 505270 698470 505322 698522
rect 505334 698470 505386 698522
rect 540822 698470 540874 698522
rect 540886 698470 540938 698522
rect 540950 698470 541002 698522
rect 541014 698470 541066 698522
rect 541078 698470 541130 698522
rect 541142 698470 541194 698522
rect 541206 698470 541258 698522
rect 541270 698470 541322 698522
rect 541334 698470 541386 698522
rect 576822 698470 576874 698522
rect 576886 698470 576938 698522
rect 576950 698470 577002 698522
rect 577014 698470 577066 698522
rect 577078 698470 577130 698522
rect 577142 698470 577194 698522
rect 577206 698470 577258 698522
rect 577270 698470 577322 698522
rect 577334 698470 577386 698522
rect 76564 698368 76616 698420
rect 578884 698368 578936 698420
rect 62304 698300 62356 698352
rect 576308 698300 576360 698352
rect 5724 698232 5776 698284
rect 351092 698232 351144 698284
rect 5816 698164 5868 698216
rect 365260 698164 365312 698216
rect 580632 698164 580684 698216
rect 209044 698096 209096 698148
rect 574560 698096 574612 698148
rect 5908 698028 5960 698080
rect 213828 698028 213880 698080
rect 579620 698028 579672 698080
rect 379520 697960 379572 698012
rect 194876 697892 194928 697944
rect 574652 697892 574704 697944
rect 6000 697824 6052 697876
rect 393688 697824 393740 697876
rect 7380 697756 7432 697808
rect 398380 697756 398432 697808
rect 180708 697688 180760 697740
rect 575388 697688 575440 697740
rect 6092 697620 6144 697672
rect 407856 697620 407908 697672
rect 407948 697620 408000 697672
rect 580816 697620 580868 697672
rect 166448 697552 166500 697604
rect 577964 697552 578016 697604
rect 6736 697484 6788 697536
rect 422116 697484 422168 697536
rect 152280 697416 152332 697468
rect 576768 697416 576820 697468
rect 6644 697348 6696 697400
rect 436284 697348 436336 697400
rect 6460 697280 6512 697332
rect 455236 697280 455288 697332
rect 6368 697212 6420 697264
rect 464712 697212 464764 697264
rect 7932 697144 7984 697196
rect 493048 697144 493100 697196
rect 7564 697076 7616 697128
rect 535644 697076 535696 697128
rect 38660 697008 38712 697060
rect 574928 697008 574980 697060
rect 24492 696940 24544 696992
rect 576216 696940 576268 696992
rect 374000 696872 374052 696924
rect 374828 696872 374880 696924
rect 3976 696736 4028 696788
rect 289728 696804 289780 696856
rect 404268 696736 404320 696788
rect 4712 696668 4764 696720
rect 360568 696668 360620 696720
rect 388996 696668 389048 696720
rect 3332 696600 3384 696652
rect 218520 696600 218572 696652
rect 578792 696600 578844 696652
rect 5448 696532 5500 696584
rect 374736 696532 374788 696584
rect 374828 696532 374880 696584
rect 580724 696532 580776 696584
rect 119712 696396 119764 696448
rect 171600 696371 171652 696380
rect 171600 696337 171609 696371
rect 171609 696337 171643 696371
rect 171643 696337 171652 696371
rect 171600 696328 171652 696337
rect 204352 696464 204404 696516
rect 579528 696464 579580 696516
rect 580448 696396 580500 696448
rect 190184 696260 190236 696312
rect 89720 696192 89772 696244
rect 580264 696192 580316 696244
rect 6828 696124 6880 696176
rect 173900 696124 173952 696176
rect 174360 696124 174412 696176
rect 412640 696124 412692 696176
rect 579436 696124 579488 696176
rect 147588 696056 147640 696108
rect 579252 696056 579304 696108
rect 124036 695988 124088 696040
rect 138480 696031 138532 696040
rect 138480 695997 138489 696031
rect 138489 695997 138523 696031
rect 138523 695997 138532 696031
rect 138480 695988 138532 695997
rect 143080 695988 143132 696040
rect 173900 695988 173952 696040
rect 174268 695988 174320 696040
rect 577780 695988 577832 696040
rect 6552 695920 6604 695972
rect 450084 695920 450136 695972
rect 5080 695852 5132 695904
rect 459652 695852 459704 695904
rect 6276 695784 6328 695836
rect 478788 695784 478840 695836
rect 3700 695648 3752 695700
rect 483388 695716 483440 695768
rect 502340 695716 502392 695768
rect 7748 695580 7800 695632
rect 4896 695512 4948 695564
rect 53288 695512 53340 695564
rect 506940 695580 506992 695632
rect 577504 695512 577556 695564
rect 7196 695444 7248 695496
rect 355508 695444 355560 695496
rect 7288 695376 7340 695428
rect 369952 695376 370004 695428
rect 3240 695308 3292 695360
rect 383844 695308 383896 695360
rect 426532 695351 426584 695360
rect 426532 695317 426541 695351
rect 426541 695317 426575 695351
rect 426575 695317 426584 695351
rect 426532 695308 426584 695317
rect 440700 695351 440752 695360
rect 440700 695317 440709 695351
rect 440709 695317 440743 695351
rect 440743 695317 440752 695351
rect 440700 695308 440752 695317
rect 469220 695351 469272 695360
rect 469220 695317 469229 695351
rect 469229 695317 469263 695351
rect 469263 695317 469272 695351
rect 469220 695308 469272 695317
rect 497556 695351 497608 695360
rect 497556 695317 497565 695351
rect 497565 695317 497599 695351
rect 497599 695317 497608 695351
rect 497556 695308 497608 695317
rect 511908 695351 511960 695360
rect 511908 695317 511917 695351
rect 511917 695317 511951 695351
rect 511951 695317 511960 695351
rect 511908 695308 511960 695317
rect 57888 695283 57940 695292
rect 57888 695249 57897 695283
rect 57897 695249 57931 695283
rect 57931 695249 57940 695283
rect 57888 695240 57940 695249
rect 67456 695283 67508 695292
rect 67456 695249 67465 695283
rect 67465 695249 67499 695283
rect 67499 695249 67508 695283
rect 67456 695240 67508 695249
rect 81348 695283 81400 695292
rect 81348 695249 81357 695283
rect 81357 695249 81391 695283
rect 81391 695249 81400 695283
rect 81348 695240 81400 695249
rect 95792 695283 95844 695292
rect 95792 695249 95801 695283
rect 95801 695249 95835 695283
rect 95835 695249 95844 695283
rect 95792 695240 95844 695249
rect 100576 695283 100628 695292
rect 100576 695249 100585 695283
rect 100585 695249 100619 695283
rect 100619 695249 100628 695283
rect 100576 695240 100628 695249
rect 109960 695283 110012 695292
rect 109960 695249 109969 695283
rect 109969 695249 110003 695283
rect 110003 695249 110012 695283
rect 109960 695240 110012 695249
rect 4068 695036 4120 695088
rect 157432 695283 157484 695292
rect 157432 695249 157441 695283
rect 157441 695249 157475 695283
rect 157475 695249 157484 695283
rect 157432 695240 157484 695249
rect 179328 695240 179380 695292
rect 185768 695240 185820 695292
rect 199936 695240 199988 695292
rect 577412 695240 577464 695292
rect 578148 695308 578200 695360
rect 578056 695104 578108 695156
rect 576032 695036 576084 695088
rect 7472 694968 7524 695020
rect 3884 694900 3936 694952
rect 3792 694764 3844 694816
rect 576676 694832 576728 694884
rect 579068 694764 579120 694816
rect 576492 694628 576544 694680
rect 578976 694560 579028 694612
rect 575296 694492 575348 694544
rect 7840 694424 7892 694476
rect 575204 694356 575256 694408
rect 575112 694288 575164 694340
rect 3608 694220 3660 694272
rect 575020 694152 575072 694204
rect 3148 693336 3200 693388
rect 578792 687148 578844 687200
rect 580908 687148 580960 687200
rect 2872 682320 2924 682372
rect 5724 682320 5776 682372
rect 575480 674772 575532 674824
rect 579804 674772 579856 674824
rect 2780 668108 2832 668160
rect 4712 668108 4764 668160
rect 3056 653556 3108 653608
rect 7196 653556 7248 653608
rect 577412 651312 577464 651364
rect 579620 651312 579672 651364
rect 575480 627852 575532 627904
rect 579804 627852 579856 627904
rect 2964 624860 3016 624912
rect 5816 624860 5868 624912
rect 2780 610988 2832 611040
rect 5448 610988 5500 611040
rect 578148 604256 578200 604308
rect 579620 604256 579672 604308
rect 3056 596028 3108 596080
rect 7288 596028 7340 596080
rect 575388 580864 575440 580916
rect 580172 580864 580224 580916
rect 2964 567468 3016 567520
rect 5908 567468 5960 567520
rect 578056 557336 578108 557388
rect 579620 557336 579672 557388
rect 577964 534012 578016 534064
rect 579712 534012 579764 534064
rect 576032 510552 576084 510604
rect 580172 510552 580224 510604
rect 3056 510348 3108 510400
rect 6000 510348 6052 510400
rect 577872 499060 577924 499112
rect 580172 499060 580224 499112
rect 576768 487092 576820 487144
rect 579988 487092 580040 487144
rect 3240 481108 3292 481160
rect 7380 481108 7432 481160
rect 577780 463632 577832 463684
rect 579620 463632 579672 463684
rect 3056 452412 3108 452464
rect 6092 452412 6144 452464
rect 3976 440240 4028 440292
rect 5356 440240 5408 440292
rect 576676 440172 576728 440224
rect 579988 440172 580040 440224
rect 3332 423920 3384 423972
rect 6828 423920 6880 423972
rect 576584 416576 576636 416628
rect 580172 416576 580224 416628
rect 3332 395700 3384 395752
rect 6736 395700 6788 395752
rect 4068 378428 4120 378480
rect 5264 378428 5316 378480
rect 3332 366188 3384 366240
rect 7472 366188 7524 366240
rect 577688 358708 577740 358760
rect 580816 358708 580868 358760
rect 576492 346332 576544 346384
rect 579988 346332 580040 346384
rect 3332 337900 3384 337952
rect 6644 337900 6696 337952
rect 2780 323892 2832 323944
rect 5172 323892 5224 323944
rect 577596 311788 577648 311840
rect 580816 311788 580868 311840
rect 575296 299412 575348 299464
rect 579620 299412 579672 299464
rect 3332 295060 3384 295112
rect 6552 295060 6604 295112
rect 2780 280032 2832 280084
rect 5080 280032 5132 280084
rect 3148 266228 3200 266280
rect 6460 266228 6512 266280
rect 576400 264800 576452 264852
rect 580172 264800 580224 264852
rect 3240 252492 3292 252544
rect 6368 252492 6420 252544
rect 575204 252492 575256 252544
rect 580172 252492 580224 252544
rect 3148 208156 3200 208208
rect 6276 208156 6328 208208
rect 575112 205504 575164 205556
rect 580172 205504 580224 205556
rect 2780 194420 2832 194472
rect 4988 194420 5040 194472
rect 575020 182112 575072 182164
rect 580172 182112 580224 182164
rect 576308 171028 576360 171080
rect 579620 171028 579672 171080
rect 1124 165656 1176 165708
rect 7932 165656 7984 165708
rect 577504 158652 577556 158704
rect 580632 158652 580684 158704
rect 2780 150832 2832 150884
rect 4896 150832 4948 150884
rect 3332 136348 3384 136400
rect 7840 136348 7892 136400
rect 3332 122068 3384 122120
rect 7748 122068 7800 122120
rect 574928 111732 574980 111784
rect 579620 111732 579672 111784
rect 3056 79840 3108 79892
rect 7656 79840 7708 79892
rect 576216 64812 576268 64864
rect 579804 64812 579856 64864
rect 2780 64540 2832 64592
rect 4804 64540 4856 64592
rect 575020 41216 575072 41268
rect 580172 41216 580224 41268
rect 3516 35776 3568 35828
rect 7564 35776 7616 35828
rect 576124 30268 576176 30320
rect 580172 30268 580224 30320
rect 575020 17824 575072 17876
rect 580172 17824 580224 17876
rect 3148 7148 3200 7200
rect 6184 7148 6236 7200
rect 484952 6808 485004 6860
rect 495348 6808 495400 6860
rect 506664 6808 506716 6860
rect 516140 6808 516192 6860
rect 519268 6808 519320 6860
rect 531044 6808 531096 6860
rect 538772 6808 538824 6860
rect 549536 6808 549588 6860
rect 560484 6808 560536 6860
rect 570144 6808 570196 6860
rect 450544 6740 450596 6792
rect 459652 6740 459704 6792
rect 494060 6740 494112 6792
rect 504732 6740 504784 6792
rect 507860 6740 507912 6792
rect 519084 6740 519136 6792
rect 520464 6740 520516 6792
rect 532240 6740 532292 6792
rect 535276 6740 535328 6792
rect 545120 6740 545172 6792
rect 546776 6740 546828 6792
rect 556160 6740 556212 6792
rect 561680 6740 561732 6792
rect 571340 6740 571392 6792
rect 458548 6672 458600 6724
rect 467932 6672 467984 6724
rect 476948 6672 477000 6724
rect 486700 6672 486752 6724
rect 492956 6672 493008 6724
rect 503628 6672 503680 6724
rect 511264 6672 511316 6724
rect 522672 6672 522724 6724
rect 527272 6672 527324 6724
rect 539324 6672 539376 6724
rect 545580 6672 545632 6724
rect 556252 6672 556304 6724
rect 558184 6672 558236 6724
rect 568212 6672 568264 6724
rect 470048 6604 470100 6656
rect 479892 6604 479944 6656
rect 486056 6604 486108 6656
rect 496544 6604 496596 6656
rect 505560 6604 505612 6656
rect 516784 6604 516836 6656
rect 526168 6604 526220 6656
rect 538128 6604 538180 6656
rect 541072 6604 541124 6656
rect 553308 6604 553360 6656
rect 557080 6604 557132 6656
rect 568396 6604 568448 6656
rect 468852 6536 468904 6588
rect 478696 6536 478748 6588
rect 479156 6536 479208 6588
rect 489368 6536 489420 6588
rect 490656 6536 490708 6588
rect 501236 6536 501288 6588
rect 504364 6536 504416 6588
rect 515588 6536 515640 6588
rect 521568 6536 521620 6588
rect 531320 6536 531372 6588
rect 543372 6536 543424 6588
rect 553400 6536 553452 6588
rect 559380 6536 559432 6588
rect 572628 6536 572680 6588
rect 119436 6468 119488 6520
rect 123024 6468 123076 6520
rect 407028 6468 407080 6520
rect 408500 6468 408552 6520
rect 466644 6468 466696 6520
rect 476304 6468 476356 6520
rect 483756 6468 483808 6520
rect 494152 6468 494204 6520
rect 495256 6468 495308 6520
rect 506020 6468 506072 6520
rect 510160 6468 510212 6520
rect 521476 6468 521528 6520
rect 524972 6468 525024 6520
rect 536748 6468 536800 6520
rect 537576 6468 537628 6520
rect 546592 6468 546644 6520
rect 550180 6468 550232 6520
rect 560392 6468 560444 6520
rect 563980 6468 564032 6520
rect 575480 6468 575532 6520
rect 88524 6400 88576 6452
rect 93308 6400 93360 6452
rect 102784 6400 102836 6452
rect 107016 6400 107068 6452
rect 120632 6400 120684 6452
rect 124220 6400 124272 6452
rect 464344 6400 464396 6452
rect 473912 6400 473964 6452
rect 475752 6400 475804 6452
rect 485688 6400 485740 6452
rect 502064 6400 502116 6452
rect 510988 6400 511040 6452
rect 512368 6400 512420 6452
rect 523868 6400 523920 6452
rect 530768 6400 530820 6452
rect 541532 6400 541584 6452
rect 544476 6400 544528 6452
rect 554872 6400 554924 6452
rect 565084 6400 565136 6452
rect 577688 6400 577740 6452
rect 151544 6332 151596 6384
rect 153936 6332 153988 6384
rect 313188 6332 313240 6384
rect 314660 6332 314712 6384
rect 340604 6332 340656 6384
rect 342720 6332 342772 6384
rect 370412 6332 370464 6384
rect 372620 6332 372672 6384
rect 379612 6332 379664 6384
rect 382372 6332 382424 6384
rect 416228 6332 416280 6384
rect 418160 6332 418212 6384
rect 442540 6332 442592 6384
rect 445484 6332 445536 6384
rect 449440 6332 449492 6384
rect 458456 6332 458508 6384
rect 463148 6332 463200 6384
rect 472716 6332 472768 6384
rect 474648 6332 474700 6384
rect 484584 6332 484636 6384
rect 489460 6332 489512 6384
rect 500132 6332 500184 6384
rect 500224 6332 500276 6384
rect 510804 6332 510856 6384
rect 513564 6332 513616 6384
rect 525064 6332 525116 6384
rect 529572 6332 529624 6384
rect 539968 6332 540020 6384
rect 542176 6332 542228 6384
rect 552020 6332 552072 6384
rect 562784 6332 562836 6384
rect 576216 6332 576268 6384
rect 93308 6264 93360 6316
rect 97816 6264 97868 6316
rect 418528 6264 418580 6316
rect 420920 6264 420972 6316
rect 465448 6264 465500 6316
rect 475108 6264 475160 6316
rect 481456 6264 481508 6316
rect 491760 6264 491812 6316
rect 496360 6264 496412 6316
rect 507216 6264 507268 6316
rect 514668 6264 514720 6316
rect 524420 6264 524472 6316
rect 528468 6264 528520 6316
rect 539416 6264 539468 6316
rect 539876 6264 539928 6316
rect 550640 6264 550692 6316
rect 554780 6264 554832 6316
rect 564440 6264 564492 6316
rect 566188 6264 566240 6316
rect 579804 6264 579856 6316
rect 161112 6196 161164 6248
rect 163136 6196 163188 6248
rect 361212 6196 361264 6248
rect 362960 6196 363012 6248
rect 415032 6196 415084 6248
rect 416964 6196 417016 6248
rect 427636 6196 427688 6248
rect 429844 6196 429896 6248
rect 433432 6196 433484 6248
rect 436100 6196 436152 6248
rect 437940 6196 437992 6248
rect 440332 6196 440384 6248
rect 448244 6196 448296 6248
rect 457260 6196 457312 6248
rect 462044 6196 462096 6248
rect 471520 6196 471572 6248
rect 473452 6196 473504 6248
rect 483480 6196 483532 6248
rect 487252 6196 487304 6248
rect 490748 6196 490800 6248
rect 497556 6196 497608 6248
rect 508412 6196 508464 6248
rect 508964 6196 509016 6248
rect 520188 6196 520240 6248
rect 524144 6196 524196 6248
rect 535368 6196 535420 6248
rect 536472 6196 536524 6248
rect 546500 6196 546552 6248
rect 551376 6196 551428 6248
rect 561772 6196 561824 6248
rect 567384 6196 567436 6248
rect 581000 6196 581052 6248
rect 5540 6128 5592 6180
rect 10784 6128 10836 6180
rect 17592 6128 17644 6180
rect 18880 6128 18932 6180
rect 86132 6128 86184 6180
rect 91008 6128 91060 6180
rect 112352 6128 112404 6180
rect 116216 6128 116268 6180
rect 270776 6128 270828 6180
rect 272892 6128 272944 6180
rect 307392 6128 307444 6180
rect 309140 6128 309192 6180
rect 322296 6128 322348 6180
rect 324320 6128 324372 6180
rect 342904 6128 342956 6180
rect 346124 6128 346176 6180
rect 434536 6128 434588 6180
rect 443000 6128 443052 6180
rect 455144 6128 455196 6180
rect 464436 6128 464488 6180
rect 467748 6128 467800 6180
rect 477500 6128 477552 6180
rect 482652 6128 482704 6180
rect 492956 6128 493008 6180
rect 498660 6128 498712 6180
rect 509608 6128 509660 6180
rect 515864 6128 515916 6180
rect 527088 6128 527140 6180
rect 534172 6128 534224 6180
rect 546408 6128 546460 6180
rect 553676 6128 553728 6180
rect 564624 6128 564676 6180
rect 568488 6128 568540 6180
rect 582196 6128 582248 6180
rect 341800 6060 341852 6112
rect 343640 6060 343692 6112
rect 350908 6060 350960 6112
rect 353300 6060 353352 6112
rect 355508 6060 355560 6112
rect 358176 6060 358228 6112
rect 360108 6060 360160 6112
rect 362224 6060 362276 6112
rect 369216 6060 369268 6112
rect 371608 6060 371660 6112
rect 388720 6060 388772 6112
rect 391112 6060 391164 6112
rect 419632 6060 419684 6112
rect 423588 6060 423640 6112
rect 436836 6060 436888 6112
rect 439228 6060 439280 6112
rect 447140 6060 447192 6112
rect 449900 6060 449952 6112
rect 454040 6060 454092 6112
rect 457536 6060 457588 6112
rect 460848 6060 460900 6112
rect 470324 6060 470376 6112
rect 478052 6060 478104 6112
rect 488172 6060 488224 6112
rect 500960 6060 501012 6112
rect 511908 6060 511960 6112
rect 522580 6060 522632 6112
rect 531504 6060 531556 6112
rect 552480 6060 552532 6112
rect 561680 6060 561732 6112
rect 18822 5958 18874 6010
rect 18886 5958 18938 6010
rect 18950 5958 19002 6010
rect 19014 5958 19066 6010
rect 19078 5958 19130 6010
rect 19142 5958 19194 6010
rect 19206 5958 19258 6010
rect 19270 5958 19322 6010
rect 19334 5958 19386 6010
rect 54822 5958 54874 6010
rect 54886 5958 54938 6010
rect 54950 5958 55002 6010
rect 55014 5958 55066 6010
rect 55078 5958 55130 6010
rect 55142 5958 55194 6010
rect 55206 5958 55258 6010
rect 55270 5958 55322 6010
rect 55334 5958 55386 6010
rect 90822 5958 90874 6010
rect 90886 5958 90938 6010
rect 90950 5958 91002 6010
rect 91014 5958 91066 6010
rect 91078 5958 91130 6010
rect 91142 5958 91194 6010
rect 91206 5958 91258 6010
rect 91270 5958 91322 6010
rect 91334 5958 91386 6010
rect 126822 5958 126874 6010
rect 126886 5958 126938 6010
rect 126950 5958 127002 6010
rect 127014 5958 127066 6010
rect 127078 5958 127130 6010
rect 127142 5958 127194 6010
rect 127206 5958 127258 6010
rect 127270 5958 127322 6010
rect 127334 5958 127386 6010
rect 162822 5958 162874 6010
rect 162886 5958 162938 6010
rect 162950 5958 163002 6010
rect 163014 5958 163066 6010
rect 163078 5958 163130 6010
rect 163142 5958 163194 6010
rect 163206 5958 163258 6010
rect 163270 5958 163322 6010
rect 163334 5958 163386 6010
rect 198822 5958 198874 6010
rect 198886 5958 198938 6010
rect 198950 5958 199002 6010
rect 199014 5958 199066 6010
rect 199078 5958 199130 6010
rect 199142 5958 199194 6010
rect 199206 5958 199258 6010
rect 199270 5958 199322 6010
rect 199334 5958 199386 6010
rect 234822 5958 234874 6010
rect 234886 5958 234938 6010
rect 234950 5958 235002 6010
rect 235014 5958 235066 6010
rect 235078 5958 235130 6010
rect 235142 5958 235194 6010
rect 235206 5958 235258 6010
rect 235270 5958 235322 6010
rect 235334 5958 235386 6010
rect 270822 5958 270874 6010
rect 270886 5958 270938 6010
rect 270950 5958 271002 6010
rect 271014 5958 271066 6010
rect 271078 5958 271130 6010
rect 271142 5958 271194 6010
rect 271206 5958 271258 6010
rect 271270 5958 271322 6010
rect 271334 5958 271386 6010
rect 306822 5958 306874 6010
rect 306886 5958 306938 6010
rect 306950 5958 307002 6010
rect 307014 5958 307066 6010
rect 307078 5958 307130 6010
rect 307142 5958 307194 6010
rect 307206 5958 307258 6010
rect 307270 5958 307322 6010
rect 307334 5958 307386 6010
rect 342822 5958 342874 6010
rect 342886 5958 342938 6010
rect 342950 5958 343002 6010
rect 343014 5958 343066 6010
rect 343078 5958 343130 6010
rect 343142 5958 343194 6010
rect 343206 5958 343258 6010
rect 343270 5958 343322 6010
rect 343334 5958 343386 6010
rect 378822 5958 378874 6010
rect 378886 5958 378938 6010
rect 378950 5958 379002 6010
rect 379014 5958 379066 6010
rect 379078 5958 379130 6010
rect 379142 5958 379194 6010
rect 379206 5958 379258 6010
rect 379270 5958 379322 6010
rect 379334 5958 379386 6010
rect 414822 5958 414874 6010
rect 414886 5958 414938 6010
rect 414950 5958 415002 6010
rect 415014 5958 415066 6010
rect 415078 5958 415130 6010
rect 415142 5958 415194 6010
rect 415206 5958 415258 6010
rect 415270 5958 415322 6010
rect 415334 5958 415386 6010
rect 450822 5958 450874 6010
rect 450886 5958 450938 6010
rect 450950 5958 451002 6010
rect 451014 5958 451066 6010
rect 451078 5958 451130 6010
rect 451142 5958 451194 6010
rect 451206 5958 451258 6010
rect 451270 5958 451322 6010
rect 451334 5958 451386 6010
rect 486822 5958 486874 6010
rect 486886 5958 486938 6010
rect 486950 5958 487002 6010
rect 487014 5958 487066 6010
rect 487078 5958 487130 6010
rect 487142 5958 487194 6010
rect 487206 5958 487258 6010
rect 487270 5958 487322 6010
rect 487334 5958 487386 6010
rect 522822 5958 522874 6010
rect 522886 5958 522938 6010
rect 522950 5958 523002 6010
rect 523014 5958 523066 6010
rect 523078 5958 523130 6010
rect 523142 5958 523194 6010
rect 523206 5958 523258 6010
rect 523270 5958 523322 6010
rect 523334 5958 523386 6010
rect 558822 5958 558874 6010
rect 558886 5958 558938 6010
rect 558950 5958 559002 6010
rect 559014 5958 559066 6010
rect 559078 5958 559130 6010
rect 559142 5958 559194 6010
rect 559206 5958 559258 6010
rect 559270 5958 559322 6010
rect 559334 5958 559386 6010
rect 331496 5856 331548 5908
rect 333980 5856 334032 5908
rect 402428 5856 402480 5908
rect 405648 5856 405700 5908
rect 410524 5856 410576 5908
rect 413744 5856 413796 5908
rect 421932 5856 421984 5908
rect 424508 5856 424560 5908
rect 431132 5856 431184 5908
rect 434168 5856 434220 5908
rect 440240 5856 440292 5908
rect 443828 5856 443880 5908
rect 480352 5856 480404 5908
rect 490564 5856 490616 5908
rect 491668 5856 491720 5908
rect 502248 5856 502300 5908
rect 516968 5856 517020 5908
rect 525800 5856 525852 5908
rect 531872 5856 531924 5908
rect 541440 5856 541492 5908
rect 555884 5856 555936 5908
rect 564532 5856 564584 5908
rect 105176 5788 105228 5840
rect 109316 5788 109368 5840
rect 283380 5788 283432 5840
rect 285956 5788 286008 5840
rect 292580 5788 292632 5840
rect 295524 5788 295576 5840
rect 306288 5788 306340 5840
rect 307944 5788 307996 5840
rect 321192 5788 321244 5840
rect 324136 5788 324188 5840
rect 324596 5788 324648 5840
rect 327172 5788 327224 5840
rect 333796 5788 333848 5840
rect 336648 5788 336700 5840
rect 339500 5788 339552 5840
rect 342260 5788 342312 5840
rect 349804 5788 349856 5840
rect 352288 5788 352340 5840
rect 353208 5788 353260 5840
rect 355508 5788 355560 5840
rect 368112 5788 368164 5840
rect 371056 5788 371108 5840
rect 373816 5788 373868 5840
rect 376668 5788 376720 5840
rect 380716 5788 380768 5840
rect 382280 5788 382332 5840
rect 383016 5788 383068 5840
rect 386144 5788 386196 5840
rect 387616 5788 387668 5840
rect 389180 5788 389232 5840
rect 392124 5788 392176 5840
rect 395344 5788 395396 5840
rect 396724 5788 396776 5840
rect 399852 5788 399904 5840
rect 401324 5788 401376 5840
rect 403900 5788 403952 5840
rect 408224 5788 408276 5840
rect 410432 5788 410484 5840
rect 420828 5788 420880 5840
rect 423312 5788 423364 5840
rect 425336 5788 425388 5840
rect 427820 5788 427872 5840
rect 441436 5788 441488 5840
rect 443460 5788 443512 5840
rect 443736 5788 443788 5840
rect 445852 5788 445904 5840
rect 445944 5788 445996 5840
rect 448612 5788 448664 5840
rect 456340 5788 456392 5840
rect 458640 5788 458692 5840
rect 12532 5720 12584 5772
rect 13820 5720 13872 5772
rect 94504 5720 94556 5772
rect 99012 5720 99064 5772
rect 107568 5720 107620 5772
rect 111616 5720 111668 5772
rect 113548 5720 113600 5772
rect 117320 5720 117372 5772
rect 118240 5720 118292 5772
rect 121920 5720 121972 5772
rect 123024 5720 123076 5772
rect 126520 5720 126572 5772
rect 143264 5720 143316 5772
rect 145932 5720 145984 5772
rect 152740 5720 152792 5772
rect 155132 5720 155184 5772
rect 277676 5720 277728 5772
rect 280068 5720 280120 5772
rect 282184 5720 282236 5772
rect 284760 5720 284812 5772
rect 291384 5720 291436 5772
rect 294328 5720 294380 5772
rect 297088 5720 297140 5772
rect 300308 5720 300360 5772
rect 302884 5720 302936 5772
rect 306196 5720 306248 5772
rect 308588 5720 308640 5772
rect 311808 5720 311860 5772
rect 317696 5720 317748 5772
rect 321468 5720 321520 5772
rect 332600 5720 332652 5772
rect 335820 5720 335872 5772
rect 338304 5720 338356 5772
rect 340880 5720 340932 5772
rect 365812 5720 365864 5772
rect 368664 5720 368716 5772
rect 399024 5720 399076 5772
rect 401600 5720 401652 5772
rect 12440 5652 12492 5704
rect 15384 5652 15436 5704
rect 18696 5652 18748 5704
rect 21088 5652 21140 5704
rect 22100 5652 22152 5704
rect 24584 5652 24636 5704
rect 29000 5652 29052 5704
rect 31392 5652 31444 5704
rect 79048 5652 79100 5704
rect 84108 5652 84160 5704
rect 96896 5652 96948 5704
rect 101312 5652 101364 5704
rect 101588 5652 101640 5704
rect 105912 5652 105964 5704
rect 109960 5652 110012 5704
rect 113916 5652 113968 5704
rect 114744 5652 114796 5704
rect 118424 5652 118476 5704
rect 125416 5652 125468 5704
rect 128728 5652 128780 5704
rect 129004 5652 129056 5704
rect 132224 5652 132276 5704
rect 132592 5652 132644 5704
rect 135628 5652 135680 5704
rect 136088 5652 136140 5704
rect 139124 5652 139176 5704
rect 139676 5652 139728 5704
rect 142528 5652 142580 5704
rect 144460 5652 144512 5704
rect 147128 5652 147180 5704
rect 148048 5652 148100 5704
rect 150532 5652 150584 5704
rect 157524 5652 157576 5704
rect 159732 5652 159784 5704
rect 171784 5652 171836 5704
rect 173440 5652 173492 5704
rect 184756 5652 184808 5704
rect 186044 5652 186096 5704
rect 248972 5652 249024 5704
rect 250352 5652 250404 5704
rect 266176 5652 266228 5704
rect 268108 5652 268160 5704
rect 276480 5652 276532 5704
rect 278872 5652 278924 5704
rect 281080 5652 281132 5704
rect 283656 5652 283708 5704
rect 286784 5652 286836 5704
rect 289544 5652 289596 5704
rect 290280 5652 290332 5704
rect 293132 5652 293184 5704
rect 295984 5652 296036 5704
rect 299112 5652 299164 5704
rect 300584 5652 300636 5704
rect 303528 5652 303580 5704
rect 311992 5652 312044 5704
rect 315764 5652 315816 5704
rect 319996 5652 320048 5704
rect 322020 5652 322072 5704
rect 328000 5652 328052 5704
rect 330116 5652 330168 5704
rect 337200 5652 337252 5704
rect 339500 5652 339552 5704
rect 345204 5652 345256 5704
rect 347780 5652 347832 5704
rect 348608 5652 348660 5704
rect 351092 5652 351144 5704
rect 354404 5652 354456 5704
rect 357256 5652 357308 5704
rect 358912 5652 358964 5704
rect 361580 5652 361632 5704
rect 363512 5652 363564 5704
rect 366548 5652 366600 5704
rect 372712 5652 372764 5704
rect 375840 5652 375892 5704
rect 376116 5652 376168 5704
rect 379428 5652 379480 5704
rect 386420 5652 386472 5704
rect 389640 5652 389692 5704
rect 395620 5652 395672 5704
rect 398748 5652 398800 5704
rect 405924 5652 405976 5704
rect 409420 5652 409472 5704
rect 413928 5652 413980 5704
rect 416688 5652 416740 5704
rect 428832 5652 428884 5704
rect 430580 5652 430632 5704
rect 444840 5652 444892 5704
rect 448060 5652 448112 5704
rect 457444 5652 457496 5704
rect 459560 5652 459612 5704
rect 471152 5652 471204 5704
rect 473360 5652 473412 5704
rect 488356 5652 488408 5704
rect 490380 5652 490432 5704
rect 13820 5584 13872 5636
rect 16580 5584 16632 5636
rect 19432 5584 19484 5636
rect 22284 5584 22336 5636
rect 28264 5584 28316 5636
rect 30288 5584 30340 5636
rect 31760 5584 31812 5636
rect 33140 5584 33192 5636
rect 34520 5584 34572 5636
rect 37188 5584 37240 5636
rect 37648 5584 37700 5636
rect 39488 5584 39540 5636
rect 44180 5584 44232 5636
rect 46296 5584 46348 5636
rect 81440 5584 81492 5636
rect 86408 5584 86460 5636
rect 87328 5584 87380 5636
rect 92112 5584 92164 5636
rect 98092 5584 98144 5636
rect 102416 5584 102468 5636
rect 103980 5584 104032 5636
rect 108120 5584 108172 5636
rect 108672 5584 108724 5636
rect 112720 5584 112772 5636
rect 115940 5584 115992 5636
rect 119620 5584 119672 5636
rect 124220 5584 124272 5636
rect 127624 5584 127676 5636
rect 127808 5584 127860 5636
rect 131028 5584 131080 5636
rect 131396 5584 131448 5636
rect 134524 5584 134576 5636
rect 134892 5584 134944 5636
rect 137928 5584 137980 5636
rect 138480 5584 138532 5636
rect 141332 5584 141384 5636
rect 142068 5584 142120 5636
rect 144828 5584 144880 5636
rect 146852 5584 146904 5636
rect 149428 5584 149480 5636
rect 150440 5584 150492 5636
rect 152832 5584 152884 5636
rect 155132 5584 155184 5636
rect 157432 5584 157484 5636
rect 158720 5584 158772 5636
rect 160836 5584 160888 5636
rect 163504 5584 163556 5636
rect 165436 5584 165488 5636
rect 165896 5584 165948 5636
rect 167736 5584 167788 5636
rect 168196 5584 168248 5636
rect 170036 5584 170088 5636
rect 170588 5584 170640 5636
rect 172336 5584 172388 5636
rect 174176 5584 174228 5636
rect 175740 5584 175792 5636
rect 176568 5584 176620 5636
rect 178040 5584 178092 5636
rect 178960 5584 179012 5636
rect 180340 5584 180392 5636
rect 181536 5584 181588 5636
rect 182640 5584 182692 5636
rect 247868 5584 247920 5636
rect 249156 5584 249208 5636
rect 251272 5584 251324 5636
rect 252652 5584 252704 5636
rect 253572 5584 253624 5636
rect 255044 5584 255096 5636
rect 255872 5584 255924 5636
rect 257436 5584 257488 5636
rect 258172 5584 258224 5636
rect 259828 5584 259880 5636
rect 260472 5584 260524 5636
rect 262220 5584 262272 5636
rect 262772 5584 262824 5636
rect 264612 5584 264664 5636
rect 265072 5584 265124 5636
rect 267004 5584 267056 5636
rect 268476 5584 268528 5636
rect 270500 5584 270552 5636
rect 273076 5584 273128 5636
rect 275284 5584 275336 5636
rect 275376 5584 275428 5636
rect 277676 5584 277728 5636
rect 279976 5584 280028 5636
rect 282460 5584 282512 5636
rect 285680 5584 285732 5636
rect 288348 5584 288400 5636
rect 289084 5584 289136 5636
rect 291936 5584 291988 5636
rect 294788 5584 294840 5636
rect 297916 5584 297968 5636
rect 299388 5584 299440 5636
rect 301044 5584 301096 5636
rect 301688 5584 301740 5636
rect 304908 5584 304960 5636
rect 305092 5584 305144 5636
rect 308588 5584 308640 5636
rect 310888 5584 310940 5636
rect 314568 5584 314620 5636
rect 315396 5584 315448 5636
rect 317696 5584 317748 5636
rect 318892 5584 318944 5636
rect 322848 5584 322900 5636
rect 325700 5584 325752 5636
rect 329748 5584 329800 5636
rect 330300 5584 330352 5636
rect 332600 5584 332652 5636
rect 334900 5584 334952 5636
rect 337292 5584 337344 5636
rect 346400 5584 346452 5636
rect 349160 5584 349212 5636
rect 352104 5584 352156 5636
rect 355600 5584 355652 5636
rect 357808 5584 357860 5636
rect 360568 5584 360620 5636
rect 364708 5584 364760 5636
rect 367468 5584 367520 5636
rect 377312 5584 377364 5636
rect 380440 5584 380492 5636
rect 384120 5584 384172 5636
rect 387340 5584 387392 5636
rect 389916 5584 389968 5636
rect 391940 5584 391992 5636
rect 393320 5584 393372 5636
rect 396540 5584 396592 5636
rect 397920 5584 397972 5636
rect 400496 5584 400548 5636
rect 403624 5584 403676 5636
rect 407028 5584 407080 5636
rect 409328 5584 409380 5636
rect 411260 5584 411312 5636
rect 412732 5584 412784 5636
rect 416504 5584 416556 5636
rect 423128 5584 423180 5636
rect 426256 5584 426308 5636
rect 432236 5584 432288 5636
rect 436008 5584 436060 5636
rect 451740 5584 451792 5636
rect 455328 5584 455380 5636
rect 518164 5584 518216 5636
rect 521568 5584 521620 5636
rect 547880 5584 547932 5636
rect 551928 5584 551980 5636
rect 15200 5516 15252 5568
rect 17684 5516 17736 5568
rect 18328 5516 18380 5568
rect 19984 5516 20036 5568
rect 20812 5516 20864 5568
rect 23388 5516 23440 5568
rect 23480 5516 23532 5568
rect 25688 5516 25740 5568
rect 26608 5516 26660 5568
rect 29184 5516 29236 5568
rect 30380 5516 30432 5568
rect 32588 5516 32640 5568
rect 36728 5516 36780 5568
rect 38292 5516 38344 5568
rect 40040 5516 40092 5568
rect 41420 5516 41472 5568
rect 42800 5516 42852 5568
rect 45192 5516 45244 5568
rect 53840 5516 53892 5568
rect 55496 5516 55548 5568
rect 62120 5516 62172 5568
rect 63500 5516 63552 5568
rect 71872 5516 71924 5568
rect 77208 5516 77260 5568
rect 80244 5516 80296 5568
rect 85212 5516 85264 5568
rect 89720 5516 89772 5568
rect 94412 5516 94464 5568
rect 95700 5516 95752 5568
rect 100116 5516 100168 5568
rect 100484 5516 100536 5568
rect 104716 5516 104768 5568
rect 106372 5516 106424 5568
rect 110420 5516 110472 5568
rect 111156 5516 111208 5568
rect 115020 5516 115072 5568
rect 117136 5516 117188 5568
rect 120724 5516 120776 5568
rect 121828 5516 121880 5568
rect 125324 5516 125376 5568
rect 126612 5516 126664 5568
rect 129924 5516 129976 5568
rect 130200 5516 130252 5568
rect 133328 5516 133380 5568
rect 133788 5516 133840 5568
rect 136824 5516 136876 5568
rect 137284 5516 137336 5568
rect 140228 5516 140280 5568
rect 140872 5516 140924 5568
rect 143632 5516 143684 5568
rect 145656 5516 145708 5568
rect 148232 5516 148284 5568
rect 149244 5516 149296 5568
rect 151636 5516 151688 5568
rect 153936 5516 153988 5568
rect 156236 5516 156288 5568
rect 156328 5516 156380 5568
rect 158536 5516 158588 5568
rect 159916 5516 159968 5568
rect 161940 5516 161992 5568
rect 162308 5516 162360 5568
rect 164240 5516 164292 5568
rect 164700 5516 164752 5568
rect 166540 5516 166592 5568
rect 167092 5516 167144 5568
rect 168840 5516 168892 5568
rect 169392 5516 169444 5568
rect 171140 5516 171192 5568
rect 172980 5516 173032 5568
rect 174544 5516 174596 5568
rect 175372 5516 175424 5568
rect 176844 5516 176896 5568
rect 177764 5516 177816 5568
rect 179144 5516 179196 5568
rect 180156 5516 180208 5568
rect 181444 5516 181496 5568
rect 182548 5516 182600 5568
rect 183744 5516 183796 5568
rect 186044 5516 186096 5568
rect 187148 5516 187200 5568
rect 187240 5516 187292 5568
rect 188344 5516 188396 5568
rect 188436 5516 188488 5568
rect 189448 5516 189500 5568
rect 189632 5516 189684 5568
rect 190644 5516 190696 5568
rect 194416 5516 194468 5568
rect 195152 5516 195204 5568
rect 196808 5516 196860 5568
rect 197452 5516 197504 5568
rect 202696 5516 202748 5568
rect 203248 5516 203300 5568
rect 232964 5516 233016 5568
rect 233700 5516 233752 5568
rect 238668 5516 238720 5568
rect 239588 5516 239640 5568
rect 239864 5516 239916 5568
rect 240784 5516 240836 5568
rect 240968 5516 241020 5568
rect 241980 5516 242032 5568
rect 242164 5516 242216 5568
rect 243176 5516 243228 5568
rect 243268 5516 243320 5568
rect 244372 5516 244424 5568
rect 245568 5516 245620 5568
rect 246672 5516 246724 5568
rect 246764 5516 246816 5568
rect 247960 5516 248012 5568
rect 250168 5516 250220 5568
rect 251456 5516 251508 5568
rect 252468 5516 252520 5568
rect 253848 5516 253900 5568
rect 254768 5516 254820 5568
rect 256240 5516 256292 5568
rect 257068 5516 257120 5568
rect 258632 5516 258684 5568
rect 259368 5516 259420 5568
rect 261024 5516 261076 5568
rect 261576 5516 261628 5568
rect 263416 5516 263468 5568
rect 263876 5516 263928 5568
rect 265808 5516 265860 5568
rect 267372 5516 267424 5568
rect 269304 5516 269356 5568
rect 269672 5516 269724 5568
rect 271696 5516 271748 5568
rect 271880 5516 271932 5568
rect 274088 5516 274140 5568
rect 274180 5516 274232 5568
rect 276480 5516 276532 5568
rect 278780 5516 278832 5568
rect 281264 5516 281316 5568
rect 284484 5516 284536 5568
rect 287152 5516 287204 5568
rect 287980 5516 288032 5568
rect 290740 5516 290792 5568
rect 293684 5516 293736 5568
rect 296628 5516 296680 5568
rect 298284 5516 298336 5568
rect 301412 5516 301464 5568
rect 303988 5516 304040 5568
rect 307484 5516 307536 5568
rect 309692 5516 309744 5568
rect 313188 5516 313240 5568
rect 314292 5516 314344 5568
rect 316500 5516 316552 5568
rect 316592 5516 316644 5568
rect 320088 5516 320140 5568
rect 323492 5516 323544 5568
rect 326528 5516 326580 5568
rect 326896 5516 326948 5568
rect 329012 5516 329064 5568
rect 329196 5516 329248 5568
rect 331312 5516 331364 5568
rect 336096 5516 336148 5568
rect 338304 5516 338356 5568
rect 344100 5516 344152 5568
rect 346860 5516 346912 5568
rect 347504 5516 347556 5568
rect 349988 5516 350040 5568
rect 356704 5516 356756 5568
rect 359372 5516 359424 5568
rect 362408 5516 362460 5568
rect 365628 5516 365680 5568
rect 367008 5516 367060 5568
rect 369768 5516 369820 5568
rect 371516 5516 371568 5568
rect 374736 5516 374788 5568
rect 375012 5516 375064 5568
rect 378048 5516 378100 5568
rect 378416 5516 378468 5568
rect 380900 5516 380952 5568
rect 381820 5516 381872 5568
rect 384948 5516 385000 5568
rect 385316 5516 385368 5568
rect 388536 5516 388588 5568
rect 391020 5516 391072 5568
rect 393596 5516 393648 5568
rect 394424 5516 394476 5568
rect 396724 5516 396776 5568
rect 400220 5516 400272 5568
rect 404084 5516 404136 5568
rect 404728 5516 404780 5568
rect 408408 5516 408460 5568
rect 411628 5516 411680 5568
rect 414664 5516 414716 5568
rect 417332 5516 417384 5568
rect 419816 5516 419868 5568
rect 424232 5516 424284 5568
rect 426440 5516 426492 5568
rect 426532 5516 426584 5568
rect 429200 5516 429252 5568
rect 429936 5516 429988 5568
rect 432696 5516 432748 5568
rect 435640 5516 435692 5568
rect 438584 5516 438636 5568
rect 439136 5516 439188 5568
rect 442080 5516 442132 5568
rect 452844 5516 452896 5568
rect 455420 5516 455472 5568
rect 459744 5516 459796 5568
rect 463608 5516 463660 5568
rect 472348 5516 472400 5568
rect 474740 5516 474792 5568
rect 503260 5516 503312 5568
rect 506296 5516 506348 5568
rect 532976 5516 533028 5568
rect 535460 5516 535512 5568
rect 549076 5516 549128 5568
rect 550732 5516 550784 5568
rect 36822 5414 36874 5466
rect 36886 5414 36938 5466
rect 36950 5414 37002 5466
rect 37014 5414 37066 5466
rect 37078 5414 37130 5466
rect 37142 5414 37194 5466
rect 37206 5414 37258 5466
rect 37270 5414 37322 5466
rect 37334 5414 37386 5466
rect 72822 5414 72874 5466
rect 72886 5414 72938 5466
rect 72950 5414 73002 5466
rect 73014 5414 73066 5466
rect 73078 5414 73130 5466
rect 73142 5414 73194 5466
rect 73206 5414 73258 5466
rect 73270 5414 73322 5466
rect 73334 5414 73386 5466
rect 108822 5414 108874 5466
rect 108886 5414 108938 5466
rect 108950 5414 109002 5466
rect 109014 5414 109066 5466
rect 109078 5414 109130 5466
rect 109142 5414 109194 5466
rect 109206 5414 109258 5466
rect 109270 5414 109322 5466
rect 109334 5414 109386 5466
rect 144822 5414 144874 5466
rect 144886 5414 144938 5466
rect 144950 5414 145002 5466
rect 145014 5414 145066 5466
rect 145078 5414 145130 5466
rect 145142 5414 145194 5466
rect 145206 5414 145258 5466
rect 145270 5414 145322 5466
rect 145334 5414 145386 5466
rect 180822 5414 180874 5466
rect 180886 5414 180938 5466
rect 180950 5414 181002 5466
rect 181014 5414 181066 5466
rect 181078 5414 181130 5466
rect 181142 5414 181194 5466
rect 181206 5414 181258 5466
rect 181270 5414 181322 5466
rect 181334 5414 181386 5466
rect 216822 5414 216874 5466
rect 216886 5414 216938 5466
rect 216950 5414 217002 5466
rect 217014 5414 217066 5466
rect 217078 5414 217130 5466
rect 217142 5414 217194 5466
rect 217206 5414 217258 5466
rect 217270 5414 217322 5466
rect 217334 5414 217386 5466
rect 252822 5414 252874 5466
rect 252886 5414 252938 5466
rect 252950 5414 253002 5466
rect 253014 5414 253066 5466
rect 253078 5414 253130 5466
rect 253142 5414 253194 5466
rect 253206 5414 253258 5466
rect 253270 5414 253322 5466
rect 253334 5414 253386 5466
rect 288822 5414 288874 5466
rect 288886 5414 288938 5466
rect 288950 5414 289002 5466
rect 289014 5414 289066 5466
rect 289078 5414 289130 5466
rect 289142 5414 289194 5466
rect 289206 5414 289258 5466
rect 289270 5414 289322 5466
rect 289334 5414 289386 5466
rect 324822 5414 324874 5466
rect 324886 5414 324938 5466
rect 324950 5414 325002 5466
rect 325014 5414 325066 5466
rect 325078 5414 325130 5466
rect 325142 5414 325194 5466
rect 325206 5414 325258 5466
rect 325270 5414 325322 5466
rect 325334 5414 325386 5466
rect 360822 5414 360874 5466
rect 360886 5414 360938 5466
rect 360950 5414 361002 5466
rect 361014 5414 361066 5466
rect 361078 5414 361130 5466
rect 361142 5414 361194 5466
rect 361206 5414 361258 5466
rect 361270 5414 361322 5466
rect 361334 5414 361386 5466
rect 396822 5414 396874 5466
rect 396886 5414 396938 5466
rect 396950 5414 397002 5466
rect 397014 5414 397066 5466
rect 397078 5414 397130 5466
rect 397142 5414 397194 5466
rect 397206 5414 397258 5466
rect 397270 5414 397322 5466
rect 397334 5414 397386 5466
rect 432822 5414 432874 5466
rect 432886 5414 432938 5466
rect 432950 5414 433002 5466
rect 433014 5414 433066 5466
rect 433078 5414 433130 5466
rect 433142 5414 433194 5466
rect 433206 5414 433258 5466
rect 433270 5414 433322 5466
rect 433334 5414 433386 5466
rect 468822 5414 468874 5466
rect 468886 5414 468938 5466
rect 468950 5414 469002 5466
rect 469014 5414 469066 5466
rect 469078 5414 469130 5466
rect 469142 5414 469194 5466
rect 469206 5414 469258 5466
rect 469270 5414 469322 5466
rect 469334 5414 469386 5466
rect 504822 5414 504874 5466
rect 504886 5414 504938 5466
rect 504950 5414 505002 5466
rect 505014 5414 505066 5466
rect 505078 5414 505130 5466
rect 505142 5414 505194 5466
rect 505206 5414 505258 5466
rect 505270 5414 505322 5466
rect 505334 5414 505386 5466
rect 540822 5414 540874 5466
rect 540886 5414 540938 5466
rect 540950 5414 541002 5466
rect 541014 5414 541066 5466
rect 541078 5414 541130 5466
rect 541142 5414 541194 5466
rect 541206 5414 541258 5466
rect 541270 5414 541322 5466
rect 541334 5414 541386 5466
rect 576822 5414 576874 5466
rect 576886 5414 576938 5466
rect 576950 5414 577002 5466
rect 577014 5414 577066 5466
rect 577078 5414 577130 5466
rect 577142 5414 577194 5466
rect 577206 5414 577258 5466
rect 577270 5414 577322 5466
rect 577334 5414 577386 5466
rect 18822 4870 18874 4922
rect 18886 4870 18938 4922
rect 18950 4870 19002 4922
rect 19014 4870 19066 4922
rect 19078 4870 19130 4922
rect 19142 4870 19194 4922
rect 19206 4870 19258 4922
rect 19270 4870 19322 4922
rect 19334 4870 19386 4922
rect 54822 4870 54874 4922
rect 54886 4870 54938 4922
rect 54950 4870 55002 4922
rect 55014 4870 55066 4922
rect 55078 4870 55130 4922
rect 55142 4870 55194 4922
rect 55206 4870 55258 4922
rect 55270 4870 55322 4922
rect 55334 4870 55386 4922
rect 90822 4870 90874 4922
rect 90886 4870 90938 4922
rect 90950 4870 91002 4922
rect 91014 4870 91066 4922
rect 91078 4870 91130 4922
rect 91142 4870 91194 4922
rect 91206 4870 91258 4922
rect 91270 4870 91322 4922
rect 91334 4870 91386 4922
rect 126822 4870 126874 4922
rect 126886 4870 126938 4922
rect 126950 4870 127002 4922
rect 127014 4870 127066 4922
rect 127078 4870 127130 4922
rect 127142 4870 127194 4922
rect 127206 4870 127258 4922
rect 127270 4870 127322 4922
rect 127334 4870 127386 4922
rect 162822 4870 162874 4922
rect 162886 4870 162938 4922
rect 162950 4870 163002 4922
rect 163014 4870 163066 4922
rect 163078 4870 163130 4922
rect 163142 4870 163194 4922
rect 163206 4870 163258 4922
rect 163270 4870 163322 4922
rect 163334 4870 163386 4922
rect 198822 4870 198874 4922
rect 198886 4870 198938 4922
rect 198950 4870 199002 4922
rect 199014 4870 199066 4922
rect 199078 4870 199130 4922
rect 199142 4870 199194 4922
rect 199206 4870 199258 4922
rect 199270 4870 199322 4922
rect 199334 4870 199386 4922
rect 234822 4870 234874 4922
rect 234886 4870 234938 4922
rect 234950 4870 235002 4922
rect 235014 4870 235066 4922
rect 235078 4870 235130 4922
rect 235142 4870 235194 4922
rect 235206 4870 235258 4922
rect 235270 4870 235322 4922
rect 235334 4870 235386 4922
rect 270822 4870 270874 4922
rect 270886 4870 270938 4922
rect 270950 4870 271002 4922
rect 271014 4870 271066 4922
rect 271078 4870 271130 4922
rect 271142 4870 271194 4922
rect 271206 4870 271258 4922
rect 271270 4870 271322 4922
rect 271334 4870 271386 4922
rect 306822 4870 306874 4922
rect 306886 4870 306938 4922
rect 306950 4870 307002 4922
rect 307014 4870 307066 4922
rect 307078 4870 307130 4922
rect 307142 4870 307194 4922
rect 307206 4870 307258 4922
rect 307270 4870 307322 4922
rect 307334 4870 307386 4922
rect 342822 4870 342874 4922
rect 342886 4870 342938 4922
rect 342950 4870 343002 4922
rect 343014 4870 343066 4922
rect 343078 4870 343130 4922
rect 343142 4870 343194 4922
rect 343206 4870 343258 4922
rect 343270 4870 343322 4922
rect 343334 4870 343386 4922
rect 378822 4870 378874 4922
rect 378886 4870 378938 4922
rect 378950 4870 379002 4922
rect 379014 4870 379066 4922
rect 379078 4870 379130 4922
rect 379142 4870 379194 4922
rect 379206 4870 379258 4922
rect 379270 4870 379322 4922
rect 379334 4870 379386 4922
rect 414822 4870 414874 4922
rect 414886 4870 414938 4922
rect 414950 4870 415002 4922
rect 415014 4870 415066 4922
rect 415078 4870 415130 4922
rect 415142 4870 415194 4922
rect 415206 4870 415258 4922
rect 415270 4870 415322 4922
rect 415334 4870 415386 4922
rect 450822 4870 450874 4922
rect 450886 4870 450938 4922
rect 450950 4870 451002 4922
rect 451014 4870 451066 4922
rect 451078 4870 451130 4922
rect 451142 4870 451194 4922
rect 451206 4870 451258 4922
rect 451270 4870 451322 4922
rect 451334 4870 451386 4922
rect 486822 4870 486874 4922
rect 486886 4870 486938 4922
rect 486950 4870 487002 4922
rect 487014 4870 487066 4922
rect 487078 4870 487130 4922
rect 487142 4870 487194 4922
rect 487206 4870 487258 4922
rect 487270 4870 487322 4922
rect 487334 4870 487386 4922
rect 522822 4870 522874 4922
rect 522886 4870 522938 4922
rect 522950 4870 523002 4922
rect 523014 4870 523066 4922
rect 523078 4870 523130 4922
rect 523142 4870 523194 4922
rect 523206 4870 523258 4922
rect 523270 4870 523322 4922
rect 523334 4870 523386 4922
rect 558822 4870 558874 4922
rect 558886 4870 558938 4922
rect 558950 4870 559002 4922
rect 559014 4870 559066 4922
rect 559078 4870 559130 4922
rect 559142 4870 559194 4922
rect 559206 4870 559258 4922
rect 559270 4870 559322 4922
rect 559334 4870 559386 4922
rect 36822 4326 36874 4378
rect 36886 4326 36938 4378
rect 36950 4326 37002 4378
rect 37014 4326 37066 4378
rect 37078 4326 37130 4378
rect 37142 4326 37194 4378
rect 37206 4326 37258 4378
rect 37270 4326 37322 4378
rect 37334 4326 37386 4378
rect 72822 4326 72874 4378
rect 72886 4326 72938 4378
rect 72950 4326 73002 4378
rect 73014 4326 73066 4378
rect 73078 4326 73130 4378
rect 73142 4326 73194 4378
rect 73206 4326 73258 4378
rect 73270 4326 73322 4378
rect 73334 4326 73386 4378
rect 108822 4326 108874 4378
rect 108886 4326 108938 4378
rect 108950 4326 109002 4378
rect 109014 4326 109066 4378
rect 109078 4326 109130 4378
rect 109142 4326 109194 4378
rect 109206 4326 109258 4378
rect 109270 4326 109322 4378
rect 109334 4326 109386 4378
rect 144822 4326 144874 4378
rect 144886 4326 144938 4378
rect 144950 4326 145002 4378
rect 145014 4326 145066 4378
rect 145078 4326 145130 4378
rect 145142 4326 145194 4378
rect 145206 4326 145258 4378
rect 145270 4326 145322 4378
rect 145334 4326 145386 4378
rect 180822 4326 180874 4378
rect 180886 4326 180938 4378
rect 180950 4326 181002 4378
rect 181014 4326 181066 4378
rect 181078 4326 181130 4378
rect 181142 4326 181194 4378
rect 181206 4326 181258 4378
rect 181270 4326 181322 4378
rect 181334 4326 181386 4378
rect 216822 4326 216874 4378
rect 216886 4326 216938 4378
rect 216950 4326 217002 4378
rect 217014 4326 217066 4378
rect 217078 4326 217130 4378
rect 217142 4326 217194 4378
rect 217206 4326 217258 4378
rect 217270 4326 217322 4378
rect 217334 4326 217386 4378
rect 252822 4326 252874 4378
rect 252886 4326 252938 4378
rect 252950 4326 253002 4378
rect 253014 4326 253066 4378
rect 253078 4326 253130 4378
rect 253142 4326 253194 4378
rect 253206 4326 253258 4378
rect 253270 4326 253322 4378
rect 253334 4326 253386 4378
rect 288822 4326 288874 4378
rect 288886 4326 288938 4378
rect 288950 4326 289002 4378
rect 289014 4326 289066 4378
rect 289078 4326 289130 4378
rect 289142 4326 289194 4378
rect 289206 4326 289258 4378
rect 289270 4326 289322 4378
rect 289334 4326 289386 4378
rect 324822 4326 324874 4378
rect 324886 4326 324938 4378
rect 324950 4326 325002 4378
rect 325014 4326 325066 4378
rect 325078 4326 325130 4378
rect 325142 4326 325194 4378
rect 325206 4326 325258 4378
rect 325270 4326 325322 4378
rect 325334 4326 325386 4378
rect 360822 4326 360874 4378
rect 360886 4326 360938 4378
rect 360950 4326 361002 4378
rect 361014 4326 361066 4378
rect 361078 4326 361130 4378
rect 361142 4326 361194 4378
rect 361206 4326 361258 4378
rect 361270 4326 361322 4378
rect 361334 4326 361386 4378
rect 396822 4326 396874 4378
rect 396886 4326 396938 4378
rect 396950 4326 397002 4378
rect 397014 4326 397066 4378
rect 397078 4326 397130 4378
rect 397142 4326 397194 4378
rect 397206 4326 397258 4378
rect 397270 4326 397322 4378
rect 397334 4326 397386 4378
rect 432822 4326 432874 4378
rect 432886 4326 432938 4378
rect 432950 4326 433002 4378
rect 433014 4326 433066 4378
rect 433078 4326 433130 4378
rect 433142 4326 433194 4378
rect 433206 4326 433258 4378
rect 433270 4326 433322 4378
rect 433334 4326 433386 4378
rect 468822 4326 468874 4378
rect 468886 4326 468938 4378
rect 468950 4326 469002 4378
rect 469014 4326 469066 4378
rect 469078 4326 469130 4378
rect 469142 4326 469194 4378
rect 469206 4326 469258 4378
rect 469270 4326 469322 4378
rect 469334 4326 469386 4378
rect 504822 4326 504874 4378
rect 504886 4326 504938 4378
rect 504950 4326 505002 4378
rect 505014 4326 505066 4378
rect 505078 4326 505130 4378
rect 505142 4326 505194 4378
rect 505206 4326 505258 4378
rect 505270 4326 505322 4378
rect 505334 4326 505386 4378
rect 540822 4326 540874 4378
rect 540886 4326 540938 4378
rect 540950 4326 541002 4378
rect 541014 4326 541066 4378
rect 541078 4326 541130 4378
rect 541142 4326 541194 4378
rect 541206 4326 541258 4378
rect 541270 4326 541322 4378
rect 541334 4326 541386 4378
rect 576822 4326 576874 4378
rect 576886 4326 576938 4378
rect 576950 4326 577002 4378
rect 577014 4326 577066 4378
rect 577078 4326 577130 4378
rect 577142 4326 577194 4378
rect 577206 4326 577258 4378
rect 577270 4326 577322 4378
rect 577334 4326 577386 4378
rect 51632 4088 51684 4140
rect 57796 4088 57848 4140
rect 70676 4088 70728 4140
rect 76104 4088 76156 4140
rect 355508 4088 355560 4140
rect 358544 4088 358596 4140
rect 366548 4088 366600 4140
rect 369216 4088 369268 4140
rect 371608 4088 371660 4140
rect 375196 4088 375248 4140
rect 375840 4088 375892 4140
rect 378692 4088 378744 4140
rect 380900 4088 380952 4140
rect 384672 4088 384724 4140
rect 391112 4088 391164 4140
rect 395436 4088 395488 4140
rect 404084 4088 404136 4140
rect 407304 4088 407356 4140
rect 408500 4088 408552 4140
rect 414480 4088 414532 4140
rect 448060 4088 448112 4140
rect 453672 4088 453724 4140
rect 539416 4088 539468 4140
rect 540520 4088 540572 4140
rect 546500 4088 546552 4140
rect 548892 4088 548944 4140
rect 568212 4088 568264 4140
rect 571432 4088 571484 4140
rect 572 4020 624 4072
rect 8576 4020 8628 4072
rect 20720 4020 20772 4072
rect 27528 4020 27580 4072
rect 31484 4020 31536 4072
rect 36728 4020 36780 4072
rect 40960 4020 41012 4072
rect 46848 4020 46900 4072
rect 50528 4020 50580 4072
rect 56508 4020 56560 4072
rect 60004 4020 60056 4072
rect 65800 4020 65852 4072
rect 69480 4020 69532 4072
rect 74908 4020 74960 4072
rect 90732 4020 90784 4072
rect 95608 4020 95660 4072
rect 99288 4020 99340 4072
rect 103612 4020 103664 4072
rect 307944 4020 307996 4072
rect 309784 4020 309836 4072
rect 324320 4020 324372 4072
rect 326436 4020 326488 4072
rect 343640 4020 343692 4072
rect 346676 4020 346728 4072
rect 352288 4020 352340 4072
rect 354956 4020 355008 4072
rect 362960 4020 363012 4072
rect 366916 4020 366968 4072
rect 371056 4020 371108 4072
rect 374000 4020 374052 4072
rect 382372 4020 382424 4072
rect 385868 4020 385920 4072
rect 393596 4020 393648 4072
rect 397828 4020 397880 4072
rect 400496 4020 400548 4072
rect 404912 4020 404964 4072
rect 409420 4020 409472 4072
rect 413284 4020 413336 4072
rect 418160 4020 418212 4072
rect 423956 4020 424008 4072
rect 429200 4020 429252 4072
rect 434628 4020 434680 4072
rect 438584 4020 438636 4072
rect 444196 4020 444248 4072
rect 457536 4020 457588 4072
rect 463240 4020 463292 4072
rect 564440 4020 564492 4072
rect 567844 4020 567896 4072
rect 570144 4020 570196 4072
rect 573824 4020 573876 4072
rect 11244 3952 11296 4004
rect 17592 3952 17644 4004
rect 55404 3952 55456 4004
rect 61200 3952 61252 4004
rect 74264 3952 74316 4004
rect 79508 3952 79560 4004
rect 314660 3952 314712 4004
rect 316960 3952 317012 4004
rect 399852 3952 399904 4004
rect 403716 3952 403768 4004
rect 571340 3952 571392 4004
rect 575020 3952 575072 4004
rect 14832 3884 14884 3936
rect 19432 3884 19484 3936
rect 25504 3884 25556 3936
rect 30380 3884 30432 3936
rect 52828 3884 52880 3936
rect 58900 3884 58952 3936
rect 63592 3884 63644 3936
rect 69204 3884 69256 3936
rect 316500 3884 316552 3936
rect 318064 3884 318116 3936
rect 335820 3884 335872 3936
rect 337108 3884 337160 3936
rect 361580 3884 361632 3936
rect 364524 3884 364576 3936
rect 442080 3884 442132 3936
rect 447784 3884 447836 3936
rect 448612 3884 448664 3936
rect 454868 3884 454920 3936
rect 490380 3884 490432 3936
rect 498936 3884 498988 3936
rect 18822 3782 18874 3834
rect 18886 3782 18938 3834
rect 18950 3782 19002 3834
rect 19014 3782 19066 3834
rect 19078 3782 19130 3834
rect 19142 3782 19194 3834
rect 19206 3782 19258 3834
rect 19270 3782 19322 3834
rect 19334 3782 19386 3834
rect 54822 3782 54874 3834
rect 54886 3782 54938 3834
rect 54950 3782 55002 3834
rect 55014 3782 55066 3834
rect 55078 3782 55130 3834
rect 55142 3782 55194 3834
rect 55206 3782 55258 3834
rect 55270 3782 55322 3834
rect 55334 3782 55386 3834
rect 90822 3782 90874 3834
rect 90886 3782 90938 3834
rect 90950 3782 91002 3834
rect 91014 3782 91066 3834
rect 91078 3782 91130 3834
rect 91142 3782 91194 3834
rect 91206 3782 91258 3834
rect 91270 3782 91322 3834
rect 91334 3782 91386 3834
rect 126822 3782 126874 3834
rect 126886 3782 126938 3834
rect 126950 3782 127002 3834
rect 127014 3782 127066 3834
rect 127078 3782 127130 3834
rect 127142 3782 127194 3834
rect 127206 3782 127258 3834
rect 127270 3782 127322 3834
rect 127334 3782 127386 3834
rect 162822 3782 162874 3834
rect 162886 3782 162938 3834
rect 162950 3782 163002 3834
rect 163014 3782 163066 3834
rect 163078 3782 163130 3834
rect 163142 3782 163194 3834
rect 163206 3782 163258 3834
rect 163270 3782 163322 3834
rect 163334 3782 163386 3834
rect 198822 3782 198874 3834
rect 198886 3782 198938 3834
rect 198950 3782 199002 3834
rect 199014 3782 199066 3834
rect 199078 3782 199130 3834
rect 199142 3782 199194 3834
rect 199206 3782 199258 3834
rect 199270 3782 199322 3834
rect 199334 3782 199386 3834
rect 234822 3782 234874 3834
rect 234886 3782 234938 3834
rect 234950 3782 235002 3834
rect 235014 3782 235066 3834
rect 235078 3782 235130 3834
rect 235142 3782 235194 3834
rect 235206 3782 235258 3834
rect 235270 3782 235322 3834
rect 235334 3782 235386 3834
rect 270822 3782 270874 3834
rect 270886 3782 270938 3834
rect 270950 3782 271002 3834
rect 271014 3782 271066 3834
rect 271078 3782 271130 3834
rect 271142 3782 271194 3834
rect 271206 3782 271258 3834
rect 271270 3782 271322 3834
rect 271334 3782 271386 3834
rect 306822 3782 306874 3834
rect 306886 3782 306938 3834
rect 306950 3782 307002 3834
rect 307014 3782 307066 3834
rect 307078 3782 307130 3834
rect 307142 3782 307194 3834
rect 307206 3782 307258 3834
rect 307270 3782 307322 3834
rect 307334 3782 307386 3834
rect 342822 3782 342874 3834
rect 342886 3782 342938 3834
rect 342950 3782 343002 3834
rect 343014 3782 343066 3834
rect 343078 3782 343130 3834
rect 343142 3782 343194 3834
rect 343206 3782 343258 3834
rect 343270 3782 343322 3834
rect 343334 3782 343386 3834
rect 378822 3782 378874 3834
rect 378886 3782 378938 3834
rect 378950 3782 379002 3834
rect 379014 3782 379066 3834
rect 379078 3782 379130 3834
rect 379142 3782 379194 3834
rect 379206 3782 379258 3834
rect 379270 3782 379322 3834
rect 379334 3782 379386 3834
rect 414822 3782 414874 3834
rect 414886 3782 414938 3834
rect 414950 3782 415002 3834
rect 415014 3782 415066 3834
rect 415078 3782 415130 3834
rect 415142 3782 415194 3834
rect 415206 3782 415258 3834
rect 415270 3782 415322 3834
rect 415334 3782 415386 3834
rect 450822 3782 450874 3834
rect 450886 3782 450938 3834
rect 450950 3782 451002 3834
rect 451014 3782 451066 3834
rect 451078 3782 451130 3834
rect 451142 3782 451194 3834
rect 451206 3782 451258 3834
rect 451270 3782 451322 3834
rect 451334 3782 451386 3834
rect 486822 3782 486874 3834
rect 486886 3782 486938 3834
rect 486950 3782 487002 3834
rect 487014 3782 487066 3834
rect 487078 3782 487130 3834
rect 487142 3782 487194 3834
rect 487206 3782 487258 3834
rect 487270 3782 487322 3834
rect 487334 3782 487386 3834
rect 522822 3782 522874 3834
rect 522886 3782 522938 3834
rect 522950 3782 523002 3834
rect 523014 3782 523066 3834
rect 523078 3782 523130 3834
rect 523142 3782 523194 3834
rect 523206 3782 523258 3834
rect 523270 3782 523322 3834
rect 523334 3782 523386 3834
rect 558822 3782 558874 3834
rect 558886 3782 558938 3834
rect 558950 3782 559002 3834
rect 559014 3782 559066 3834
rect 559078 3782 559130 3834
rect 559142 3782 559194 3834
rect 559206 3782 559258 3834
rect 559270 3782 559322 3834
rect 559334 3782 559386 3834
rect 5264 3680 5316 3732
rect 12348 3680 12400 3732
rect 44548 3680 44600 3732
rect 50896 3680 50948 3732
rect 61200 3680 61252 3732
rect 66904 3680 66956 3732
rect 353300 3680 353352 3732
rect 356152 3680 356204 3732
rect 374736 3680 374788 3732
rect 377588 3680 377640 3732
rect 384948 3680 385000 3732
rect 388260 3680 388312 3732
rect 403900 3680 403952 3732
rect 408500 3680 408552 3732
rect 420920 3680 420972 3732
rect 426348 3680 426400 3732
rect 449900 3680 449952 3732
rect 456064 3680 456116 3732
rect 553400 3680 553452 3732
rect 555976 3680 556028 3732
rect 6460 3612 6512 3664
rect 12532 3612 12584 3664
rect 16028 3612 16080 3664
rect 20812 3612 20864 3664
rect 36176 3612 36228 3664
rect 42616 3612 42668 3664
rect 43352 3612 43404 3664
rect 49608 3612 49660 3664
rect 54024 3612 54076 3664
rect 60096 3612 60148 3664
rect 401600 3612 401652 3664
rect 406108 3612 406160 3664
rect 429844 3612 429896 3664
rect 435824 3612 435876 3664
rect 440332 3612 440384 3664
rect 446588 3612 446640 3664
rect 27896 3544 27948 3596
rect 34336 3544 34388 3596
rect 34980 3544 35032 3596
rect 40040 3544 40092 3596
rect 57612 3544 57664 3596
rect 62120 3544 62172 3596
rect 67180 3544 67232 3596
rect 72332 3544 72384 3596
rect 72700 3544 72752 3596
rect 78404 3544 78456 3596
rect 82636 3544 82688 3596
rect 87512 3544 87564 3596
rect 342720 3544 342772 3596
rect 345480 3544 345532 3596
rect 347780 3544 347832 3596
rect 350264 3544 350316 3596
rect 358176 3544 358228 3596
rect 360752 3544 360804 3596
rect 362224 3544 362276 3596
rect 365720 3544 365772 3596
rect 369768 3544 369820 3596
rect 372804 3544 372856 3596
rect 379428 3544 379480 3596
rect 382372 3544 382424 3596
rect 389180 3544 389232 3596
rect 394240 3544 394292 3596
rect 396540 3544 396592 3596
rect 400220 3544 400272 3596
rect 408408 3544 408460 3596
rect 412088 3544 412140 3596
rect 416504 3544 416556 3596
rect 420368 3544 420420 3596
rect 430580 3544 430632 3596
rect 437020 3544 437072 3596
rect 516140 3544 516192 3596
rect 517888 3544 517940 3596
rect 531320 3544 531372 3596
rect 533436 3544 533488 3596
rect 545120 3544 545172 3596
rect 547696 3544 547748 3596
rect 556160 3544 556212 3596
rect 559564 3544 559616 3596
rect 4068 3476 4120 3528
rect 11980 3476 12032 3528
rect 17224 3476 17276 3528
rect 22100 3476 22152 3528
rect 24308 3476 24360 3528
rect 29000 3476 29052 3528
rect 37464 3476 37516 3528
rect 43996 3476 44048 3528
rect 46940 3476 46992 3528
rect 53196 3476 53248 3528
rect 56416 3476 56468 3528
rect 61936 3476 61988 3528
rect 62396 3476 62448 3528
rect 68100 3476 68152 3528
rect 68284 3476 68336 3528
rect 73804 3476 73856 3528
rect 76656 3476 76708 3528
rect 81808 3476 81860 3528
rect 83832 3476 83884 3528
rect 88708 3476 88760 3528
rect 92112 3476 92164 3528
rect 96712 3476 96764 3528
rect 183744 3476 183796 3528
rect 184848 3476 184900 3528
rect 190828 3476 190880 3528
rect 191748 3476 191800 3528
rect 192024 3476 192076 3528
rect 192944 3476 192996 3528
rect 193220 3476 193272 3528
rect 194048 3476 194100 3528
rect 236460 3476 236512 3528
rect 237196 3476 237248 3528
rect 237564 3476 237616 3528
rect 238392 3476 238444 3528
rect 244464 3476 244516 3528
rect 245568 3476 245620 3528
rect 301044 3476 301096 3528
rect 302608 3476 302660 3528
rect 322020 3476 322072 3528
rect 324044 3476 324096 3528
rect 324136 3476 324188 3528
rect 325424 3476 325476 3528
rect 331312 3476 331364 3528
rect 333612 3476 333664 3528
rect 338304 3476 338356 3528
rect 340696 3476 340748 3528
rect 342260 3476 342312 3528
rect 344284 3476 344336 3528
rect 349160 3476 349212 3528
rect 351368 3476 351420 3528
rect 359372 3476 359424 3528
rect 362132 3476 362184 3528
rect 367468 3476 367520 3528
rect 370412 3476 370464 3528
rect 378048 3476 378100 3528
rect 381176 3476 381228 3528
rect 382280 3476 382332 3528
rect 387064 3476 387116 3528
rect 387340 3476 387392 3528
rect 390652 3476 390704 3528
rect 391940 3476 391992 3528
rect 396632 3476 396684 3528
rect 398748 3476 398800 3528
rect 402520 3476 402572 3528
rect 410432 3476 410484 3528
rect 415676 3476 415728 3528
rect 419816 3476 419868 3528
rect 425152 3476 425204 3528
rect 426256 3476 426308 3528
rect 431132 3476 431184 3528
rect 436008 3476 436060 3528
rect 440608 3476 440660 3528
rect 459560 3476 459612 3528
rect 466828 3476 466880 3528
rect 551928 3476 551980 3528
rect 560760 3476 560812 3528
rect 7656 3408 7708 3460
rect 12440 3408 12492 3460
rect 26700 3408 26752 3460
rect 31760 3408 31812 3460
rect 33876 3408 33928 3460
rect 39856 3408 39908 3460
rect 48136 3408 48188 3460
rect 53748 3408 53800 3460
rect 58808 3408 58860 3460
rect 64604 3408 64656 3460
rect 64788 3408 64840 3460
rect 70216 3408 70268 3460
rect 77852 3408 77904 3460
rect 83004 3408 83056 3460
rect 329012 3408 329064 3460
rect 331220 3408 331272 3460
rect 333980 3408 334032 3460
rect 335912 3408 335964 3460
rect 340880 3408 340932 3460
rect 342720 3408 342772 3460
rect 360568 3408 360620 3460
rect 363328 3408 363380 3460
rect 372620 3408 372672 3460
rect 376392 3408 376444 3460
rect 380440 3408 380492 3460
rect 383568 3408 383620 3460
rect 388536 3408 388588 3460
rect 391848 3408 391900 3460
rect 396724 3408 396776 3460
rect 401324 3408 401376 3460
rect 407028 3408 407080 3460
rect 410892 3408 410944 3460
rect 411260 3408 411312 3460
rect 416872 3408 416924 3460
rect 416964 3408 417016 3460
rect 422760 3408 422812 3460
rect 427820 3408 427872 3460
rect 433524 3408 433576 3460
rect 439228 3408 439280 3460
rect 445392 3408 445444 3460
rect 445484 3408 445536 3460
rect 451464 3408 451516 3460
rect 458640 3408 458692 3460
rect 465632 3408 465684 3460
rect 473360 3408 473412 3460
rect 481088 3408 481140 3460
rect 506296 3408 506348 3460
rect 514392 3408 514444 3460
rect 521568 3408 521620 3460
rect 529848 3408 529900 3460
rect 535460 3408 535512 3460
rect 545304 3408 545356 3460
rect 546592 3408 546644 3460
rect 550088 3408 550140 3460
rect 550732 3408 550784 3460
rect 561956 3408 562008 3460
rect 568396 3408 568448 3460
rect 570236 3408 570288 3460
rect 38568 3340 38620 3392
rect 42800 3340 42852 3392
rect 332600 3340 332652 3392
rect 334716 3340 334768 3392
rect 339500 3340 339552 3392
rect 341892 3340 341944 3392
rect 389640 3340 389692 3392
rect 393044 3340 393096 3392
rect 416688 3340 416740 3392
rect 421564 3340 421616 3392
rect 436100 3340 436152 3392
rect 441804 3340 441856 3392
rect 474740 3340 474792 3392
rect 482284 3340 482336 3392
rect 541532 3340 541584 3392
rect 542912 3340 542964 3392
rect 549536 3340 549588 3392
rect 551192 3340 551244 3392
rect 556252 3340 556304 3392
rect 558368 3340 558420 3392
rect 560392 3340 560444 3392
rect 563152 3340 563204 3392
rect 36822 3238 36874 3290
rect 36886 3238 36938 3290
rect 36950 3238 37002 3290
rect 37014 3238 37066 3290
rect 37078 3238 37130 3290
rect 37142 3238 37194 3290
rect 37206 3238 37258 3290
rect 37270 3238 37322 3290
rect 37334 3238 37386 3290
rect 72822 3238 72874 3290
rect 72886 3238 72938 3290
rect 72950 3238 73002 3290
rect 73014 3238 73066 3290
rect 73078 3238 73130 3290
rect 73142 3238 73194 3290
rect 73206 3238 73258 3290
rect 73270 3238 73322 3290
rect 73334 3238 73386 3290
rect 108822 3238 108874 3290
rect 108886 3238 108938 3290
rect 108950 3238 109002 3290
rect 109014 3238 109066 3290
rect 109078 3238 109130 3290
rect 109142 3238 109194 3290
rect 109206 3238 109258 3290
rect 109270 3238 109322 3290
rect 109334 3238 109386 3290
rect 144822 3238 144874 3290
rect 144886 3238 144938 3290
rect 144950 3238 145002 3290
rect 145014 3238 145066 3290
rect 145078 3238 145130 3290
rect 145142 3238 145194 3290
rect 145206 3238 145258 3290
rect 145270 3238 145322 3290
rect 145334 3238 145386 3290
rect 180822 3238 180874 3290
rect 180886 3238 180938 3290
rect 180950 3238 181002 3290
rect 181014 3238 181066 3290
rect 181078 3238 181130 3290
rect 181142 3238 181194 3290
rect 181206 3238 181258 3290
rect 181270 3238 181322 3290
rect 181334 3238 181386 3290
rect 216822 3238 216874 3290
rect 216886 3238 216938 3290
rect 216950 3238 217002 3290
rect 217014 3238 217066 3290
rect 217078 3238 217130 3290
rect 217142 3238 217194 3290
rect 217206 3238 217258 3290
rect 217270 3238 217322 3290
rect 217334 3238 217386 3290
rect 252822 3238 252874 3290
rect 252886 3238 252938 3290
rect 252950 3238 253002 3290
rect 253014 3238 253066 3290
rect 253078 3238 253130 3290
rect 253142 3238 253194 3290
rect 253206 3238 253258 3290
rect 253270 3238 253322 3290
rect 253334 3238 253386 3290
rect 288822 3238 288874 3290
rect 288886 3238 288938 3290
rect 288950 3238 289002 3290
rect 289014 3238 289066 3290
rect 289078 3238 289130 3290
rect 289142 3238 289194 3290
rect 289206 3238 289258 3290
rect 289270 3238 289322 3290
rect 289334 3238 289386 3290
rect 324822 3238 324874 3290
rect 324886 3238 324938 3290
rect 324950 3238 325002 3290
rect 325014 3238 325066 3290
rect 325078 3238 325130 3290
rect 325142 3238 325194 3290
rect 325206 3238 325258 3290
rect 325270 3238 325322 3290
rect 325334 3238 325386 3290
rect 360822 3238 360874 3290
rect 360886 3238 360938 3290
rect 360950 3238 361002 3290
rect 361014 3238 361066 3290
rect 361078 3238 361130 3290
rect 361142 3238 361194 3290
rect 361206 3238 361258 3290
rect 361270 3238 361322 3290
rect 361334 3238 361386 3290
rect 396822 3238 396874 3290
rect 396886 3238 396938 3290
rect 396950 3238 397002 3290
rect 397014 3238 397066 3290
rect 397078 3238 397130 3290
rect 397142 3238 397194 3290
rect 397206 3238 397258 3290
rect 397270 3238 397322 3290
rect 397334 3238 397386 3290
rect 432822 3238 432874 3290
rect 432886 3238 432938 3290
rect 432950 3238 433002 3290
rect 433014 3238 433066 3290
rect 433078 3238 433130 3290
rect 433142 3238 433194 3290
rect 433206 3238 433258 3290
rect 433270 3238 433322 3290
rect 433334 3238 433386 3290
rect 468822 3238 468874 3290
rect 468886 3238 468938 3290
rect 468950 3238 469002 3290
rect 469014 3238 469066 3290
rect 469078 3238 469130 3290
rect 469142 3238 469194 3290
rect 469206 3238 469258 3290
rect 469270 3238 469322 3290
rect 469334 3238 469386 3290
rect 504822 3238 504874 3290
rect 504886 3238 504938 3290
rect 504950 3238 505002 3290
rect 505014 3238 505066 3290
rect 505078 3238 505130 3290
rect 505142 3238 505194 3290
rect 505206 3238 505258 3290
rect 505270 3238 505322 3290
rect 505334 3238 505386 3290
rect 540822 3238 540874 3290
rect 540886 3238 540938 3290
rect 540950 3238 541002 3290
rect 541014 3238 541066 3290
rect 541078 3238 541130 3290
rect 541142 3238 541194 3290
rect 541206 3238 541258 3290
rect 541270 3238 541322 3290
rect 541334 3238 541386 3290
rect 576822 3238 576874 3290
rect 576886 3238 576938 3290
rect 576950 3238 577002 3290
rect 577014 3238 577066 3290
rect 577078 3238 577130 3290
rect 577142 3238 577194 3290
rect 577206 3238 577258 3290
rect 577270 3238 577322 3290
rect 577334 3238 577386 3290
rect 23112 3136 23164 3188
rect 28264 3136 28316 3188
rect 45744 3136 45796 3188
rect 52092 3136 52144 3188
rect 65984 3136 66036 3188
rect 71504 3136 71556 3188
rect 75460 3136 75512 3188
rect 80704 3136 80756 3188
rect 309140 3136 309192 3188
rect 310980 3136 311032 3188
rect 330116 3136 330168 3188
rect 332416 3136 332468 3188
rect 349988 3136 350040 3188
rect 352564 3136 352616 3188
rect 368664 3136 368716 3188
rect 371608 3136 371660 3188
rect 376668 3136 376720 3188
rect 379980 3136 380032 3188
rect 405648 3136 405700 3188
rect 409696 3136 409748 3188
rect 423588 3136 423640 3188
rect 427544 3136 427596 3188
rect 445852 3136 445904 3188
rect 452476 3136 452528 3188
rect 463608 3136 463660 3188
rect 468668 3136 468720 3188
rect 510988 3136 511040 3188
rect 513196 3136 513248 3188
rect 524420 3136 524472 3188
rect 526260 3136 526312 3188
rect 541440 3136 541492 3188
rect 544108 3136 544160 3188
rect 550640 3136 550692 3188
rect 552388 3136 552440 3188
rect 554872 3136 554924 3188
rect 557172 3136 557224 3188
rect 561680 3136 561732 3188
rect 565544 3136 565596 3188
rect 575480 3136 575532 3188
rect 577412 3136 577464 3188
rect 577688 3136 577740 3188
rect 578608 3136 578660 3188
rect 12440 3068 12492 3120
rect 18328 3068 18380 3120
rect 32680 3068 32732 3120
rect 37648 3068 37700 3120
rect 42156 3068 42208 3120
rect 48228 3068 48280 3120
rect 346124 3068 346176 3120
rect 347872 3068 347924 3120
rect 351092 3068 351144 3120
rect 353760 3068 353812 3120
rect 426440 3068 426492 3120
rect 432328 3068 432380 3120
rect 455420 3068 455472 3120
rect 462044 3068 462096 3120
rect 490748 3068 490800 3120
rect 497740 3068 497792 3120
rect 539968 3068 540020 3120
rect 541716 3068 541768 3120
rect 552020 3068 552072 3120
rect 554780 3068 554832 3120
rect 561772 3068 561824 3120
rect 564348 3068 564400 3120
rect 564624 3068 564676 3120
rect 566740 3068 566792 3120
rect 1676 3000 1728 3052
rect 9588 3000 9640 3052
rect 19524 3000 19576 3052
rect 26148 3000 26200 3052
rect 326528 3000 326580 3052
rect 327632 3000 327684 3052
rect 365628 3000 365680 3052
rect 368020 3000 368072 3052
rect 386144 3000 386196 3052
rect 389456 3000 389508 3052
rect 413744 3000 413796 3052
rect 417976 3000 418028 3052
rect 434168 3000 434220 3052
rect 439412 3000 439464 3052
rect 455328 3000 455380 3052
rect 460848 3000 460900 3052
rect 525800 3000 525852 3052
rect 528652 3000 528704 3052
rect 531504 3000 531556 3052
rect 534540 3000 534592 3052
rect 564532 3000 564584 3052
rect 569040 3000 569092 3052
rect 8852 2932 8904 2984
rect 13820 2932 13872 2984
rect 18328 2932 18380 2984
rect 23480 2932 23532 2984
rect 84936 2932 84988 2984
rect 89812 2932 89864 2984
rect 336648 2932 336700 2984
rect 338304 2932 338356 2984
rect 424508 2932 424560 2984
rect 429936 2932 429988 2984
rect 443828 2932 443880 2984
rect 448980 2932 449032 2984
rect 2872 2864 2924 2916
rect 5540 2864 5592 2916
rect 10048 2864 10100 2916
rect 15200 2864 15252 2916
rect 21916 2864 21968 2916
rect 26608 2864 26660 2916
rect 29092 2864 29144 2916
rect 35808 2864 35860 2916
rect 327172 2864 327224 2916
rect 328828 2864 328880 2916
rect 337292 2864 337344 2916
rect 339500 2864 339552 2916
rect 357256 2864 357308 2916
rect 359740 2864 359792 2916
rect 395344 2864 395396 2916
rect 399024 2864 399076 2916
rect 423312 2864 423364 2916
rect 428740 2864 428792 2916
rect 432696 2864 432748 2916
rect 438216 2864 438268 2916
rect 443460 2864 443512 2916
rect 450176 2864 450228 2916
rect 13636 2796 13688 2848
rect 18696 2796 18748 2848
rect 30288 2796 30340 2848
rect 34520 2796 34572 2848
rect 39764 2796 39816 2848
rect 44180 2796 44232 2848
rect 49332 2796 49384 2848
rect 53840 2796 53892 2848
rect 317696 2796 317748 2848
rect 319260 2796 319312 2848
rect 346860 2796 346912 2848
rect 349068 2796 349120 2848
rect 355600 2796 355652 2848
rect 357348 2796 357400 2848
rect 414664 2796 414716 2848
rect 419172 2796 419224 2848
rect 18822 2694 18874 2746
rect 18886 2694 18938 2746
rect 18950 2694 19002 2746
rect 19014 2694 19066 2746
rect 19078 2694 19130 2746
rect 19142 2694 19194 2746
rect 19206 2694 19258 2746
rect 19270 2694 19322 2746
rect 19334 2694 19386 2746
rect 54822 2694 54874 2746
rect 54886 2694 54938 2746
rect 54950 2694 55002 2746
rect 55014 2694 55066 2746
rect 55078 2694 55130 2746
rect 55142 2694 55194 2746
rect 55206 2694 55258 2746
rect 55270 2694 55322 2746
rect 55334 2694 55386 2746
rect 90822 2694 90874 2746
rect 90886 2694 90938 2746
rect 90950 2694 91002 2746
rect 91014 2694 91066 2746
rect 91078 2694 91130 2746
rect 91142 2694 91194 2746
rect 91206 2694 91258 2746
rect 91270 2694 91322 2746
rect 91334 2694 91386 2746
rect 126822 2694 126874 2746
rect 126886 2694 126938 2746
rect 126950 2694 127002 2746
rect 127014 2694 127066 2746
rect 127078 2694 127130 2746
rect 127142 2694 127194 2746
rect 127206 2694 127258 2746
rect 127270 2694 127322 2746
rect 127334 2694 127386 2746
rect 162822 2694 162874 2746
rect 162886 2694 162938 2746
rect 162950 2694 163002 2746
rect 163014 2694 163066 2746
rect 163078 2694 163130 2746
rect 163142 2694 163194 2746
rect 163206 2694 163258 2746
rect 163270 2694 163322 2746
rect 163334 2694 163386 2746
rect 198822 2694 198874 2746
rect 198886 2694 198938 2746
rect 198950 2694 199002 2746
rect 199014 2694 199066 2746
rect 199078 2694 199130 2746
rect 199142 2694 199194 2746
rect 199206 2694 199258 2746
rect 199270 2694 199322 2746
rect 199334 2694 199386 2746
rect 234822 2694 234874 2746
rect 234886 2694 234938 2746
rect 234950 2694 235002 2746
rect 235014 2694 235066 2746
rect 235078 2694 235130 2746
rect 235142 2694 235194 2746
rect 235206 2694 235258 2746
rect 235270 2694 235322 2746
rect 235334 2694 235386 2746
rect 270822 2694 270874 2746
rect 270886 2694 270938 2746
rect 270950 2694 271002 2746
rect 271014 2694 271066 2746
rect 271078 2694 271130 2746
rect 271142 2694 271194 2746
rect 271206 2694 271258 2746
rect 271270 2694 271322 2746
rect 271334 2694 271386 2746
rect 306822 2694 306874 2746
rect 306886 2694 306938 2746
rect 306950 2694 307002 2746
rect 307014 2694 307066 2746
rect 307078 2694 307130 2746
rect 307142 2694 307194 2746
rect 307206 2694 307258 2746
rect 307270 2694 307322 2746
rect 307334 2694 307386 2746
rect 342822 2694 342874 2746
rect 342886 2694 342938 2746
rect 342950 2694 343002 2746
rect 343014 2694 343066 2746
rect 343078 2694 343130 2746
rect 343142 2694 343194 2746
rect 343206 2694 343258 2746
rect 343270 2694 343322 2746
rect 343334 2694 343386 2746
rect 378822 2694 378874 2746
rect 378886 2694 378938 2746
rect 378950 2694 379002 2746
rect 379014 2694 379066 2746
rect 379078 2694 379130 2746
rect 379142 2694 379194 2746
rect 379206 2694 379258 2746
rect 379270 2694 379322 2746
rect 379334 2694 379386 2746
rect 414822 2694 414874 2746
rect 414886 2694 414938 2746
rect 414950 2694 415002 2746
rect 415014 2694 415066 2746
rect 415078 2694 415130 2746
rect 415142 2694 415194 2746
rect 415206 2694 415258 2746
rect 415270 2694 415322 2746
rect 415334 2694 415386 2746
rect 450822 2694 450874 2746
rect 450886 2694 450938 2746
rect 450950 2694 451002 2746
rect 451014 2694 451066 2746
rect 451078 2694 451130 2746
rect 451142 2694 451194 2746
rect 451206 2694 451258 2746
rect 451270 2694 451322 2746
rect 451334 2694 451386 2746
rect 486822 2694 486874 2746
rect 486886 2694 486938 2746
rect 486950 2694 487002 2746
rect 487014 2694 487066 2746
rect 487078 2694 487130 2746
rect 487142 2694 487194 2746
rect 487206 2694 487258 2746
rect 487270 2694 487322 2746
rect 487334 2694 487386 2746
rect 522822 2694 522874 2746
rect 522886 2694 522938 2746
rect 522950 2694 523002 2746
rect 523014 2694 523066 2746
rect 523078 2694 523130 2746
rect 523142 2694 523194 2746
rect 523206 2694 523258 2746
rect 523270 2694 523322 2746
rect 523334 2694 523386 2746
rect 558822 2694 558874 2746
rect 558886 2694 558938 2746
rect 558950 2694 559002 2746
rect 559014 2694 559066 2746
rect 559078 2694 559130 2746
rect 559142 2694 559194 2746
rect 559206 2694 559258 2746
rect 559270 2694 559322 2746
rect 559334 2694 559386 2746
rect 36822 2150 36874 2202
rect 36886 2150 36938 2202
rect 36950 2150 37002 2202
rect 37014 2150 37066 2202
rect 37078 2150 37130 2202
rect 37142 2150 37194 2202
rect 37206 2150 37258 2202
rect 37270 2150 37322 2202
rect 37334 2150 37386 2202
rect 72822 2150 72874 2202
rect 72886 2150 72938 2202
rect 72950 2150 73002 2202
rect 73014 2150 73066 2202
rect 73078 2150 73130 2202
rect 73142 2150 73194 2202
rect 73206 2150 73258 2202
rect 73270 2150 73322 2202
rect 73334 2150 73386 2202
rect 108822 2150 108874 2202
rect 108886 2150 108938 2202
rect 108950 2150 109002 2202
rect 109014 2150 109066 2202
rect 109078 2150 109130 2202
rect 109142 2150 109194 2202
rect 109206 2150 109258 2202
rect 109270 2150 109322 2202
rect 109334 2150 109386 2202
rect 144822 2150 144874 2202
rect 144886 2150 144938 2202
rect 144950 2150 145002 2202
rect 145014 2150 145066 2202
rect 145078 2150 145130 2202
rect 145142 2150 145194 2202
rect 145206 2150 145258 2202
rect 145270 2150 145322 2202
rect 145334 2150 145386 2202
rect 180822 2150 180874 2202
rect 180886 2150 180938 2202
rect 180950 2150 181002 2202
rect 181014 2150 181066 2202
rect 181078 2150 181130 2202
rect 181142 2150 181194 2202
rect 181206 2150 181258 2202
rect 181270 2150 181322 2202
rect 181334 2150 181386 2202
rect 216822 2150 216874 2202
rect 216886 2150 216938 2202
rect 216950 2150 217002 2202
rect 217014 2150 217066 2202
rect 217078 2150 217130 2202
rect 217142 2150 217194 2202
rect 217206 2150 217258 2202
rect 217270 2150 217322 2202
rect 217334 2150 217386 2202
rect 252822 2150 252874 2202
rect 252886 2150 252938 2202
rect 252950 2150 253002 2202
rect 253014 2150 253066 2202
rect 253078 2150 253130 2202
rect 253142 2150 253194 2202
rect 253206 2150 253258 2202
rect 253270 2150 253322 2202
rect 253334 2150 253386 2202
rect 288822 2150 288874 2202
rect 288886 2150 288938 2202
rect 288950 2150 289002 2202
rect 289014 2150 289066 2202
rect 289078 2150 289130 2202
rect 289142 2150 289194 2202
rect 289206 2150 289258 2202
rect 289270 2150 289322 2202
rect 289334 2150 289386 2202
rect 324822 2150 324874 2202
rect 324886 2150 324938 2202
rect 324950 2150 325002 2202
rect 325014 2150 325066 2202
rect 325078 2150 325130 2202
rect 325142 2150 325194 2202
rect 325206 2150 325258 2202
rect 325270 2150 325322 2202
rect 325334 2150 325386 2202
rect 360822 2150 360874 2202
rect 360886 2150 360938 2202
rect 360950 2150 361002 2202
rect 361014 2150 361066 2202
rect 361078 2150 361130 2202
rect 361142 2150 361194 2202
rect 361206 2150 361258 2202
rect 361270 2150 361322 2202
rect 361334 2150 361386 2202
rect 396822 2150 396874 2202
rect 396886 2150 396938 2202
rect 396950 2150 397002 2202
rect 397014 2150 397066 2202
rect 397078 2150 397130 2202
rect 397142 2150 397194 2202
rect 397206 2150 397258 2202
rect 397270 2150 397322 2202
rect 397334 2150 397386 2202
rect 432822 2150 432874 2202
rect 432886 2150 432938 2202
rect 432950 2150 433002 2202
rect 433014 2150 433066 2202
rect 433078 2150 433130 2202
rect 433142 2150 433194 2202
rect 433206 2150 433258 2202
rect 433270 2150 433322 2202
rect 433334 2150 433386 2202
rect 468822 2150 468874 2202
rect 468886 2150 468938 2202
rect 468950 2150 469002 2202
rect 469014 2150 469066 2202
rect 469078 2150 469130 2202
rect 469142 2150 469194 2202
rect 469206 2150 469258 2202
rect 469270 2150 469322 2202
rect 469334 2150 469386 2202
rect 504822 2150 504874 2202
rect 504886 2150 504938 2202
rect 504950 2150 505002 2202
rect 505014 2150 505066 2202
rect 505078 2150 505130 2202
rect 505142 2150 505194 2202
rect 505206 2150 505258 2202
rect 505270 2150 505322 2202
rect 505334 2150 505386 2202
rect 540822 2150 540874 2202
rect 540886 2150 540938 2202
rect 540950 2150 541002 2202
rect 541014 2150 541066 2202
rect 541078 2150 541130 2202
rect 541142 2150 541194 2202
rect 541206 2150 541258 2202
rect 541270 2150 541322 2202
rect 541334 2150 541386 2202
rect 576822 2150 576874 2202
rect 576886 2150 576938 2202
rect 576950 2150 577002 2202
rect 577014 2150 577066 2202
rect 577078 2150 577130 2202
rect 577142 2150 577194 2202
rect 577206 2150 577258 2202
rect 577270 2150 577322 2202
rect 577334 2150 577386 2202
rect 226340 552 226392 604
rect 226524 552 226576 604
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 700369 8156 703520
rect 18822 701244 19386 701264
rect 18822 701242 18836 701244
rect 18892 701242 18916 701244
rect 18972 701242 18996 701244
rect 19052 701242 19076 701244
rect 19132 701242 19156 701244
rect 19212 701242 19236 701244
rect 19292 701242 19316 701244
rect 19372 701242 19386 701244
rect 19066 701190 19076 701242
rect 19132 701190 19142 701242
rect 18822 701188 18836 701190
rect 18892 701188 18916 701190
rect 18972 701188 18996 701190
rect 19052 701188 19076 701190
rect 19132 701188 19156 701190
rect 19212 701188 19236 701190
rect 19292 701188 19316 701190
rect 19372 701188 19386 701190
rect 18822 701168 19386 701188
rect 24320 700505 24348 703520
rect 36822 701788 37386 701808
rect 36822 701786 36836 701788
rect 36892 701786 36916 701788
rect 36972 701786 36996 701788
rect 37052 701786 37076 701788
rect 37132 701786 37156 701788
rect 37212 701786 37236 701788
rect 37292 701786 37316 701788
rect 37372 701786 37386 701788
rect 37066 701734 37076 701786
rect 37132 701734 37142 701786
rect 36822 701732 36836 701734
rect 36892 701732 36916 701734
rect 36972 701732 36996 701734
rect 37052 701732 37076 701734
rect 37132 701732 37156 701734
rect 37212 701732 37236 701734
rect 37292 701732 37316 701734
rect 37372 701732 37386 701734
rect 36822 701712 37386 701732
rect 40512 701049 40540 703520
rect 72988 701978 73016 703520
rect 72712 701950 73016 701978
rect 54822 701244 55386 701264
rect 54822 701242 54836 701244
rect 54892 701242 54916 701244
rect 54972 701242 54996 701244
rect 55052 701242 55076 701244
rect 55132 701242 55156 701244
rect 55212 701242 55236 701244
rect 55292 701242 55316 701244
rect 55372 701242 55386 701244
rect 55066 701190 55076 701242
rect 55132 701190 55142 701242
rect 54822 701188 54836 701190
rect 54892 701188 54916 701190
rect 54972 701188 54996 701190
rect 55052 701188 55076 701190
rect 55132 701188 55156 701190
rect 55212 701188 55236 701190
rect 55292 701188 55316 701190
rect 55372 701188 55386 701190
rect 54822 701168 55386 701188
rect 40498 701040 40554 701049
rect 40498 700975 40554 700984
rect 36822 700700 37386 700720
rect 36822 700698 36836 700700
rect 36892 700698 36916 700700
rect 36972 700698 36996 700700
rect 37052 700698 37076 700700
rect 37132 700698 37156 700700
rect 37212 700698 37236 700700
rect 37292 700698 37316 700700
rect 37372 700698 37386 700700
rect 37066 700646 37076 700698
rect 37132 700646 37142 700698
rect 36822 700644 36836 700646
rect 36892 700644 36916 700646
rect 36972 700644 36996 700646
rect 37052 700644 37076 700646
rect 37132 700644 37156 700646
rect 37212 700644 37236 700646
rect 37292 700644 37316 700646
rect 37372 700644 37386 700646
rect 36822 700624 37386 700644
rect 24306 700496 24362 700505
rect 24306 700431 24362 700440
rect 8114 700360 8170 700369
rect 72712 700330 72740 701950
rect 72822 701788 73386 701808
rect 72822 701786 72836 701788
rect 72892 701786 72916 701788
rect 72972 701786 72996 701788
rect 73052 701786 73076 701788
rect 73132 701786 73156 701788
rect 73212 701786 73236 701788
rect 73292 701786 73316 701788
rect 73372 701786 73386 701788
rect 73066 701734 73076 701786
rect 73132 701734 73142 701786
rect 72822 701732 72836 701734
rect 72892 701732 72916 701734
rect 72972 701732 72996 701734
rect 73052 701732 73076 701734
rect 73132 701732 73156 701734
rect 73212 701732 73236 701734
rect 73292 701732 73316 701734
rect 73372 701732 73386 701734
rect 72822 701712 73386 701732
rect 72822 700700 73386 700720
rect 72822 700698 72836 700700
rect 72892 700698 72916 700700
rect 72972 700698 72996 700700
rect 73052 700698 73076 700700
rect 73132 700698 73156 700700
rect 73212 700698 73236 700700
rect 73292 700698 73316 700700
rect 73372 700698 73386 700700
rect 73066 700646 73076 700698
rect 73132 700646 73142 700698
rect 72822 700644 72836 700646
rect 72892 700644 72916 700646
rect 72972 700644 72996 700646
rect 73052 700644 73076 700646
rect 73132 700644 73156 700646
rect 73212 700644 73236 700646
rect 73292 700644 73316 700646
rect 73372 700644 73386 700646
rect 72822 700624 73386 700644
rect 89180 700466 89208 703520
rect 90822 701244 91386 701264
rect 90822 701242 90836 701244
rect 90892 701242 90916 701244
rect 90972 701242 90996 701244
rect 91052 701242 91076 701244
rect 91132 701242 91156 701244
rect 91212 701242 91236 701244
rect 91292 701242 91316 701244
rect 91372 701242 91386 701244
rect 91066 701190 91076 701242
rect 91132 701190 91142 701242
rect 90822 701188 90836 701190
rect 90892 701188 90916 701190
rect 90972 701188 90996 701190
rect 91052 701188 91076 701190
rect 91132 701188 91156 701190
rect 91212 701188 91236 701190
rect 91292 701188 91316 701190
rect 91372 701188 91386 701190
rect 90822 701168 91386 701188
rect 105464 700806 105492 703520
rect 108822 701788 109386 701808
rect 108822 701786 108836 701788
rect 108892 701786 108916 701788
rect 108972 701786 108996 701788
rect 109052 701786 109076 701788
rect 109132 701786 109156 701788
rect 109212 701786 109236 701788
rect 109292 701786 109316 701788
rect 109372 701786 109386 701788
rect 109066 701734 109076 701786
rect 109132 701734 109142 701786
rect 108822 701732 108836 701734
rect 108892 701732 108916 701734
rect 108972 701732 108996 701734
rect 109052 701732 109076 701734
rect 109132 701732 109156 701734
rect 109212 701732 109236 701734
rect 109292 701732 109316 701734
rect 109372 701732 109386 701734
rect 108822 701712 109386 701732
rect 126822 701244 127386 701264
rect 126822 701242 126836 701244
rect 126892 701242 126916 701244
rect 126972 701242 126996 701244
rect 127052 701242 127076 701244
rect 127132 701242 127156 701244
rect 127212 701242 127236 701244
rect 127292 701242 127316 701244
rect 127372 701242 127386 701244
rect 127066 701190 127076 701242
rect 127132 701190 127142 701242
rect 126822 701188 126836 701190
rect 126892 701188 126916 701190
rect 126972 701188 126996 701190
rect 127052 701188 127076 701190
rect 127132 701188 127156 701190
rect 127212 701188 127236 701190
rect 127292 701188 127316 701190
rect 127372 701188 127386 701190
rect 126822 701168 127386 701188
rect 137848 700874 137876 703520
rect 144822 701788 145386 701808
rect 144822 701786 144836 701788
rect 144892 701786 144916 701788
rect 144972 701786 144996 701788
rect 145052 701786 145076 701788
rect 145132 701786 145156 701788
rect 145212 701786 145236 701788
rect 145292 701786 145316 701788
rect 145372 701786 145386 701788
rect 145066 701734 145076 701786
rect 145132 701734 145142 701786
rect 144822 701732 144836 701734
rect 144892 701732 144916 701734
rect 144972 701732 144996 701734
rect 145052 701732 145076 701734
rect 145132 701732 145156 701734
rect 145212 701732 145236 701734
rect 145292 701732 145316 701734
rect 145372 701732 145386 701734
rect 144822 701712 145386 701732
rect 154132 700942 154160 703520
rect 162822 701244 163386 701264
rect 162822 701242 162836 701244
rect 162892 701242 162916 701244
rect 162972 701242 162996 701244
rect 163052 701242 163076 701244
rect 163132 701242 163156 701244
rect 163212 701242 163236 701244
rect 163292 701242 163316 701244
rect 163372 701242 163386 701244
rect 163066 701190 163076 701242
rect 163132 701190 163142 701242
rect 162822 701188 162836 701190
rect 162892 701188 162916 701190
rect 162972 701188 162996 701190
rect 163052 701188 163076 701190
rect 163132 701188 163156 701190
rect 163212 701188 163236 701190
rect 163292 701188 163316 701190
rect 163372 701188 163386 701190
rect 162822 701168 163386 701188
rect 154120 700936 154172 700942
rect 154120 700878 154172 700884
rect 137836 700868 137888 700874
rect 137836 700810 137888 700816
rect 105452 700800 105504 700806
rect 105452 700742 105504 700748
rect 108822 700700 109386 700720
rect 108822 700698 108836 700700
rect 108892 700698 108916 700700
rect 108972 700698 108996 700700
rect 109052 700698 109076 700700
rect 109132 700698 109156 700700
rect 109212 700698 109236 700700
rect 109292 700698 109316 700700
rect 109372 700698 109386 700700
rect 109066 700646 109076 700698
rect 109132 700646 109142 700698
rect 108822 700644 108836 700646
rect 108892 700644 108916 700646
rect 108972 700644 108996 700646
rect 109052 700644 109076 700646
rect 109132 700644 109156 700646
rect 109212 700644 109236 700646
rect 109292 700644 109316 700646
rect 109372 700644 109386 700646
rect 108822 700624 109386 700644
rect 144822 700700 145386 700720
rect 144822 700698 144836 700700
rect 144892 700698 144916 700700
rect 144972 700698 144996 700700
rect 145052 700698 145076 700700
rect 145132 700698 145156 700700
rect 145212 700698 145236 700700
rect 145292 700698 145316 700700
rect 145372 700698 145386 700700
rect 145066 700646 145076 700698
rect 145132 700646 145142 700698
rect 144822 700644 144836 700646
rect 144892 700644 144916 700646
rect 144972 700644 144996 700646
rect 145052 700644 145076 700646
rect 145132 700644 145156 700646
rect 145212 700644 145236 700646
rect 145292 700644 145316 700646
rect 145372 700644 145386 700646
rect 144822 700624 145386 700644
rect 89168 700460 89220 700466
rect 89168 700402 89220 700408
rect 8114 700295 8170 700304
rect 72700 700324 72752 700330
rect 72700 700266 72752 700272
rect 170324 700262 170352 703520
rect 180822 701788 181386 701808
rect 180822 701786 180836 701788
rect 180892 701786 180916 701788
rect 180972 701786 180996 701788
rect 181052 701786 181076 701788
rect 181132 701786 181156 701788
rect 181212 701786 181236 701788
rect 181292 701786 181316 701788
rect 181372 701786 181386 701788
rect 181066 701734 181076 701786
rect 181132 701734 181142 701786
rect 180822 701732 180836 701734
rect 180892 701732 180916 701734
rect 180972 701732 180996 701734
rect 181052 701732 181076 701734
rect 181132 701732 181156 701734
rect 181212 701732 181236 701734
rect 181292 701732 181316 701734
rect 181372 701732 181386 701734
rect 180822 701712 181386 701732
rect 198822 701244 199386 701264
rect 198822 701242 198836 701244
rect 198892 701242 198916 701244
rect 198972 701242 198996 701244
rect 199052 701242 199076 701244
rect 199132 701242 199156 701244
rect 199212 701242 199236 701244
rect 199292 701242 199316 701244
rect 199372 701242 199386 701244
rect 199066 701190 199076 701242
rect 199132 701190 199142 701242
rect 198822 701188 198836 701190
rect 198892 701188 198916 701190
rect 198972 701188 198996 701190
rect 199052 701188 199076 701190
rect 199132 701188 199156 701190
rect 199212 701188 199236 701190
rect 199292 701188 199316 701190
rect 199372 701188 199386 701190
rect 198822 701168 199386 701188
rect 180822 700700 181386 700720
rect 180822 700698 180836 700700
rect 180892 700698 180916 700700
rect 180972 700698 180996 700700
rect 181052 700698 181076 700700
rect 181132 700698 181156 700700
rect 181212 700698 181236 700700
rect 181292 700698 181316 700700
rect 181372 700698 181386 700700
rect 181066 700646 181076 700698
rect 181132 700646 181142 700698
rect 180822 700644 180836 700646
rect 180892 700644 180916 700646
rect 180972 700644 180996 700646
rect 181052 700644 181076 700646
rect 181132 700644 181156 700646
rect 181212 700644 181236 700646
rect 181292 700644 181316 700646
rect 181372 700644 181386 700646
rect 180822 700624 181386 700644
rect 202800 700398 202828 703520
rect 216822 701788 217386 701808
rect 216822 701786 216836 701788
rect 216892 701786 216916 701788
rect 216972 701786 216996 701788
rect 217052 701786 217076 701788
rect 217132 701786 217156 701788
rect 217212 701786 217236 701788
rect 217292 701786 217316 701788
rect 217372 701786 217386 701788
rect 217066 701734 217076 701786
rect 217132 701734 217142 701786
rect 216822 701732 216836 701734
rect 216892 701732 216916 701734
rect 216972 701732 216996 701734
rect 217052 701732 217076 701734
rect 217132 701732 217156 701734
rect 217212 701732 217236 701734
rect 217292 701732 217316 701734
rect 217372 701732 217386 701734
rect 216822 701712 217386 701732
rect 216822 700700 217386 700720
rect 216822 700698 216836 700700
rect 216892 700698 216916 700700
rect 216972 700698 216996 700700
rect 217052 700698 217076 700700
rect 217132 700698 217156 700700
rect 217212 700698 217236 700700
rect 217292 700698 217316 700700
rect 217372 700698 217386 700700
rect 217066 700646 217076 700698
rect 217132 700646 217142 700698
rect 216822 700644 216836 700646
rect 216892 700644 216916 700646
rect 216972 700644 216996 700646
rect 217052 700644 217076 700646
rect 217132 700644 217156 700646
rect 217212 700644 217236 700646
rect 217292 700644 217316 700646
rect 217372 700644 217386 700646
rect 216822 700624 217386 700644
rect 202788 700392 202840 700398
rect 202788 700334 202840 700340
rect 170312 700256 170364 700262
rect 170312 700198 170364 700204
rect 18822 700156 19386 700176
rect 18822 700154 18836 700156
rect 18892 700154 18916 700156
rect 18972 700154 18996 700156
rect 19052 700154 19076 700156
rect 19132 700154 19156 700156
rect 19212 700154 19236 700156
rect 19292 700154 19316 700156
rect 19372 700154 19386 700156
rect 19066 700102 19076 700154
rect 19132 700102 19142 700154
rect 18822 700100 18836 700102
rect 18892 700100 18916 700102
rect 18972 700100 18996 700102
rect 19052 700100 19076 700102
rect 19132 700100 19156 700102
rect 19212 700100 19236 700102
rect 19292 700100 19316 700102
rect 19372 700100 19386 700102
rect 18822 700080 19386 700100
rect 54822 700156 55386 700176
rect 54822 700154 54836 700156
rect 54892 700154 54916 700156
rect 54972 700154 54996 700156
rect 55052 700154 55076 700156
rect 55132 700154 55156 700156
rect 55212 700154 55236 700156
rect 55292 700154 55316 700156
rect 55372 700154 55386 700156
rect 55066 700102 55076 700154
rect 55132 700102 55142 700154
rect 54822 700100 54836 700102
rect 54892 700100 54916 700102
rect 54972 700100 54996 700102
rect 55052 700100 55076 700102
rect 55132 700100 55156 700102
rect 55212 700100 55236 700102
rect 55292 700100 55316 700102
rect 55372 700100 55386 700102
rect 54822 700080 55386 700100
rect 90822 700156 91386 700176
rect 90822 700154 90836 700156
rect 90892 700154 90916 700156
rect 90972 700154 90996 700156
rect 91052 700154 91076 700156
rect 91132 700154 91156 700156
rect 91212 700154 91236 700156
rect 91292 700154 91316 700156
rect 91372 700154 91386 700156
rect 91066 700102 91076 700154
rect 91132 700102 91142 700154
rect 90822 700100 90836 700102
rect 90892 700100 90916 700102
rect 90972 700100 90996 700102
rect 91052 700100 91076 700102
rect 91132 700100 91156 700102
rect 91212 700100 91236 700102
rect 91292 700100 91316 700102
rect 91372 700100 91386 700102
rect 90822 700080 91386 700100
rect 126822 700156 127386 700176
rect 126822 700154 126836 700156
rect 126892 700154 126916 700156
rect 126972 700154 126996 700156
rect 127052 700154 127076 700156
rect 127132 700154 127156 700156
rect 127212 700154 127236 700156
rect 127292 700154 127316 700156
rect 127372 700154 127386 700156
rect 127066 700102 127076 700154
rect 127132 700102 127142 700154
rect 126822 700100 126836 700102
rect 126892 700100 126916 700102
rect 126972 700100 126996 700102
rect 127052 700100 127076 700102
rect 127132 700100 127156 700102
rect 127212 700100 127236 700102
rect 127292 700100 127316 700102
rect 127372 700100 127386 700102
rect 126822 700080 127386 700100
rect 162822 700156 163386 700176
rect 162822 700154 162836 700156
rect 162892 700154 162916 700156
rect 162972 700154 162996 700156
rect 163052 700154 163076 700156
rect 163132 700154 163156 700156
rect 163212 700154 163236 700156
rect 163292 700154 163316 700156
rect 163372 700154 163386 700156
rect 163066 700102 163076 700154
rect 163132 700102 163142 700154
rect 162822 700100 162836 700102
rect 162892 700100 162916 700102
rect 162972 700100 162996 700102
rect 163052 700100 163076 700102
rect 163132 700100 163156 700102
rect 163212 700100 163236 700102
rect 163292 700100 163316 700102
rect 163372 700100 163386 700102
rect 162822 700080 163386 700100
rect 198822 700156 199386 700176
rect 198822 700154 198836 700156
rect 198892 700154 198916 700156
rect 198972 700154 198996 700156
rect 199052 700154 199076 700156
rect 199132 700154 199156 700156
rect 199212 700154 199236 700156
rect 199292 700154 199316 700156
rect 199372 700154 199386 700156
rect 199066 700102 199076 700154
rect 199132 700102 199142 700154
rect 198822 700100 198836 700102
rect 198892 700100 198916 700102
rect 198972 700100 198996 700102
rect 199052 700100 199076 700102
rect 199132 700100 199156 700102
rect 199212 700100 199236 700102
rect 199292 700100 199316 700102
rect 199372 700100 199386 700102
rect 198822 700080 199386 700100
rect 218992 699922 219020 703520
rect 223304 701888 223356 701894
rect 223304 701830 223356 701836
rect 218980 699916 219032 699922
rect 218980 699858 219032 699864
rect 179328 699712 179380 699718
rect 179328 699654 179380 699660
rect 36822 699612 37386 699632
rect 36822 699610 36836 699612
rect 36892 699610 36916 699612
rect 36972 699610 36996 699612
rect 37052 699610 37076 699612
rect 37132 699610 37156 699612
rect 37212 699610 37236 699612
rect 37292 699610 37316 699612
rect 37372 699610 37386 699612
rect 37066 699558 37076 699610
rect 37132 699558 37142 699610
rect 36822 699556 36836 699558
rect 36892 699556 36916 699558
rect 36972 699556 36996 699558
rect 37052 699556 37076 699558
rect 37132 699556 37156 699558
rect 37212 699556 37236 699558
rect 37292 699556 37316 699558
rect 37372 699556 37386 699558
rect 36822 699536 37386 699556
rect 72822 699612 73386 699632
rect 72822 699610 72836 699612
rect 72892 699610 72916 699612
rect 72972 699610 72996 699612
rect 73052 699610 73076 699612
rect 73132 699610 73156 699612
rect 73212 699610 73236 699612
rect 73292 699610 73316 699612
rect 73372 699610 73386 699612
rect 73066 699558 73076 699610
rect 73132 699558 73142 699610
rect 72822 699556 72836 699558
rect 72892 699556 72916 699558
rect 72972 699556 72996 699558
rect 73052 699556 73076 699558
rect 73132 699556 73156 699558
rect 73212 699556 73236 699558
rect 73292 699556 73316 699558
rect 73372 699556 73386 699558
rect 72822 699536 73386 699556
rect 108822 699612 109386 699632
rect 108822 699610 108836 699612
rect 108892 699610 108916 699612
rect 108972 699610 108996 699612
rect 109052 699610 109076 699612
rect 109132 699610 109156 699612
rect 109212 699610 109236 699612
rect 109292 699610 109316 699612
rect 109372 699610 109386 699612
rect 109066 699558 109076 699610
rect 109132 699558 109142 699610
rect 108822 699556 108836 699558
rect 108892 699556 108916 699558
rect 108972 699556 108996 699558
rect 109052 699556 109076 699558
rect 109132 699556 109156 699558
rect 109212 699556 109236 699558
rect 109292 699556 109316 699558
rect 109372 699556 109386 699558
rect 108822 699536 109386 699556
rect 144822 699612 145386 699632
rect 144822 699610 144836 699612
rect 144892 699610 144916 699612
rect 144972 699610 144996 699612
rect 145052 699610 145076 699612
rect 145132 699610 145156 699612
rect 145212 699610 145236 699612
rect 145292 699610 145316 699612
rect 145372 699610 145386 699612
rect 145066 699558 145076 699610
rect 145132 699558 145142 699610
rect 144822 699556 144836 699558
rect 144892 699556 144916 699558
rect 144972 699556 144996 699558
rect 145052 699556 145076 699558
rect 145132 699556 145156 699558
rect 145212 699556 145236 699558
rect 145292 699556 145316 699558
rect 145372 699556 145386 699558
rect 144822 699536 145386 699556
rect 86040 699508 86092 699514
rect 86040 699450 86092 699456
rect 71780 699440 71832 699446
rect 71780 699382 71832 699388
rect 4802 699272 4858 699281
rect 4802 699207 4858 699216
rect 5172 699236 5224 699242
rect 3976 696788 4028 696794
rect 3976 696730 4028 696736
rect 3332 696652 3384 696658
rect 3332 696594 3384 696600
rect 3240 695360 3292 695366
rect 3240 695302 3292 695308
rect 3148 693388 3200 693394
rect 3148 693330 3200 693336
rect 2872 682372 2924 682378
rect 2872 682314 2924 682320
rect 2884 682281 2912 682314
rect 2870 682272 2926 682281
rect 2870 682207 2926 682216
rect 2780 668160 2832 668166
rect 2780 668102 2832 668108
rect 2792 668001 2820 668102
rect 2778 667992 2834 668001
rect 2778 667927 2834 667936
rect 3056 653608 3108 653614
rect 3054 653576 3056 653585
rect 3108 653576 3110 653585
rect 3054 653511 3110 653520
rect 2964 624912 3016 624918
rect 2962 624880 2964 624889
rect 3016 624880 3018 624889
rect 2962 624815 3018 624824
rect 2780 611040 2832 611046
rect 2780 610982 2832 610988
rect 2792 610473 2820 610982
rect 2778 610464 2834 610473
rect 2778 610399 2834 610408
rect 3056 596080 3108 596086
rect 3054 596048 3056 596057
rect 3108 596048 3110 596057
rect 3054 595983 3110 595992
rect 2964 567520 3016 567526
rect 2964 567462 3016 567468
rect 2976 567361 3004 567462
rect 2962 567352 3018 567361
rect 2962 567287 3018 567296
rect 3160 553081 3188 693330
rect 3146 553072 3202 553081
rect 3146 553007 3202 553016
rect 3252 538665 3280 695302
rect 3238 538656 3294 538665
rect 3238 538591 3294 538600
rect 3056 510400 3108 510406
rect 3056 510342 3108 510348
rect 3068 509969 3096 510342
rect 3054 509960 3110 509969
rect 3054 509895 3110 509904
rect 3240 481160 3292 481166
rect 3238 481128 3240 481137
rect 3292 481128 3294 481137
rect 3238 481063 3294 481072
rect 3056 452464 3108 452470
rect 3054 452432 3056 452441
rect 3108 452432 3110 452441
rect 3054 452367 3110 452376
rect 3344 438025 3372 696594
rect 3422 695736 3478 695745
rect 3422 695671 3478 695680
rect 3700 695700 3752 695706
rect 3330 438016 3386 438025
rect 3330 437951 3386 437960
rect 3332 423972 3384 423978
rect 3332 423914 3384 423920
rect 3344 423745 3372 423914
rect 3330 423736 3386 423745
rect 3330 423671 3386 423680
rect 3332 395752 3384 395758
rect 3332 395694 3384 395700
rect 3344 395049 3372 395694
rect 3330 395040 3386 395049
rect 3330 394975 3386 394984
rect 3332 366240 3384 366246
rect 3330 366208 3332 366217
rect 3384 366208 3386 366217
rect 3330 366143 3386 366152
rect 3332 337952 3384 337958
rect 3332 337894 3384 337900
rect 3344 337521 3372 337894
rect 3330 337512 3386 337521
rect 3330 337447 3386 337456
rect 2780 323944 2832 323950
rect 2780 323886 2832 323892
rect 2792 323105 2820 323886
rect 2778 323096 2834 323105
rect 2778 323031 2834 323040
rect 3332 295112 3384 295118
rect 3332 295054 3384 295060
rect 3344 294409 3372 295054
rect 3330 294400 3386 294409
rect 3330 294335 3386 294344
rect 2778 280120 2834 280129
rect 2778 280055 2780 280064
rect 2832 280055 2834 280064
rect 2780 280026 2832 280032
rect 3148 266280 3200 266286
rect 3148 266222 3200 266228
rect 3160 265713 3188 266222
rect 3146 265704 3202 265713
rect 3146 265639 3202 265648
rect 3240 252544 3292 252550
rect 3240 252486 3292 252492
rect 3252 251297 3280 252486
rect 3238 251288 3294 251297
rect 3238 251223 3294 251232
rect 3148 208208 3200 208214
rect 3146 208176 3148 208185
rect 3200 208176 3202 208185
rect 3146 208111 3202 208120
rect 2780 194472 2832 194478
rect 2780 194414 2832 194420
rect 2792 193905 2820 194414
rect 2778 193896 2834 193905
rect 2778 193831 2834 193840
rect 1124 165708 1176 165714
rect 1124 165650 1176 165656
rect 1136 165073 1164 165650
rect 1122 165064 1178 165073
rect 1122 164999 1178 165008
rect 2780 150884 2832 150890
rect 2780 150826 2832 150832
rect 2792 150793 2820 150826
rect 2778 150784 2834 150793
rect 2778 150719 2834 150728
rect 3332 136400 3384 136406
rect 3330 136368 3332 136377
rect 3384 136368 3386 136377
rect 3330 136303 3386 136312
rect 3332 122120 3384 122126
rect 3330 122088 3332 122097
rect 3384 122088 3386 122097
rect 3330 122023 3386 122032
rect 3056 79892 3108 79898
rect 3056 79834 3108 79840
rect 3068 78985 3096 79834
rect 3054 78976 3110 78985
rect 3054 78911 3110 78920
rect 2780 64592 2832 64598
rect 2778 64560 2780 64569
rect 2832 64560 2834 64569
rect 2778 64495 2834 64504
rect 3436 21457 3464 695671
rect 3700 695642 3752 695648
rect 3608 694272 3660 694278
rect 3608 694214 3660 694220
rect 3514 693968 3570 693977
rect 3514 693903 3570 693912
rect 3528 50153 3556 693903
rect 3620 93265 3648 694214
rect 3712 179489 3740 695642
rect 3884 694952 3936 694958
rect 3884 694894 3936 694900
rect 3792 694816 3844 694822
rect 3792 694758 3844 694764
rect 3804 222601 3832 694758
rect 3896 308825 3924 694894
rect 3988 495553 4016 696730
rect 4712 696720 4764 696726
rect 4712 696662 4764 696668
rect 4068 695088 4120 695094
rect 4068 695030 4120 695036
rect 3974 495544 4030 495553
rect 3974 495479 4030 495488
rect 3976 440292 4028 440298
rect 3976 440234 4028 440240
rect 3882 308816 3938 308825
rect 3882 308751 3938 308760
rect 3790 222592 3846 222601
rect 3790 222527 3846 222536
rect 3698 179480 3754 179489
rect 3698 179415 3754 179424
rect 3988 107681 4016 440234
rect 4080 380633 4108 695030
rect 4724 668166 4752 696662
rect 4712 668160 4764 668166
rect 4712 668102 4764 668108
rect 4066 380624 4122 380633
rect 4066 380559 4122 380568
rect 4068 378480 4120 378486
rect 4068 378422 4120 378428
rect 4080 237017 4108 378422
rect 4066 237008 4122 237017
rect 4066 236943 4122 236952
rect 3974 107672 4030 107681
rect 3974 107607 4030 107616
rect 3606 93256 3662 93265
rect 3606 93191 3662 93200
rect 4816 64598 4844 699207
rect 5172 699178 5224 699184
rect 4988 698692 5040 698698
rect 4988 698634 5040 698640
rect 4896 695564 4948 695570
rect 4896 695506 4948 695512
rect 4908 150890 4936 695506
rect 5000 194478 5028 698634
rect 5080 695904 5132 695910
rect 5080 695846 5132 695852
rect 5092 280090 5120 695846
rect 5184 323950 5212 699178
rect 18822 699068 19386 699088
rect 18822 699066 18836 699068
rect 18892 699066 18916 699068
rect 18972 699066 18996 699068
rect 19052 699066 19076 699068
rect 19132 699066 19156 699068
rect 19212 699066 19236 699068
rect 19292 699066 19316 699068
rect 19372 699066 19386 699068
rect 19066 699014 19076 699066
rect 19132 699014 19142 699066
rect 18822 699012 18836 699014
rect 18892 699012 18916 699014
rect 18972 699012 18996 699014
rect 19052 699012 19076 699014
rect 19132 699012 19156 699014
rect 19212 699012 19236 699014
rect 19292 699012 19316 699014
rect 19372 699012 19386 699014
rect 18822 698992 19386 699012
rect 54822 699068 55386 699088
rect 54822 699066 54836 699068
rect 54892 699066 54916 699068
rect 54972 699066 54996 699068
rect 55052 699066 55076 699068
rect 55132 699066 55156 699068
rect 55212 699066 55236 699068
rect 55292 699066 55316 699068
rect 55372 699066 55386 699068
rect 55066 699014 55076 699066
rect 55132 699014 55142 699066
rect 54822 699012 54836 699014
rect 54892 699012 54916 699014
rect 54972 699012 54996 699014
rect 55052 699012 55076 699014
rect 55132 699012 55156 699014
rect 55212 699012 55236 699014
rect 55292 699012 55316 699014
rect 55372 699012 55386 699014
rect 54822 698992 55386 699012
rect 48136 698964 48188 698970
rect 48136 698906 48188 698912
rect 43442 698864 43498 698873
rect 5264 698828 5316 698834
rect 43442 698799 43498 698808
rect 5264 698770 5316 698776
rect 5276 378486 5304 698770
rect 33968 698760 34020 698766
rect 5354 698728 5410 698737
rect 33968 698702 34020 698708
rect 5354 698663 5410 698672
rect 5368 440298 5396 698663
rect 29182 698320 29238 698329
rect 5724 698284 5776 698290
rect 29182 698255 29238 698264
rect 5724 698226 5776 698232
rect 5448 696584 5500 696590
rect 5448 696526 5500 696532
rect 5460 611046 5488 696526
rect 5736 682378 5764 698226
rect 5816 698216 5868 698222
rect 5816 698158 5868 698164
rect 5724 682372 5776 682378
rect 5724 682314 5776 682320
rect 5828 624918 5856 698158
rect 5908 698080 5960 698086
rect 5908 698022 5960 698028
rect 5816 624912 5868 624918
rect 5816 624854 5868 624860
rect 5448 611040 5500 611046
rect 5448 610982 5500 610988
rect 5920 567526 5948 698022
rect 6000 697876 6052 697882
rect 6000 697818 6052 697824
rect 5908 567520 5960 567526
rect 5908 567462 5960 567468
rect 6012 510406 6040 697818
rect 7380 697808 7432 697814
rect 7380 697750 7432 697756
rect 6092 697672 6144 697678
rect 6092 697614 6144 697620
rect 6000 510400 6052 510406
rect 6000 510342 6052 510348
rect 6104 452470 6132 697614
rect 6736 697536 6788 697542
rect 6736 697478 6788 697484
rect 6644 697400 6696 697406
rect 6644 697342 6696 697348
rect 6460 697332 6512 697338
rect 6460 697274 6512 697280
rect 6368 697264 6420 697270
rect 6368 697206 6420 697212
rect 6182 697096 6238 697105
rect 6182 697031 6238 697040
rect 6092 452464 6144 452470
rect 6092 452406 6144 452412
rect 5356 440292 5408 440298
rect 5356 440234 5408 440240
rect 5264 378480 5316 378486
rect 5264 378422 5316 378428
rect 5172 323944 5224 323950
rect 5172 323886 5224 323892
rect 5080 280084 5132 280090
rect 5080 280026 5132 280032
rect 4988 194472 5040 194478
rect 4988 194414 5040 194420
rect 4896 150884 4948 150890
rect 4896 150826 4948 150832
rect 4804 64592 4856 64598
rect 4804 64534 4856 64540
rect 3514 50144 3570 50153
rect 3514 50079 3570 50088
rect 3514 35864 3570 35873
rect 3514 35799 3516 35808
rect 3568 35799 3570 35808
rect 3516 35770 3568 35776
rect 3422 21448 3478 21457
rect 3422 21383 3478 21392
rect 6196 7206 6224 697031
rect 6276 695836 6328 695842
rect 6276 695778 6328 695784
rect 6288 208214 6316 695778
rect 6380 252550 6408 697206
rect 6472 266286 6500 697274
rect 6552 695972 6604 695978
rect 6552 695914 6604 695920
rect 6564 295118 6592 695914
rect 6656 337958 6684 697342
rect 6748 395758 6776 697478
rect 6828 696176 6880 696182
rect 6828 696118 6880 696124
rect 6840 423978 6868 696118
rect 7196 695496 7248 695502
rect 7196 695438 7248 695444
rect 7208 653614 7236 695438
rect 7288 695428 7340 695434
rect 7288 695370 7340 695376
rect 7196 653608 7248 653614
rect 7196 653550 7248 653556
rect 7300 596086 7328 695370
rect 7288 596080 7340 596086
rect 7288 596022 7340 596028
rect 7392 481166 7420 697750
rect 7932 697196 7984 697202
rect 7932 697138 7984 697144
rect 7564 697128 7616 697134
rect 7564 697070 7616 697076
rect 7472 695020 7524 695026
rect 7472 694962 7524 694968
rect 7380 481160 7432 481166
rect 7380 481102 7432 481108
rect 6828 423972 6880 423978
rect 6828 423914 6880 423920
rect 6736 395752 6788 395758
rect 6736 395694 6788 395700
rect 7484 366246 7512 694962
rect 7472 366240 7524 366246
rect 7472 366182 7524 366188
rect 6644 337952 6696 337958
rect 6644 337894 6696 337900
rect 6552 295112 6604 295118
rect 6552 295054 6604 295060
rect 6460 266280 6512 266286
rect 6460 266222 6512 266228
rect 6368 252544 6420 252550
rect 6368 252486 6420 252492
rect 6276 208208 6328 208214
rect 6276 208150 6328 208156
rect 7576 35834 7604 697070
rect 7748 695632 7800 695638
rect 7748 695574 7800 695580
rect 7654 693696 7710 693705
rect 7654 693631 7710 693640
rect 7668 79898 7696 693631
rect 7760 122126 7788 695574
rect 7840 694476 7892 694482
rect 7840 694418 7892 694424
rect 7852 136406 7880 694418
rect 7944 165714 7972 697138
rect 24492 696992 24544 696998
rect 10322 696960 10378 696969
rect 24492 696934 24544 696940
rect 10322 696895 10378 696904
rect 10336 695980 10364 696895
rect 24504 695980 24532 696934
rect 29196 695980 29224 698255
rect 33980 695980 34008 698702
rect 36822 698524 37386 698544
rect 36822 698522 36836 698524
rect 36892 698522 36916 698524
rect 36972 698522 36996 698524
rect 37052 698522 37076 698524
rect 37132 698522 37156 698524
rect 37212 698522 37236 698524
rect 37292 698522 37316 698524
rect 37372 698522 37386 698524
rect 37066 698470 37076 698522
rect 37132 698470 37142 698522
rect 36822 698468 36836 698470
rect 36892 698468 36916 698470
rect 36972 698468 36996 698470
rect 37052 698468 37076 698470
rect 37132 698468 37156 698470
rect 37212 698468 37236 698470
rect 37292 698468 37316 698470
rect 37372 698468 37386 698470
rect 36822 698448 37386 698468
rect 38660 697060 38712 697066
rect 38660 697002 38712 697008
rect 38672 695980 38700 697002
rect 43456 695980 43484 698799
rect 48148 695980 48176 698906
rect 62304 698352 62356 698358
rect 62304 698294 62356 698300
rect 62316 695980 62344 698294
rect 71792 695980 71820 699382
rect 72822 698524 73386 698544
rect 72822 698522 72836 698524
rect 72892 698522 72916 698524
rect 72972 698522 72996 698524
rect 73052 698522 73076 698524
rect 73132 698522 73156 698524
rect 73212 698522 73236 698524
rect 73292 698522 73316 698524
rect 73372 698522 73386 698524
rect 73066 698470 73076 698522
rect 73132 698470 73142 698522
rect 72822 698468 72836 698470
rect 72892 698468 72916 698470
rect 72972 698468 72996 698470
rect 73052 698468 73076 698470
rect 73132 698468 73156 698470
rect 73212 698468 73236 698470
rect 73292 698468 73316 698470
rect 73372 698468 73386 698470
rect 72822 698448 73386 698468
rect 76564 698420 76616 698426
rect 76564 698362 76616 698368
rect 76576 695980 76604 698362
rect 86052 695980 86080 699450
rect 114376 699372 114428 699378
rect 114376 699314 114428 699320
rect 90822 699068 91386 699088
rect 90822 699066 90836 699068
rect 90892 699066 90916 699068
rect 90972 699066 90996 699068
rect 91052 699066 91076 699068
rect 91132 699066 91156 699068
rect 91212 699066 91236 699068
rect 91292 699066 91316 699068
rect 91372 699066 91386 699068
rect 91066 699014 91076 699066
rect 91132 699014 91142 699066
rect 90822 699012 90836 699014
rect 90892 699012 90916 699014
rect 90972 699012 90996 699014
rect 91052 699012 91076 699014
rect 91132 699012 91156 699014
rect 91212 699012 91236 699014
rect 91292 699012 91316 699014
rect 91372 699012 91386 699014
rect 90822 698992 91386 699012
rect 89720 698760 89772 698766
rect 89720 698702 89772 698708
rect 104992 698760 105044 698766
rect 104992 698702 105044 698708
rect 89732 696250 89760 698702
rect 90732 698624 90784 698630
rect 90732 698566 90784 698572
rect 89720 696244 89772 696250
rect 89720 696186 89772 696192
rect 90744 695980 90772 698566
rect 105004 695980 105032 698702
rect 108822 698524 109386 698544
rect 108822 698522 108836 698524
rect 108892 698522 108916 698524
rect 108972 698522 108996 698524
rect 109052 698522 109076 698524
rect 109132 698522 109156 698524
rect 109212 698522 109236 698524
rect 109292 698522 109316 698524
rect 109372 698522 109386 698524
rect 109066 698470 109076 698522
rect 109132 698470 109142 698522
rect 108822 698468 108836 698470
rect 108892 698468 108916 698470
rect 108972 698468 108996 698470
rect 109052 698468 109076 698470
rect 109132 698468 109156 698470
rect 109212 698468 109236 698470
rect 109292 698468 109316 698470
rect 109372 698468 109386 698470
rect 108822 698448 109386 698468
rect 114388 695980 114416 699314
rect 161756 699304 161808 699310
rect 161756 699246 161808 699252
rect 133328 699168 133380 699174
rect 133328 699110 133380 699116
rect 126822 699068 127386 699088
rect 126822 699066 126836 699068
rect 126892 699066 126916 699068
rect 126972 699066 126996 699068
rect 127052 699066 127076 699068
rect 127132 699066 127156 699068
rect 127212 699066 127236 699068
rect 127292 699066 127316 699068
rect 127372 699066 127386 699068
rect 127066 699014 127076 699066
rect 127132 699014 127142 699066
rect 126822 699012 126836 699014
rect 126892 699012 126916 699014
rect 126972 699012 126996 699014
rect 127052 699012 127076 699014
rect 127132 699012 127156 699014
rect 127212 699012 127236 699014
rect 127292 699012 127316 699014
rect 127372 699012 127386 699014
rect 126822 698992 127386 699012
rect 119712 698964 119764 698970
rect 119712 698906 119764 698912
rect 128636 698964 128688 698970
rect 128636 698906 128688 698912
rect 119160 698896 119212 698902
rect 119160 698838 119212 698844
rect 119172 695980 119200 698838
rect 119724 696454 119752 698906
rect 119712 696448 119764 696454
rect 119712 696390 119764 696396
rect 124036 696040 124088 696046
rect 123878 695988 124036 695994
rect 123878 695982 124088 695988
rect 123878 695966 124076 695982
rect 128648 695980 128676 698906
rect 133340 695980 133368 699110
rect 144822 698524 145386 698544
rect 144822 698522 144836 698524
rect 144892 698522 144916 698524
rect 144972 698522 144996 698524
rect 145052 698522 145076 698524
rect 145132 698522 145156 698524
rect 145212 698522 145236 698524
rect 145292 698522 145316 698524
rect 145372 698522 145386 698524
rect 145066 698470 145076 698522
rect 145132 698470 145142 698522
rect 144822 698468 144836 698470
rect 144892 698468 144916 698470
rect 144972 698468 144996 698470
rect 145052 698468 145076 698470
rect 145132 698468 145156 698470
rect 145212 698468 145236 698470
rect 145292 698468 145316 698470
rect 145372 698468 145386 698470
rect 144822 698448 145386 698468
rect 152280 697468 152332 697474
rect 152280 697410 152332 697416
rect 147588 696108 147640 696114
rect 147588 696050 147640 696056
rect 138480 696040 138532 696046
rect 138138 695988 138480 695994
rect 143080 696040 143132 696046
rect 138138 695982 138532 695988
rect 142830 695988 143080 695994
rect 142830 695982 143132 695988
rect 138138 695966 138520 695982
rect 142830 695966 143120 695982
rect 147600 695980 147628 696050
rect 152292 695980 152320 697410
rect 161768 695980 161796 699246
rect 162822 699068 163386 699088
rect 162822 699066 162836 699068
rect 162892 699066 162916 699068
rect 162972 699066 162996 699068
rect 163052 699066 163076 699068
rect 163132 699066 163156 699068
rect 163212 699066 163236 699068
rect 163292 699066 163316 699068
rect 163372 699066 163386 699068
rect 163066 699014 163076 699066
rect 163132 699014 163142 699066
rect 162822 699012 162836 699014
rect 162892 699012 162916 699014
rect 162972 699012 162996 699014
rect 163052 699012 163076 699014
rect 163132 699012 163156 699014
rect 163212 699012 163236 699014
rect 163292 699012 163316 699014
rect 163372 699012 163386 699014
rect 162822 698992 163386 699012
rect 166448 697604 166500 697610
rect 166448 697546 166500 697552
rect 166460 695980 166488 697546
rect 171600 696380 171652 696386
rect 171600 696322 171652 696328
rect 171612 695994 171640 696322
rect 173912 696238 174400 696266
rect 173912 696182 173940 696238
rect 174372 696182 174400 696238
rect 173900 696176 173952 696182
rect 173900 696118 173952 696124
rect 174360 696176 174412 696182
rect 174360 696118 174412 696124
rect 173900 696040 173952 696046
rect 171258 695966 171640 695994
rect 173898 696008 173900 696017
rect 174268 696040 174320 696046
rect 173952 696008 173954 696017
rect 173898 695943 173954 695952
rect 174266 696008 174268 696017
rect 174320 696008 174322 696017
rect 174266 695943 174322 695952
rect 19982 695600 20038 695609
rect 19734 695558 19982 695586
rect 52946 695570 53328 695586
rect 52946 695564 53340 695570
rect 52946 695558 53288 695564
rect 19982 695535 20038 695544
rect 53288 695506 53340 695512
rect 15290 695328 15346 695337
rect 15042 695286 15290 695314
rect 176198 695328 176254 695337
rect 57638 695298 57928 695314
rect 67114 695298 67496 695314
rect 81282 695298 81388 695314
rect 95542 695298 95832 695314
rect 100234 695298 100616 695314
rect 109710 695298 110000 695314
rect 156998 695298 157472 695314
rect 57638 695292 57940 695298
rect 57638 695286 57888 695292
rect 15290 695263 15346 695272
rect 67114 695292 67508 695298
rect 67114 695286 67456 695292
rect 57888 695234 57940 695240
rect 81282 695292 81400 695298
rect 81282 695286 81348 695292
rect 67456 695234 67508 695240
rect 95542 695292 95844 695298
rect 95542 695286 95792 695292
rect 81348 695234 81400 695240
rect 100234 695292 100628 695298
rect 100234 695286 100576 695292
rect 95792 695234 95844 695240
rect 109710 695292 110012 695298
rect 109710 695286 109960 695292
rect 100576 695234 100628 695240
rect 156998 695292 157484 695298
rect 156998 695286 157432 695292
rect 109960 695234 110012 695240
rect 175950 695286 176198 695314
rect 179340 695298 179368 699654
rect 180822 699612 181386 699632
rect 180822 699610 180836 699612
rect 180892 699610 180916 699612
rect 180972 699610 180996 699612
rect 181052 699610 181076 699612
rect 181132 699610 181156 699612
rect 181212 699610 181236 699612
rect 181292 699610 181316 699612
rect 181372 699610 181386 699612
rect 181066 699558 181076 699610
rect 181132 699558 181142 699610
rect 180822 699556 180836 699558
rect 180892 699556 180916 699558
rect 180972 699556 180996 699558
rect 181052 699556 181076 699558
rect 181132 699556 181156 699558
rect 181212 699556 181236 699558
rect 181292 699556 181316 699558
rect 181372 699556 181386 699558
rect 180822 699536 181386 699556
rect 216822 699612 217386 699632
rect 216822 699610 216836 699612
rect 216892 699610 216916 699612
rect 216972 699610 216996 699612
rect 217052 699610 217076 699612
rect 217132 699610 217156 699612
rect 217212 699610 217236 699612
rect 217292 699610 217316 699612
rect 217372 699610 217386 699612
rect 217066 699558 217076 699610
rect 217132 699558 217142 699610
rect 216822 699556 216836 699558
rect 216892 699556 216916 699558
rect 216972 699556 216996 699558
rect 217052 699556 217076 699558
rect 217132 699556 217156 699558
rect 217212 699556 217236 699558
rect 217292 699556 217316 699558
rect 217372 699556 217386 699558
rect 216822 699536 217386 699556
rect 190458 699408 190514 699417
rect 190458 699343 190514 699352
rect 200026 699408 200082 699417
rect 200026 699343 200082 699352
rect 190472 699174 190500 699343
rect 200040 699174 200068 699343
rect 180800 699168 180852 699174
rect 180798 699136 180800 699145
rect 190368 699168 190420 699174
rect 180852 699136 180854 699145
rect 180798 699071 180854 699080
rect 190366 699136 190368 699145
rect 190460 699168 190512 699174
rect 190420 699136 190422 699145
rect 190460 699110 190512 699116
rect 200028 699168 200080 699174
rect 209780 699168 209832 699174
rect 200028 699110 200080 699116
rect 209778 699136 209780 699145
rect 219348 699168 219400 699174
rect 209832 699136 209834 699145
rect 190366 699071 190422 699080
rect 198822 699068 199386 699088
rect 209778 699071 209834 699080
rect 219346 699136 219348 699145
rect 219400 699136 219402 699145
rect 219346 699071 219402 699080
rect 198822 699066 198836 699068
rect 198892 699066 198916 699068
rect 198972 699066 198996 699068
rect 199052 699066 199076 699068
rect 199132 699066 199156 699068
rect 199212 699066 199236 699068
rect 199292 699066 199316 699068
rect 199372 699066 199386 699068
rect 199066 699014 199076 699066
rect 199132 699014 199142 699066
rect 198822 699012 198836 699014
rect 198892 699012 198916 699014
rect 198972 699012 198996 699014
rect 199052 699012 199076 699014
rect 199132 699012 199156 699014
rect 199212 699012 199236 699014
rect 199292 699012 199316 699014
rect 199372 699012 199386 699014
rect 198822 698992 199386 699012
rect 180822 698524 181386 698544
rect 180822 698522 180836 698524
rect 180892 698522 180916 698524
rect 180972 698522 180996 698524
rect 181052 698522 181076 698524
rect 181132 698522 181156 698524
rect 181212 698522 181236 698524
rect 181292 698522 181316 698524
rect 181372 698522 181386 698524
rect 181066 698470 181076 698522
rect 181132 698470 181142 698522
rect 180822 698468 180836 698470
rect 180892 698468 180916 698470
rect 180972 698468 180996 698470
rect 181052 698468 181076 698470
rect 181132 698468 181156 698470
rect 181212 698468 181236 698470
rect 181292 698468 181316 698470
rect 181372 698468 181386 698470
rect 180822 698448 181386 698468
rect 216822 698524 217386 698544
rect 216822 698522 216836 698524
rect 216892 698522 216916 698524
rect 216972 698522 216996 698524
rect 217052 698522 217076 698524
rect 217132 698522 217156 698524
rect 217212 698522 217236 698524
rect 217292 698522 217316 698524
rect 217372 698522 217386 698524
rect 217066 698470 217076 698522
rect 217132 698470 217142 698522
rect 216822 698468 216836 698470
rect 216892 698468 216916 698470
rect 216972 698468 216996 698470
rect 217052 698468 217076 698470
rect 217132 698468 217156 698470
rect 217212 698468 217236 698470
rect 217292 698468 217316 698470
rect 217372 698468 217386 698470
rect 216822 698448 217386 698468
rect 209044 698148 209096 698154
rect 209044 698090 209096 698096
rect 194876 697944 194928 697950
rect 194876 697886 194928 697892
rect 180708 697740 180760 697746
rect 180708 697682 180760 697688
rect 180720 695980 180748 697682
rect 190184 696312 190236 696318
rect 190184 696254 190236 696260
rect 190196 695980 190224 696254
rect 194888 695980 194916 697886
rect 204352 696516 204404 696522
rect 204352 696458 204404 696464
rect 204364 695980 204392 696458
rect 209056 695980 209084 698090
rect 213828 698080 213880 698086
rect 213828 698022 213880 698028
rect 213840 695980 213868 698022
rect 218520 696652 218572 696658
rect 218520 696594 218572 696600
rect 218532 695980 218560 696594
rect 223316 695980 223344 701830
rect 235184 701690 235212 703520
rect 251640 702024 251692 702030
rect 251640 701966 251692 701972
rect 237472 701956 237524 701962
rect 237472 701898 237524 701904
rect 235172 701684 235224 701690
rect 235172 701626 235224 701632
rect 234822 701244 235386 701264
rect 234822 701242 234836 701244
rect 234892 701242 234916 701244
rect 234972 701242 234996 701244
rect 235052 701242 235076 701244
rect 235132 701242 235156 701244
rect 235212 701242 235236 701244
rect 235292 701242 235316 701244
rect 235372 701242 235386 701244
rect 235066 701190 235076 701242
rect 235132 701190 235142 701242
rect 234822 701188 234836 701190
rect 234892 701188 234916 701190
rect 234972 701188 234996 701190
rect 235052 701188 235076 701190
rect 235132 701188 235156 701190
rect 235212 701188 235236 701190
rect 235292 701188 235316 701190
rect 235372 701188 235386 701190
rect 234822 701168 235386 701188
rect 227994 700904 228050 700913
rect 227994 700839 228050 700848
rect 228008 695980 228036 700839
rect 234822 700156 235386 700176
rect 234822 700154 234836 700156
rect 234892 700154 234916 700156
rect 234972 700154 234996 700156
rect 235052 700154 235076 700156
rect 235132 700154 235156 700156
rect 235212 700154 235236 700156
rect 235292 700154 235316 700156
rect 235372 700154 235386 700156
rect 235066 700102 235076 700154
rect 235132 700102 235142 700154
rect 234822 700100 234836 700102
rect 234892 700100 234916 700102
rect 234972 700100 234996 700102
rect 235052 700100 235076 700102
rect 235132 700100 235156 700102
rect 235212 700100 235236 700102
rect 235292 700100 235316 700102
rect 235372 700100 235386 700102
rect 234822 700080 235386 700100
rect 229098 699408 229154 699417
rect 229098 699343 229154 699352
rect 229112 699174 229140 699343
rect 234712 699236 234764 699242
rect 234712 699178 234764 699184
rect 229100 699168 229152 699174
rect 229100 699110 229152 699116
rect 234724 698873 234752 699178
rect 234822 699068 235386 699088
rect 234822 699066 234836 699068
rect 234892 699066 234916 699068
rect 234972 699066 234996 699068
rect 235052 699066 235076 699068
rect 235132 699066 235156 699068
rect 235212 699066 235236 699068
rect 235292 699066 235316 699068
rect 235372 699066 235386 699068
rect 235066 699014 235076 699066
rect 235132 699014 235142 699066
rect 234822 699012 234836 699014
rect 234892 699012 234916 699014
rect 234972 699012 234996 699014
rect 235052 699012 235076 699014
rect 235132 699012 235156 699014
rect 235212 699012 235236 699014
rect 235292 699012 235316 699014
rect 235372 699012 235386 699014
rect 234822 698992 235386 699012
rect 233054 698864 233110 698873
rect 233054 698799 233110 698808
rect 234710 698864 234766 698873
rect 234710 698799 234766 698808
rect 233068 695994 233096 698799
rect 232806 695966 233096 695994
rect 237484 695980 237512 701898
rect 242256 700596 242308 700602
rect 242256 700538 242308 700544
rect 241520 699780 241572 699786
rect 241520 699722 241572 699728
rect 241532 699689 241560 699722
rect 241518 699680 241574 699689
rect 241518 699615 241574 699624
rect 242268 695980 242296 700538
rect 246948 700528 247000 700534
rect 246948 700470 247000 700476
rect 244186 700088 244242 700097
rect 244186 700023 244242 700032
rect 244200 699990 244228 700023
rect 244188 699984 244240 699990
rect 244188 699926 244240 699932
rect 244186 699408 244242 699417
rect 244186 699343 244242 699352
rect 244200 699174 244228 699343
rect 244096 699168 244148 699174
rect 244096 699110 244148 699116
rect 244188 699168 244240 699174
rect 244188 699110 244240 699116
rect 244108 699009 244136 699110
rect 244094 699000 244150 699009
rect 244094 698935 244150 698944
rect 246960 695980 246988 700470
rect 251086 700088 251142 700097
rect 251086 700023 251142 700032
rect 251100 699990 251128 700023
rect 251088 699984 251140 699990
rect 251088 699926 251140 699932
rect 251088 699780 251140 699786
rect 251088 699722 251140 699728
rect 251100 699689 251128 699722
rect 251086 699680 251142 699689
rect 251086 699615 251142 699624
rect 251652 695980 251680 701966
rect 252822 701788 253386 701808
rect 252822 701786 252836 701788
rect 252892 701786 252916 701788
rect 252972 701786 252996 701788
rect 253052 701786 253076 701788
rect 253132 701786 253156 701788
rect 253212 701786 253236 701788
rect 253292 701786 253316 701788
rect 253372 701786 253386 701788
rect 253066 701734 253076 701786
rect 253132 701734 253142 701786
rect 252822 701732 252836 701734
rect 252892 701732 252916 701734
rect 252972 701732 252996 701734
rect 253052 701732 253076 701734
rect 253132 701732 253156 701734
rect 253212 701732 253236 701734
rect 253292 701732 253316 701734
rect 253372 701732 253386 701734
rect 252822 701712 253386 701732
rect 256424 701004 256476 701010
rect 256424 700946 256476 700952
rect 252822 700700 253386 700720
rect 252822 700698 252836 700700
rect 252892 700698 252916 700700
rect 252972 700698 252996 700700
rect 253052 700698 253076 700700
rect 253132 700698 253156 700700
rect 253212 700698 253236 700700
rect 253292 700698 253316 700700
rect 253372 700698 253386 700700
rect 253066 700646 253076 700698
rect 253132 700646 253142 700698
rect 252822 700644 252836 700646
rect 252892 700644 252916 700646
rect 252972 700644 252996 700646
rect 253052 700644 253076 700646
rect 253132 700644 253156 700646
rect 253212 700644 253236 700646
rect 253292 700644 253316 700646
rect 253372 700644 253386 700646
rect 252822 700624 253386 700644
rect 253848 699984 253900 699990
rect 253848 699926 253900 699932
rect 252822 699612 253386 699632
rect 252822 699610 252836 699612
rect 252892 699610 252916 699612
rect 252972 699610 252996 699612
rect 253052 699610 253076 699612
rect 253132 699610 253156 699612
rect 253212 699610 253236 699612
rect 253292 699610 253316 699612
rect 253372 699610 253386 699612
rect 253066 699558 253076 699610
rect 253132 699558 253142 699610
rect 252822 699556 252836 699558
rect 252892 699556 252916 699558
rect 252972 699556 252996 699558
rect 253052 699556 253076 699558
rect 253132 699556 253156 699558
rect 253212 699556 253236 699558
rect 253292 699556 253316 699558
rect 253372 699556 253386 699558
rect 252822 699536 253386 699556
rect 253860 699242 253888 699926
rect 253848 699236 253900 699242
rect 253848 699178 253900 699184
rect 253664 699168 253716 699174
rect 253662 699136 253664 699145
rect 253716 699136 253718 699145
rect 253662 699071 253718 699080
rect 253846 699000 253902 699009
rect 253846 698935 253902 698944
rect 253860 698902 253888 698935
rect 253756 698896 253808 698902
rect 253754 698864 253756 698873
rect 253848 698896 253900 698902
rect 253808 698864 253810 698873
rect 253848 698838 253900 698844
rect 253754 698799 253810 698808
rect 252822 698524 253386 698544
rect 252822 698522 252836 698524
rect 252892 698522 252916 698524
rect 252972 698522 252996 698524
rect 253052 698522 253076 698524
rect 253132 698522 253156 698524
rect 253212 698522 253236 698524
rect 253292 698522 253316 698524
rect 253372 698522 253386 698524
rect 253066 698470 253076 698522
rect 253132 698470 253142 698522
rect 252822 698468 252836 698470
rect 252892 698468 252916 698470
rect 252972 698468 252996 698470
rect 253052 698468 253076 698470
rect 253132 698468 253156 698470
rect 253212 698468 253236 698470
rect 253292 698468 253316 698470
rect 253372 698468 253386 698470
rect 252822 698448 253386 698468
rect 256436 695980 256464 700946
rect 267660 700058 267688 703520
rect 270822 701244 271386 701264
rect 270822 701242 270836 701244
rect 270892 701242 270916 701244
rect 270972 701242 270996 701244
rect 271052 701242 271076 701244
rect 271132 701242 271156 701244
rect 271212 701242 271236 701244
rect 271292 701242 271316 701244
rect 271372 701242 271386 701244
rect 271066 701190 271076 701242
rect 271132 701190 271142 701242
rect 270822 701188 270836 701190
rect 270892 701188 270916 701190
rect 270972 701188 270996 701190
rect 271052 701188 271076 701190
rect 271132 701188 271156 701190
rect 271212 701188 271236 701190
rect 271292 701188 271316 701190
rect 271372 701188 271386 701190
rect 270822 701168 271386 701188
rect 270822 700156 271386 700176
rect 270822 700154 270836 700156
rect 270892 700154 270916 700156
rect 270972 700154 270996 700156
rect 271052 700154 271076 700156
rect 271132 700154 271156 700156
rect 271212 700154 271236 700156
rect 271292 700154 271316 700156
rect 271372 700154 271386 700156
rect 271066 700102 271076 700154
rect 271132 700102 271142 700154
rect 270822 700100 270836 700102
rect 270892 700100 270916 700102
rect 270972 700100 270996 700102
rect 271052 700100 271076 700102
rect 271132 700100 271156 700102
rect 271212 700100 271236 700102
rect 271292 700100 271316 700102
rect 271372 700100 271386 700102
rect 270822 700080 271386 700100
rect 280066 700088 280122 700097
rect 267648 700052 267700 700058
rect 283852 700058 283880 703520
rect 288822 701788 289386 701808
rect 288822 701786 288836 701788
rect 288892 701786 288916 701788
rect 288972 701786 288996 701788
rect 289052 701786 289076 701788
rect 289132 701786 289156 701788
rect 289212 701786 289236 701788
rect 289292 701786 289316 701788
rect 289372 701786 289386 701788
rect 289066 701734 289076 701786
rect 289132 701734 289142 701786
rect 288822 701732 288836 701734
rect 288892 701732 288916 701734
rect 288972 701732 288996 701734
rect 289052 701732 289076 701734
rect 289132 701732 289156 701734
rect 289212 701732 289236 701734
rect 289292 701732 289316 701734
rect 289372 701732 289386 701734
rect 288822 701712 289386 701732
rect 288822 700700 289386 700720
rect 288822 700698 288836 700700
rect 288892 700698 288916 700700
rect 288972 700698 288996 700700
rect 289052 700698 289076 700700
rect 289132 700698 289156 700700
rect 289212 700698 289236 700700
rect 289292 700698 289316 700700
rect 289372 700698 289386 700700
rect 289066 700646 289076 700698
rect 289132 700646 289142 700698
rect 288822 700644 288836 700646
rect 288892 700644 288916 700646
rect 288972 700644 288996 700646
rect 289052 700644 289076 700646
rect 289132 700644 289156 700646
rect 289212 700644 289236 700646
rect 289292 700644 289316 700646
rect 289372 700644 289386 700646
rect 288822 700624 289386 700644
rect 300136 700398 300164 703520
rect 324822 701788 325386 701808
rect 324822 701786 324836 701788
rect 324892 701786 324916 701788
rect 324972 701786 324996 701788
rect 325052 701786 325076 701788
rect 325132 701786 325156 701788
rect 325212 701786 325236 701788
rect 325292 701786 325316 701788
rect 325372 701786 325386 701788
rect 325066 701734 325076 701786
rect 325132 701734 325142 701786
rect 324822 701732 324836 701734
rect 324892 701732 324916 701734
rect 324972 701732 324996 701734
rect 325052 701732 325076 701734
rect 325132 701732 325156 701734
rect 325212 701732 325236 701734
rect 325292 701732 325316 701734
rect 325372 701732 325386 701734
rect 324822 701712 325386 701732
rect 306822 701244 307386 701264
rect 306822 701242 306836 701244
rect 306892 701242 306916 701244
rect 306972 701242 306996 701244
rect 307052 701242 307076 701244
rect 307132 701242 307156 701244
rect 307212 701242 307236 701244
rect 307292 701242 307316 701244
rect 307372 701242 307386 701244
rect 307066 701190 307076 701242
rect 307132 701190 307142 701242
rect 306822 701188 306836 701190
rect 306892 701188 306916 701190
rect 306972 701188 306996 701190
rect 307052 701188 307076 701190
rect 307132 701188 307156 701190
rect 307212 701188 307236 701190
rect 307292 701188 307316 701190
rect 307372 701188 307386 701190
rect 306822 701168 307386 701188
rect 317972 700936 318024 700942
rect 317972 700878 318024 700884
rect 313188 700868 313240 700874
rect 313188 700810 313240 700816
rect 292580 700392 292632 700398
rect 292580 700334 292632 700340
rect 292672 700392 292724 700398
rect 292672 700334 292724 700340
rect 300124 700392 300176 700398
rect 300124 700334 300176 700340
rect 300216 700392 300268 700398
rect 300216 700334 300268 700340
rect 292592 700233 292620 700334
rect 292578 700224 292634 700233
rect 292578 700159 292634 700168
rect 289542 700088 289598 700097
rect 280066 700023 280122 700032
rect 283748 700052 283800 700058
rect 267648 699994 267700 700000
rect 265900 699984 265952 699990
rect 265900 699926 265952 699932
rect 263876 699780 263928 699786
rect 263876 699722 263928 699728
rect 263598 699544 263654 699553
rect 263598 699479 263654 699488
rect 261390 699000 261446 699009
rect 261390 698935 261446 698944
rect 261404 695994 261432 698935
rect 263612 698902 263640 699479
rect 263690 699408 263746 699417
rect 263690 699343 263746 699352
rect 263704 699145 263732 699343
rect 263690 699136 263746 699145
rect 263690 699071 263746 699080
rect 263888 699009 263916 699722
rect 263874 699000 263930 699009
rect 263874 698935 263930 698944
rect 263600 698896 263652 698902
rect 263692 698896 263744 698902
rect 263600 698838 263652 698844
rect 263690 698864 263692 698873
rect 263744 698864 263746 698873
rect 263690 698799 263746 698808
rect 261142 695966 261432 695994
rect 265912 695980 265940 699926
rect 270500 699848 270552 699854
rect 270498 699816 270500 699825
rect 270592 699848 270644 699854
rect 270552 699816 270554 699825
rect 270592 699790 270644 699796
rect 273166 699816 273222 699825
rect 270498 699751 270554 699760
rect 270604 695980 270632 699790
rect 273166 699751 273222 699760
rect 273536 699780 273588 699786
rect 273180 699718 273208 699751
rect 273536 699722 273588 699728
rect 275744 699780 275796 699786
rect 275744 699722 275796 699728
rect 273168 699712 273220 699718
rect 273168 699654 273220 699660
rect 273260 699440 273312 699446
rect 273352 699440 273404 699446
rect 273260 699382 273312 699388
rect 273350 699408 273352 699417
rect 273404 699408 273406 699417
rect 273272 699145 273300 699382
rect 273350 699343 273406 699352
rect 273258 699136 273314 699145
rect 270822 699068 271386 699088
rect 273258 699071 273314 699080
rect 270822 699066 270836 699068
rect 270892 699066 270916 699068
rect 270972 699066 270996 699068
rect 271052 699066 271076 699068
rect 271132 699066 271156 699068
rect 271212 699066 271236 699068
rect 271292 699066 271316 699068
rect 271372 699066 271386 699068
rect 271066 699014 271076 699066
rect 271132 699014 271142 699066
rect 270822 699012 270836 699014
rect 270892 699012 270916 699014
rect 270972 699012 270996 699014
rect 271052 699012 271076 699014
rect 271132 699012 271156 699014
rect 271212 699012 271236 699014
rect 271292 699012 271316 699014
rect 271372 699012 271386 699014
rect 270822 698992 271386 699012
rect 273548 699009 273576 699722
rect 273534 699000 273590 699009
rect 273534 698935 273590 698944
rect 275756 695994 275784 699722
rect 275402 695966 275784 695994
rect 280080 695980 280108 700023
rect 283748 699994 283800 700000
rect 283840 700052 283892 700058
rect 283840 699994 283892 700000
rect 289452 700052 289504 700058
rect 292684 700074 292712 700334
rect 298650 700224 298706 700233
rect 298650 700159 298706 700168
rect 289542 700023 289544 700032
rect 289452 699994 289504 700000
rect 289596 700023 289598 700032
rect 292592 700046 292712 700074
rect 289544 699994 289596 700000
rect 283760 699938 283788 699994
rect 283760 699910 284340 699938
rect 282920 699712 282972 699718
rect 282920 699654 282972 699660
rect 282932 699553 282960 699654
rect 282734 699544 282790 699553
rect 282918 699544 282974 699553
rect 282790 699502 282868 699530
rect 282734 699479 282790 699488
rect 282734 699408 282790 699417
rect 282734 699343 282790 699352
rect 282748 699174 282776 699343
rect 282840 699174 282868 699502
rect 282918 699479 282974 699488
rect 282920 699440 282972 699446
rect 283012 699440 283064 699446
rect 282920 699382 282972 699388
rect 283010 699408 283012 699417
rect 283064 699408 283066 699417
rect 282932 699258 282960 699382
rect 283010 699343 283066 699352
rect 282932 699230 283144 699258
rect 282736 699168 282788 699174
rect 282736 699110 282788 699116
rect 282828 699168 282880 699174
rect 282828 699110 282880 699116
rect 282920 699168 282972 699174
rect 282920 699110 282972 699116
rect 283012 699168 283064 699174
rect 283012 699110 283064 699116
rect 282932 698873 282960 699110
rect 282918 698864 282974 698873
rect 282918 698799 282974 698808
rect 283024 698601 283052 699110
rect 283116 698986 283144 699230
rect 283286 699000 283342 699009
rect 283116 698958 283286 698986
rect 283286 698935 283342 698944
rect 283010 698592 283066 698601
rect 283010 698527 283066 698536
rect 284312 695994 284340 699910
rect 288440 699712 288492 699718
rect 288440 699654 288492 699660
rect 288452 699145 288480 699654
rect 288822 699612 289386 699632
rect 288822 699610 288836 699612
rect 288892 699610 288916 699612
rect 288972 699610 288996 699612
rect 289052 699610 289076 699612
rect 289132 699610 289156 699612
rect 289212 699610 289236 699612
rect 289292 699610 289316 699612
rect 289372 699610 289386 699612
rect 289066 699558 289076 699610
rect 289132 699558 289142 699610
rect 288822 699556 288836 699558
rect 288892 699556 288916 699558
rect 288972 699556 288996 699558
rect 289052 699556 289076 699558
rect 289132 699556 289156 699558
rect 289212 699556 289236 699558
rect 289292 699556 289316 699558
rect 289372 699556 289386 699558
rect 288822 699536 289386 699556
rect 288438 699136 288494 699145
rect 288438 699071 288494 699080
rect 288822 698524 289386 698544
rect 288822 698522 288836 698524
rect 288892 698522 288916 698524
rect 288972 698522 288996 698524
rect 289052 698522 289076 698524
rect 289132 698522 289156 698524
rect 289212 698522 289236 698524
rect 289292 698522 289316 698524
rect 289372 698522 289386 698524
rect 289066 698470 289076 698522
rect 289132 698470 289142 698522
rect 288822 698468 288836 698470
rect 288892 698468 288916 698470
rect 288972 698468 288996 698470
rect 289052 698468 289076 698470
rect 289132 698468 289156 698470
rect 289212 698468 289236 698470
rect 289292 698468 289316 698470
rect 289372 698468 289386 698470
rect 288822 698448 289386 698468
rect 289464 695994 289492 699994
rect 292302 699952 292358 699961
rect 292302 699887 292358 699896
rect 292316 699786 292344 699887
rect 292488 699848 292540 699854
rect 292486 699816 292488 699825
rect 292540 699816 292542 699825
rect 292304 699780 292356 699786
rect 292486 699751 292542 699760
rect 292304 699722 292356 699728
rect 292592 699718 292620 700046
rect 292670 699952 292726 699961
rect 292670 699887 292726 699896
rect 292684 699786 292712 699887
rect 292672 699780 292724 699786
rect 292672 699722 292724 699728
rect 292580 699712 292632 699718
rect 292580 699654 292632 699660
rect 289726 699544 289782 699553
rect 289726 699479 289782 699488
rect 292670 699544 292726 699553
rect 292670 699479 292726 699488
rect 289740 696862 289768 699479
rect 292684 699446 292712 699479
rect 292672 699440 292724 699446
rect 292672 699382 292724 699388
rect 294050 699408 294106 699417
rect 294050 699343 294106 699352
rect 292396 699168 292448 699174
rect 292394 699136 292396 699145
rect 292488 699168 292540 699174
rect 292448 699136 292450 699145
rect 292488 699110 292540 699116
rect 292394 699071 292450 699080
rect 292500 699009 292528 699110
rect 292486 699000 292542 699009
rect 292486 698935 292542 698944
rect 289728 696856 289780 696862
rect 289728 696798 289780 696804
rect 294064 695994 294092 699343
rect 298664 695994 298692 700159
rect 300228 698873 300256 700334
rect 308496 700256 308548 700262
rect 308496 700198 308548 700204
rect 306822 700156 307386 700176
rect 306822 700154 306836 700156
rect 306892 700154 306916 700156
rect 306972 700154 306996 700156
rect 307052 700154 307076 700156
rect 307132 700154 307156 700156
rect 307212 700154 307236 700156
rect 307292 700154 307316 700156
rect 307372 700154 307386 700156
rect 307066 700102 307076 700154
rect 307132 700102 307142 700154
rect 306822 700100 306836 700102
rect 306892 700100 306916 700102
rect 306972 700100 306996 700102
rect 307052 700100 307076 700102
rect 307132 700100 307156 700102
rect 307212 700100 307236 700102
rect 307292 700100 307316 700102
rect 307372 700100 307386 700102
rect 306822 700080 307386 700100
rect 302054 699952 302110 699961
rect 302054 699887 302056 699896
rect 302108 699887 302110 699896
rect 303618 699952 303674 699961
rect 303618 699887 303674 699896
rect 302056 699858 302108 699864
rect 301964 699848 302016 699854
rect 301962 699816 301964 699825
rect 302016 699816 302018 699825
rect 301962 699751 302018 699760
rect 302148 699440 302200 699446
rect 302148 699382 302200 699388
rect 302160 699145 302188 699382
rect 302146 699136 302202 699145
rect 302146 699071 302202 699080
rect 300214 698864 300270 698873
rect 300214 698799 300270 698808
rect 303632 695994 303660 699887
rect 306822 699068 307386 699088
rect 306822 699066 306836 699068
rect 306892 699066 306916 699068
rect 306972 699066 306996 699068
rect 307052 699066 307076 699068
rect 307132 699066 307156 699068
rect 307212 699066 307236 699068
rect 307292 699066 307316 699068
rect 307372 699066 307386 699068
rect 307066 699014 307076 699066
rect 307132 699014 307142 699066
rect 306822 699012 306836 699014
rect 306892 699012 306916 699014
rect 306972 699012 306996 699014
rect 307052 699012 307076 699014
rect 307132 699012 307156 699014
rect 307212 699012 307236 699014
rect 307292 699012 307316 699014
rect 307372 699012 307386 699014
rect 306822 698992 307386 699012
rect 306380 698896 306432 698902
rect 306378 698864 306380 698873
rect 306432 698864 306434 698873
rect 306378 698799 306434 698808
rect 284312 695966 284878 695994
rect 289464 695966 289570 695994
rect 294064 695966 294354 695994
rect 298664 695966 299046 695994
rect 303632 695966 303738 695994
rect 308508 695980 308536 700198
rect 311900 699712 311952 699718
rect 311900 699654 311952 699660
rect 311912 699145 311940 699654
rect 311898 699136 311954 699145
rect 311898 699071 311954 699080
rect 313200 695980 313228 700810
rect 317984 695980 318012 700878
rect 322664 700800 322716 700806
rect 322664 700742 322716 700748
rect 322676 695980 322704 700742
rect 324822 700700 325386 700720
rect 324822 700698 324836 700700
rect 324892 700698 324916 700700
rect 324972 700698 324996 700700
rect 325052 700698 325076 700700
rect 325132 700698 325156 700700
rect 325212 700698 325236 700700
rect 325292 700698 325316 700700
rect 325372 700698 325386 700700
rect 325066 700646 325076 700698
rect 325132 700646 325142 700698
rect 324822 700644 324836 700646
rect 324892 700644 324916 700646
rect 324972 700644 324996 700646
rect 325052 700644 325076 700646
rect 325132 700644 325156 700646
rect 325212 700644 325236 700646
rect 325292 700644 325316 700646
rect 325372 700644 325386 700646
rect 324822 700624 325386 700644
rect 332140 700460 332192 700466
rect 332140 700402 332192 700408
rect 327448 700324 327500 700330
rect 327448 700266 327500 700272
rect 324822 699612 325386 699632
rect 324822 699610 324836 699612
rect 324892 699610 324916 699612
rect 324972 699610 324996 699612
rect 325052 699610 325076 699612
rect 325132 699610 325156 699612
rect 325212 699610 325236 699612
rect 325292 699610 325316 699612
rect 325372 699610 325386 699612
rect 325066 699558 325076 699610
rect 325132 699558 325142 699610
rect 324822 699556 324836 699558
rect 324892 699556 324916 699558
rect 324972 699556 324996 699558
rect 325052 699556 325076 699558
rect 325132 699556 325156 699558
rect 325212 699556 325236 699558
rect 325292 699556 325316 699558
rect 325372 699556 325386 699558
rect 324822 699536 325386 699556
rect 325516 699168 325568 699174
rect 325514 699136 325516 699145
rect 325700 699168 325752 699174
rect 325568 699136 325570 699145
rect 325514 699071 325570 699080
rect 325698 699136 325700 699145
rect 325752 699136 325754 699145
rect 325698 699071 325754 699080
rect 325608 698896 325660 698902
rect 325606 698864 325608 698873
rect 325660 698864 325662 698873
rect 325606 698799 325662 698808
rect 324822 698524 325386 698544
rect 324822 698522 324836 698524
rect 324892 698522 324916 698524
rect 324972 698522 324996 698524
rect 325052 698522 325076 698524
rect 325132 698522 325156 698524
rect 325212 698522 325236 698524
rect 325292 698522 325316 698524
rect 325372 698522 325386 698524
rect 325066 698470 325076 698522
rect 325132 698470 325142 698522
rect 324822 698468 324836 698470
rect 324892 698468 324916 698470
rect 324972 698468 324996 698470
rect 325052 698468 325076 698470
rect 325132 698468 325156 698470
rect 325212 698468 325236 698470
rect 325292 698468 325316 698470
rect 325372 698468 325386 698470
rect 324822 698448 325386 698468
rect 327460 695980 327488 700266
rect 331220 699712 331272 699718
rect 331220 699654 331272 699660
rect 331232 699145 331260 699654
rect 331218 699136 331274 699145
rect 331218 699071 331274 699080
rect 332152 695980 332180 700402
rect 332520 699786 332548 703520
rect 342822 701244 343386 701264
rect 342822 701242 342836 701244
rect 342892 701242 342916 701244
rect 342972 701242 342996 701244
rect 343052 701242 343076 701244
rect 343132 701242 343156 701244
rect 343212 701242 343236 701244
rect 343292 701242 343316 701244
rect 343372 701242 343386 701244
rect 343066 701190 343076 701242
rect 343132 701190 343142 701242
rect 342822 701188 342836 701190
rect 342892 701188 342916 701190
rect 342972 701188 342996 701190
rect 343052 701188 343076 701190
rect 343132 701188 343156 701190
rect 343212 701188 343236 701190
rect 343292 701188 343316 701190
rect 343372 701188 343386 701190
rect 342822 701168 343386 701188
rect 336922 701040 336978 701049
rect 336922 700975 336978 700984
rect 332508 699780 332560 699786
rect 332508 699722 332560 699728
rect 336936 695980 336964 700975
rect 346306 700496 346362 700505
rect 346306 700431 346362 700440
rect 341614 700360 341670 700369
rect 341614 700295 341670 700304
rect 340788 699916 340840 699922
rect 340788 699858 340840 699864
rect 340800 699174 340828 699858
rect 340788 699168 340840 699174
rect 340788 699110 340840 699116
rect 340696 698896 340748 698902
rect 340694 698864 340696 698873
rect 340748 698864 340750 698873
rect 340694 698799 340750 698808
rect 341628 695980 341656 700295
rect 342822 700156 343386 700176
rect 342822 700154 342836 700156
rect 342892 700154 342916 700156
rect 342972 700154 342996 700156
rect 343052 700154 343076 700156
rect 343132 700154 343156 700156
rect 343212 700154 343236 700156
rect 343292 700154 343316 700156
rect 343372 700154 343386 700156
rect 343066 700102 343076 700154
rect 343132 700102 343142 700154
rect 342822 700100 342836 700102
rect 342892 700100 342916 700102
rect 342972 700100 342996 700102
rect 343052 700100 343076 700102
rect 343132 700100 343156 700102
rect 343212 700100 343236 700102
rect 343292 700100 343316 700102
rect 343372 700100 343386 700102
rect 342822 700080 343386 700100
rect 343548 699712 343600 699718
rect 343548 699654 343600 699660
rect 343560 699145 343588 699654
rect 343546 699136 343602 699145
rect 342822 699068 343386 699088
rect 343546 699071 343602 699080
rect 342822 699066 342836 699068
rect 342892 699066 342916 699068
rect 342972 699066 342996 699068
rect 343052 699066 343076 699068
rect 343132 699066 343156 699068
rect 343212 699066 343236 699068
rect 343292 699066 343316 699068
rect 343372 699066 343386 699068
rect 343066 699014 343076 699066
rect 343132 699014 343142 699066
rect 342822 699012 342836 699014
rect 342892 699012 342916 699014
rect 342972 699012 342996 699014
rect 343052 699012 343076 699014
rect 343132 699012 343156 699014
rect 343212 699012 343236 699014
rect 343292 699012 343316 699014
rect 343372 699012 343386 699014
rect 342822 698992 343386 699012
rect 346320 695980 346348 700431
rect 348804 699854 348832 703520
rect 360822 701788 361386 701808
rect 360822 701786 360836 701788
rect 360892 701786 360916 701788
rect 360972 701786 360996 701788
rect 361052 701786 361076 701788
rect 361132 701786 361156 701788
rect 361212 701786 361236 701788
rect 361292 701786 361316 701788
rect 361372 701786 361386 701788
rect 361066 701734 361076 701786
rect 361132 701734 361142 701786
rect 360822 701732 360836 701734
rect 360892 701732 360916 701734
rect 360972 701732 360996 701734
rect 361052 701732 361076 701734
rect 361132 701732 361156 701734
rect 361212 701732 361236 701734
rect 361292 701732 361316 701734
rect 361372 701732 361386 701734
rect 360822 701712 361386 701732
rect 360822 700700 361386 700720
rect 360822 700698 360836 700700
rect 360892 700698 360916 700700
rect 360972 700698 360996 700700
rect 361052 700698 361076 700700
rect 361132 700698 361156 700700
rect 361212 700698 361236 700700
rect 361292 700698 361316 700700
rect 361372 700698 361386 700700
rect 361066 700646 361076 700698
rect 361132 700646 361142 700698
rect 360822 700644 360836 700646
rect 360892 700644 360916 700646
rect 360972 700644 360996 700646
rect 361052 700644 361076 700646
rect 361132 700644 361156 700646
rect 361212 700644 361236 700646
rect 361292 700644 361316 700646
rect 361372 700644 361386 700646
rect 360822 700624 361386 700644
rect 364996 699990 365024 703520
rect 396822 701788 397386 701808
rect 396822 701786 396836 701788
rect 396892 701786 396916 701788
rect 396972 701786 396996 701788
rect 397052 701786 397076 701788
rect 397132 701786 397156 701788
rect 397212 701786 397236 701788
rect 397292 701786 397316 701788
rect 397372 701786 397386 701788
rect 397066 701734 397076 701786
rect 397132 701734 397142 701786
rect 396822 701732 396836 701734
rect 396892 701732 396916 701734
rect 396972 701732 396996 701734
rect 397052 701732 397076 701734
rect 397132 701732 397156 701734
rect 397212 701732 397236 701734
rect 397292 701732 397316 701734
rect 397372 701732 397386 701734
rect 396822 701712 397386 701732
rect 378822 701244 379386 701264
rect 378822 701242 378836 701244
rect 378892 701242 378916 701244
rect 378972 701242 378996 701244
rect 379052 701242 379076 701244
rect 379132 701242 379156 701244
rect 379212 701242 379236 701244
rect 379292 701242 379316 701244
rect 379372 701242 379386 701244
rect 379066 701190 379076 701242
rect 379132 701190 379142 701242
rect 378822 701188 378836 701190
rect 378892 701188 378916 701190
rect 378972 701188 378996 701190
rect 379052 701188 379076 701190
rect 379132 701188 379156 701190
rect 379212 701188 379236 701190
rect 379292 701188 379316 701190
rect 379372 701188 379386 701190
rect 378822 701168 379386 701188
rect 397472 701010 397500 703520
rect 397460 701004 397512 701010
rect 397460 700946 397512 700952
rect 396822 700700 397386 700720
rect 396822 700698 396836 700700
rect 396892 700698 396916 700700
rect 396972 700698 396996 700700
rect 397052 700698 397076 700700
rect 397132 700698 397156 700700
rect 397212 700698 397236 700700
rect 397292 700698 397316 700700
rect 397372 700698 397386 700700
rect 397066 700646 397076 700698
rect 397132 700646 397142 700698
rect 396822 700644 396836 700646
rect 396892 700644 396916 700646
rect 396972 700644 396996 700646
rect 397052 700644 397076 700646
rect 397132 700644 397156 700646
rect 397212 700644 397236 700646
rect 397292 700644 397316 700646
rect 397372 700644 397386 700646
rect 396822 700624 397386 700644
rect 378822 700156 379386 700176
rect 378822 700154 378836 700156
rect 378892 700154 378916 700156
rect 378972 700154 378996 700156
rect 379052 700154 379076 700156
rect 379132 700154 379156 700156
rect 379212 700154 379236 700156
rect 379292 700154 379316 700156
rect 379372 700154 379386 700156
rect 379066 700102 379076 700154
rect 379132 700102 379142 700154
rect 378822 700100 378836 700102
rect 378892 700100 378916 700102
rect 378972 700100 378996 700102
rect 379052 700100 379076 700102
rect 379132 700100 379156 700102
rect 379212 700100 379236 700102
rect 379292 700100 379316 700102
rect 379372 700100 379386 700102
rect 378822 700080 379386 700100
rect 413664 700058 413692 703520
rect 429856 702030 429884 703520
rect 429844 702024 429896 702030
rect 429844 701966 429896 701972
rect 432822 701788 433386 701808
rect 432822 701786 432836 701788
rect 432892 701786 432916 701788
rect 432972 701786 432996 701788
rect 433052 701786 433076 701788
rect 433132 701786 433156 701788
rect 433212 701786 433236 701788
rect 433292 701786 433316 701788
rect 433372 701786 433386 701788
rect 433066 701734 433076 701786
rect 433132 701734 433142 701786
rect 432822 701732 432836 701734
rect 432892 701732 432916 701734
rect 432972 701732 432996 701734
rect 433052 701732 433076 701734
rect 433132 701732 433156 701734
rect 433212 701732 433236 701734
rect 433292 701732 433316 701734
rect 433372 701732 433386 701734
rect 432822 701712 433386 701732
rect 414822 701244 415386 701264
rect 414822 701242 414836 701244
rect 414892 701242 414916 701244
rect 414972 701242 414996 701244
rect 415052 701242 415076 701244
rect 415132 701242 415156 701244
rect 415212 701242 415236 701244
rect 415292 701242 415316 701244
rect 415372 701242 415386 701244
rect 415066 701190 415076 701242
rect 415132 701190 415142 701242
rect 414822 701188 414836 701190
rect 414892 701188 414916 701190
rect 414972 701188 414996 701190
rect 415052 701188 415076 701190
rect 415132 701188 415156 701190
rect 415212 701188 415236 701190
rect 415292 701188 415316 701190
rect 415372 701188 415386 701190
rect 414822 701168 415386 701188
rect 450822 701244 451386 701264
rect 450822 701242 450836 701244
rect 450892 701242 450916 701244
rect 450972 701242 450996 701244
rect 451052 701242 451076 701244
rect 451132 701242 451156 701244
rect 451212 701242 451236 701244
rect 451292 701242 451316 701244
rect 451372 701242 451386 701244
rect 451066 701190 451076 701242
rect 451132 701190 451142 701242
rect 450822 701188 450836 701190
rect 450892 701188 450916 701190
rect 450972 701188 450996 701190
rect 451052 701188 451076 701190
rect 451132 701188 451156 701190
rect 451212 701188 451236 701190
rect 451292 701188 451316 701190
rect 451372 701188 451386 701190
rect 450822 701168 451386 701188
rect 432822 700700 433386 700720
rect 432822 700698 432836 700700
rect 432892 700698 432916 700700
rect 432972 700698 432996 700700
rect 433052 700698 433076 700700
rect 433132 700698 433156 700700
rect 433212 700698 433236 700700
rect 433292 700698 433316 700700
rect 433372 700698 433386 700700
rect 433066 700646 433076 700698
rect 433132 700646 433142 700698
rect 432822 700644 432836 700646
rect 432892 700644 432916 700646
rect 432972 700644 432996 700646
rect 433052 700644 433076 700646
rect 433132 700644 433156 700646
rect 433212 700644 433236 700646
rect 433292 700644 433316 700646
rect 433372 700644 433386 700646
rect 432822 700624 433386 700644
rect 462332 700602 462360 703520
rect 468822 701788 469386 701808
rect 468822 701786 468836 701788
rect 468892 701786 468916 701788
rect 468972 701786 468996 701788
rect 469052 701786 469076 701788
rect 469132 701786 469156 701788
rect 469212 701786 469236 701788
rect 469292 701786 469316 701788
rect 469372 701786 469386 701788
rect 469066 701734 469076 701786
rect 469132 701734 469142 701786
rect 468822 701732 468836 701734
rect 468892 701732 468916 701734
rect 468972 701732 468996 701734
rect 469052 701732 469076 701734
rect 469132 701732 469156 701734
rect 469212 701732 469236 701734
rect 469292 701732 469316 701734
rect 469372 701732 469386 701734
rect 468822 701712 469386 701732
rect 468822 700700 469386 700720
rect 468822 700698 468836 700700
rect 468892 700698 468916 700700
rect 468972 700698 468996 700700
rect 469052 700698 469076 700700
rect 469132 700698 469156 700700
rect 469212 700698 469236 700700
rect 469292 700698 469316 700700
rect 469372 700698 469386 700700
rect 469066 700646 469076 700698
rect 469132 700646 469142 700698
rect 468822 700644 468836 700646
rect 468892 700644 468916 700646
rect 468972 700644 468996 700646
rect 469052 700644 469076 700646
rect 469132 700644 469156 700646
rect 469212 700644 469236 700646
rect 469292 700644 469316 700646
rect 469372 700644 469386 700646
rect 468822 700624 469386 700644
rect 462320 700596 462372 700602
rect 462320 700538 462372 700544
rect 478524 700534 478552 703520
rect 494808 701962 494836 703520
rect 494796 701956 494848 701962
rect 494796 701898 494848 701904
rect 504822 701788 505386 701808
rect 504822 701786 504836 701788
rect 504892 701786 504916 701788
rect 504972 701786 504996 701788
rect 505052 701786 505076 701788
rect 505132 701786 505156 701788
rect 505212 701786 505236 701788
rect 505292 701786 505316 701788
rect 505372 701786 505386 701788
rect 505066 701734 505076 701786
rect 505132 701734 505142 701786
rect 504822 701732 504836 701734
rect 504892 701732 504916 701734
rect 504972 701732 504996 701734
rect 505052 701732 505076 701734
rect 505132 701732 505156 701734
rect 505212 701732 505236 701734
rect 505292 701732 505316 701734
rect 505372 701732 505386 701734
rect 504822 701712 505386 701732
rect 486822 701244 487386 701264
rect 486822 701242 486836 701244
rect 486892 701242 486916 701244
rect 486972 701242 486996 701244
rect 487052 701242 487076 701244
rect 487132 701242 487156 701244
rect 487212 701242 487236 701244
rect 487292 701242 487316 701244
rect 487372 701242 487386 701244
rect 487066 701190 487076 701242
rect 487132 701190 487142 701242
rect 486822 701188 486836 701190
rect 486892 701188 486916 701190
rect 486972 701188 486996 701190
rect 487052 701188 487076 701190
rect 487132 701188 487156 701190
rect 487212 701188 487236 701190
rect 487292 701188 487316 701190
rect 487372 701188 487386 701190
rect 486822 701168 487386 701188
rect 522822 701244 523386 701264
rect 522822 701242 522836 701244
rect 522892 701242 522916 701244
rect 522972 701242 522996 701244
rect 523052 701242 523076 701244
rect 523132 701242 523156 701244
rect 523212 701242 523236 701244
rect 523292 701242 523316 701244
rect 523372 701242 523386 701244
rect 523066 701190 523076 701242
rect 523132 701190 523142 701242
rect 522822 701188 522836 701190
rect 522892 701188 522916 701190
rect 522972 701188 522996 701190
rect 523052 701188 523076 701190
rect 523132 701188 523156 701190
rect 523212 701188 523236 701190
rect 523292 701188 523316 701190
rect 523372 701188 523386 701190
rect 522822 701168 523386 701188
rect 527192 700913 527220 703520
rect 540822 701788 541386 701808
rect 540822 701786 540836 701788
rect 540892 701786 540916 701788
rect 540972 701786 540996 701788
rect 541052 701786 541076 701788
rect 541132 701786 541156 701788
rect 541212 701786 541236 701788
rect 541292 701786 541316 701788
rect 541372 701786 541386 701788
rect 541066 701734 541076 701786
rect 541132 701734 541142 701786
rect 540822 701732 540836 701734
rect 540892 701732 540916 701734
rect 540972 701732 540996 701734
rect 541052 701732 541076 701734
rect 541132 701732 541156 701734
rect 541212 701732 541236 701734
rect 541292 701732 541316 701734
rect 541372 701732 541386 701734
rect 540822 701712 541386 701732
rect 527178 700904 527234 700913
rect 527178 700839 527234 700848
rect 504822 700700 505386 700720
rect 504822 700698 504836 700700
rect 504892 700698 504916 700700
rect 504972 700698 504996 700700
rect 505052 700698 505076 700700
rect 505132 700698 505156 700700
rect 505212 700698 505236 700700
rect 505292 700698 505316 700700
rect 505372 700698 505386 700700
rect 505066 700646 505076 700698
rect 505132 700646 505142 700698
rect 504822 700644 504836 700646
rect 504892 700644 504916 700646
rect 504972 700644 504996 700646
rect 505052 700644 505076 700646
rect 505132 700644 505156 700646
rect 505212 700644 505236 700646
rect 505292 700644 505316 700646
rect 505372 700644 505386 700646
rect 504822 700624 505386 700644
rect 540822 700700 541386 700720
rect 540822 700698 540836 700700
rect 540892 700698 540916 700700
rect 540972 700698 540996 700700
rect 541052 700698 541076 700700
rect 541132 700698 541156 700700
rect 541212 700698 541236 700700
rect 541292 700698 541316 700700
rect 541372 700698 541386 700700
rect 541066 700646 541076 700698
rect 541132 700646 541142 700698
rect 540822 700644 540836 700646
rect 540892 700644 540916 700646
rect 540972 700644 540996 700646
rect 541052 700644 541076 700646
rect 541132 700644 541156 700646
rect 541212 700644 541236 700646
rect 541292 700644 541316 700646
rect 541372 700644 541386 700646
rect 540822 700624 541386 700644
rect 478512 700528 478564 700534
rect 478512 700470 478564 700476
rect 543476 700398 543504 703520
rect 559668 701894 559696 703520
rect 559656 701888 559708 701894
rect 559656 701830 559708 701836
rect 576822 701788 577386 701808
rect 576822 701786 576836 701788
rect 576892 701786 576916 701788
rect 576972 701786 576996 701788
rect 577052 701786 577076 701788
rect 577132 701786 577156 701788
rect 577212 701786 577236 701788
rect 577292 701786 577316 701788
rect 577372 701786 577386 701788
rect 577066 701734 577076 701786
rect 577132 701734 577142 701786
rect 576822 701732 576836 701734
rect 576892 701732 576916 701734
rect 576972 701732 576996 701734
rect 577052 701732 577076 701734
rect 577132 701732 577156 701734
rect 577212 701732 577236 701734
rect 577292 701732 577316 701734
rect 577372 701732 577386 701734
rect 576822 701712 577386 701732
rect 558822 701244 559386 701264
rect 558822 701242 558836 701244
rect 558892 701242 558916 701244
rect 558972 701242 558996 701244
rect 559052 701242 559076 701244
rect 559132 701242 559156 701244
rect 559212 701242 559236 701244
rect 559292 701242 559316 701244
rect 559372 701242 559386 701244
rect 559066 701190 559076 701242
rect 559132 701190 559142 701242
rect 558822 701188 558836 701190
rect 558892 701188 558916 701190
rect 558972 701188 558996 701190
rect 559052 701188 559076 701190
rect 559132 701188 559156 701190
rect 559212 701188 559236 701190
rect 559292 701188 559316 701190
rect 559372 701188 559386 701190
rect 558822 701168 559386 701188
rect 576822 700700 577386 700720
rect 576822 700698 576836 700700
rect 576892 700698 576916 700700
rect 576972 700698 576996 700700
rect 577052 700698 577076 700700
rect 577132 700698 577156 700700
rect 577212 700698 577236 700700
rect 577292 700698 577316 700700
rect 577372 700698 577386 700700
rect 577066 700646 577076 700698
rect 577132 700646 577142 700698
rect 576822 700644 576836 700646
rect 576892 700644 576916 700646
rect 576972 700644 576996 700646
rect 577052 700644 577076 700646
rect 577132 700644 577156 700646
rect 577212 700644 577236 700646
rect 577292 700644 577316 700646
rect 577372 700644 577386 700646
rect 576822 700624 577386 700644
rect 543464 700392 543516 700398
rect 543464 700334 543516 700340
rect 414822 700156 415386 700176
rect 414822 700154 414836 700156
rect 414892 700154 414916 700156
rect 414972 700154 414996 700156
rect 415052 700154 415076 700156
rect 415132 700154 415156 700156
rect 415212 700154 415236 700156
rect 415292 700154 415316 700156
rect 415372 700154 415386 700156
rect 415066 700102 415076 700154
rect 415132 700102 415142 700154
rect 414822 700100 414836 700102
rect 414892 700100 414916 700102
rect 414972 700100 414996 700102
rect 415052 700100 415076 700102
rect 415132 700100 415156 700102
rect 415212 700100 415236 700102
rect 415292 700100 415316 700102
rect 415372 700100 415386 700102
rect 414822 700080 415386 700100
rect 450822 700156 451386 700176
rect 450822 700154 450836 700156
rect 450892 700154 450916 700156
rect 450972 700154 450996 700156
rect 451052 700154 451076 700156
rect 451132 700154 451156 700156
rect 451212 700154 451236 700156
rect 451292 700154 451316 700156
rect 451372 700154 451386 700156
rect 451066 700102 451076 700154
rect 451132 700102 451142 700154
rect 450822 700100 450836 700102
rect 450892 700100 450916 700102
rect 450972 700100 450996 700102
rect 451052 700100 451076 700102
rect 451132 700100 451156 700102
rect 451212 700100 451236 700102
rect 451292 700100 451316 700102
rect 451372 700100 451386 700102
rect 450822 700080 451386 700100
rect 486822 700156 487386 700176
rect 486822 700154 486836 700156
rect 486892 700154 486916 700156
rect 486972 700154 486996 700156
rect 487052 700154 487076 700156
rect 487132 700154 487156 700156
rect 487212 700154 487236 700156
rect 487292 700154 487316 700156
rect 487372 700154 487386 700156
rect 487066 700102 487076 700154
rect 487132 700102 487142 700154
rect 486822 700100 486836 700102
rect 486892 700100 486916 700102
rect 486972 700100 486996 700102
rect 487052 700100 487076 700102
rect 487132 700100 487156 700102
rect 487212 700100 487236 700102
rect 487292 700100 487316 700102
rect 487372 700100 487386 700102
rect 486822 700080 487386 700100
rect 522822 700156 523386 700176
rect 522822 700154 522836 700156
rect 522892 700154 522916 700156
rect 522972 700154 522996 700156
rect 523052 700154 523076 700156
rect 523132 700154 523156 700156
rect 523212 700154 523236 700156
rect 523292 700154 523316 700156
rect 523372 700154 523386 700156
rect 523066 700102 523076 700154
rect 523132 700102 523142 700154
rect 522822 700100 522836 700102
rect 522892 700100 522916 700102
rect 522972 700100 522996 700102
rect 523052 700100 523076 700102
rect 523132 700100 523156 700102
rect 523212 700100 523236 700102
rect 523292 700100 523316 700102
rect 523372 700100 523386 700102
rect 522822 700080 523386 700100
rect 558822 700156 559386 700176
rect 558822 700154 558836 700156
rect 558892 700154 558916 700156
rect 558972 700154 558996 700156
rect 559052 700154 559076 700156
rect 559132 700154 559156 700156
rect 559212 700154 559236 700156
rect 559292 700154 559316 700156
rect 559372 700154 559386 700156
rect 559066 700102 559076 700154
rect 559132 700102 559142 700154
rect 558822 700100 558836 700102
rect 558892 700100 558916 700102
rect 558972 700100 558996 700102
rect 559052 700100 559076 700102
rect 559132 700100 559156 700102
rect 559212 700100 559236 700102
rect 559292 700100 559316 700102
rect 559372 700100 559386 700102
rect 558822 700080 559386 700100
rect 413652 700052 413704 700058
rect 413652 699994 413704 700000
rect 364984 699984 365036 699990
rect 364984 699926 365036 699932
rect 348792 699848 348844 699854
rect 348792 699790 348844 699796
rect 374000 699712 374052 699718
rect 374000 699654 374052 699660
rect 360822 699612 361386 699632
rect 360822 699610 360836 699612
rect 360892 699610 360916 699612
rect 360972 699610 360996 699612
rect 361052 699610 361076 699612
rect 361132 699610 361156 699612
rect 361212 699610 361236 699612
rect 361292 699610 361316 699612
rect 361372 699610 361386 699612
rect 361066 699558 361076 699610
rect 361132 699558 361142 699610
rect 360822 699556 360836 699558
rect 360892 699556 360916 699558
rect 360972 699556 360996 699558
rect 361052 699556 361076 699558
rect 361132 699556 361156 699558
rect 361212 699556 361236 699558
rect 361292 699556 361316 699558
rect 361372 699556 361386 699558
rect 360822 699536 361386 699556
rect 354496 699168 354548 699174
rect 354494 699136 354496 699145
rect 354548 699136 354550 699145
rect 354494 699071 354550 699080
rect 354588 698896 354640 698902
rect 354586 698864 354588 698873
rect 354640 698864 354642 698873
rect 354586 698799 354642 698808
rect 360822 698524 361386 698544
rect 360822 698522 360836 698524
rect 360892 698522 360916 698524
rect 360972 698522 360996 698524
rect 361052 698522 361076 698524
rect 361132 698522 361156 698524
rect 361212 698522 361236 698524
rect 361292 698522 361316 698524
rect 361372 698522 361386 698524
rect 361066 698470 361076 698522
rect 361132 698470 361142 698522
rect 360822 698468 360836 698470
rect 360892 698468 360916 698470
rect 360972 698468 360996 698470
rect 361052 698468 361076 698470
rect 361132 698468 361156 698470
rect 361212 698468 361236 698470
rect 361292 698468 361316 698470
rect 361372 698468 361386 698470
rect 360822 698448 361386 698468
rect 351092 698284 351144 698290
rect 351092 698226 351144 698232
rect 351104 695980 351132 698226
rect 365260 698216 365312 698222
rect 365260 698158 365312 698164
rect 360568 696720 360620 696726
rect 360568 696662 360620 696668
rect 360580 695980 360608 696662
rect 365272 695980 365300 698158
rect 374012 696930 374040 699654
rect 396822 699612 397386 699632
rect 396822 699610 396836 699612
rect 396892 699610 396916 699612
rect 396972 699610 396996 699612
rect 397052 699610 397076 699612
rect 397132 699610 397156 699612
rect 397212 699610 397236 699612
rect 397292 699610 397316 699612
rect 397372 699610 397386 699612
rect 397066 699558 397076 699610
rect 397132 699558 397142 699610
rect 396822 699556 396836 699558
rect 396892 699556 396916 699558
rect 396972 699556 396996 699558
rect 397052 699556 397076 699558
rect 397132 699556 397156 699558
rect 397212 699556 397236 699558
rect 397292 699556 397316 699558
rect 397372 699556 397386 699558
rect 396822 699536 397386 699556
rect 432822 699612 433386 699632
rect 432822 699610 432836 699612
rect 432892 699610 432916 699612
rect 432972 699610 432996 699612
rect 433052 699610 433076 699612
rect 433132 699610 433156 699612
rect 433212 699610 433236 699612
rect 433292 699610 433316 699612
rect 433372 699610 433386 699612
rect 433066 699558 433076 699610
rect 433132 699558 433142 699610
rect 432822 699556 432836 699558
rect 432892 699556 432916 699558
rect 432972 699556 432996 699558
rect 433052 699556 433076 699558
rect 433132 699556 433156 699558
rect 433212 699556 433236 699558
rect 433292 699556 433316 699558
rect 433372 699556 433386 699558
rect 432822 699536 433386 699556
rect 468822 699612 469386 699632
rect 468822 699610 468836 699612
rect 468892 699610 468916 699612
rect 468972 699610 468996 699612
rect 469052 699610 469076 699612
rect 469132 699610 469156 699612
rect 469212 699610 469236 699612
rect 469292 699610 469316 699612
rect 469372 699610 469386 699612
rect 469066 699558 469076 699610
rect 469132 699558 469142 699610
rect 468822 699556 468836 699558
rect 468892 699556 468916 699558
rect 468972 699556 468996 699558
rect 469052 699556 469076 699558
rect 469132 699556 469156 699558
rect 469212 699556 469236 699558
rect 469292 699556 469316 699558
rect 469372 699556 469386 699558
rect 468822 699536 469386 699556
rect 504822 699612 505386 699632
rect 504822 699610 504836 699612
rect 504892 699610 504916 699612
rect 504972 699610 504996 699612
rect 505052 699610 505076 699612
rect 505132 699610 505156 699612
rect 505212 699610 505236 699612
rect 505292 699610 505316 699612
rect 505372 699610 505386 699612
rect 505066 699558 505076 699610
rect 505132 699558 505142 699610
rect 504822 699556 504836 699558
rect 504892 699556 504916 699558
rect 504972 699556 504996 699558
rect 505052 699556 505076 699558
rect 505132 699556 505156 699558
rect 505212 699556 505236 699558
rect 505292 699556 505316 699558
rect 505372 699556 505386 699558
rect 504822 699536 505386 699556
rect 540822 699612 541386 699632
rect 540822 699610 540836 699612
rect 540892 699610 540916 699612
rect 540972 699610 540996 699612
rect 541052 699610 541076 699612
rect 541132 699610 541156 699612
rect 541212 699610 541236 699612
rect 541292 699610 541316 699612
rect 541372 699610 541386 699612
rect 541066 699558 541076 699610
rect 541132 699558 541142 699610
rect 540822 699556 540836 699558
rect 540892 699556 540916 699558
rect 540972 699556 540996 699558
rect 541052 699556 541076 699558
rect 541132 699556 541156 699558
rect 541212 699556 541236 699558
rect 541292 699556 541316 699558
rect 541372 699556 541386 699558
rect 540822 699536 541386 699556
rect 576822 699612 577386 699632
rect 576822 699610 576836 699612
rect 576892 699610 576916 699612
rect 576972 699610 576996 699612
rect 577052 699610 577076 699612
rect 577132 699610 577156 699612
rect 577212 699610 577236 699612
rect 577292 699610 577316 699612
rect 577372 699610 577386 699612
rect 577066 699558 577076 699610
rect 577132 699558 577142 699610
rect 576822 699556 576836 699558
rect 576892 699556 576916 699558
rect 576972 699556 576996 699558
rect 577052 699556 577076 699558
rect 577132 699556 577156 699558
rect 577212 699556 577236 699558
rect 577292 699556 577316 699558
rect 577372 699556 577386 699558
rect 576822 699536 577386 699556
rect 403164 699508 403216 699514
rect 403164 699450 403216 699456
rect 404268 699508 404320 699514
rect 404268 699450 404320 699456
rect 417332 699508 417384 699514
rect 417332 699450 417384 699456
rect 378822 699068 379386 699088
rect 378822 699066 378836 699068
rect 378892 699066 378916 699068
rect 378972 699066 378996 699068
rect 379052 699066 379076 699068
rect 379132 699066 379156 699068
rect 379212 699066 379236 699068
rect 379292 699066 379316 699068
rect 379372 699066 379386 699068
rect 379066 699014 379076 699066
rect 379132 699014 379142 699066
rect 378822 699012 378836 699014
rect 378892 699012 378916 699014
rect 378972 699012 378996 699014
rect 379052 699012 379076 699014
rect 379132 699012 379156 699014
rect 379212 699012 379236 699014
rect 379292 699012 379316 699014
rect 379372 699012 379386 699014
rect 378822 698992 379386 699012
rect 396822 698524 397386 698544
rect 396822 698522 396836 698524
rect 396892 698522 396916 698524
rect 396972 698522 396996 698524
rect 397052 698522 397076 698524
rect 397132 698522 397156 698524
rect 397212 698522 397236 698524
rect 397292 698522 397316 698524
rect 397372 698522 397386 698524
rect 397066 698470 397076 698522
rect 397132 698470 397142 698522
rect 396822 698468 396836 698470
rect 396892 698468 396916 698470
rect 396972 698468 396996 698470
rect 397052 698468 397076 698470
rect 397132 698468 397156 698470
rect 397212 698468 397236 698470
rect 397292 698468 397316 698470
rect 397372 698468 397386 698470
rect 396822 698448 397386 698468
rect 379520 698012 379572 698018
rect 379520 697954 379572 697960
rect 374000 696924 374052 696930
rect 374000 696866 374052 696872
rect 374828 696924 374880 696930
rect 374828 696866 374880 696872
rect 374840 696590 374868 696866
rect 374736 696584 374788 696590
rect 374736 696526 374788 696532
rect 374828 696584 374880 696590
rect 374828 696526 374880 696532
rect 374748 695980 374776 696526
rect 379532 695980 379560 697954
rect 393688 697876 393740 697882
rect 393688 697818 393740 697824
rect 388996 696720 389048 696726
rect 388996 696662 389048 696668
rect 389008 695980 389036 696662
rect 393700 695980 393728 697818
rect 398380 697808 398432 697814
rect 398380 697750 398432 697756
rect 398392 695980 398420 697750
rect 403176 695980 403204 699450
rect 404280 696794 404308 699450
rect 407948 699372 408000 699378
rect 407948 699314 408000 699320
rect 407960 697678 407988 699314
rect 414822 699068 415386 699088
rect 414822 699066 414836 699068
rect 414892 699066 414916 699068
rect 414972 699066 414996 699068
rect 415052 699066 415076 699068
rect 415132 699066 415156 699068
rect 415212 699066 415236 699068
rect 415292 699066 415316 699068
rect 415372 699066 415386 699068
rect 415066 699014 415076 699066
rect 415132 699014 415142 699066
rect 414822 699012 414836 699014
rect 414892 699012 414916 699014
rect 414972 699012 414996 699014
rect 415052 699012 415076 699014
rect 415132 699012 415156 699014
rect 415212 699012 415236 699014
rect 415292 699012 415316 699014
rect 415372 699012 415386 699014
rect 414822 698992 415386 699012
rect 407856 697672 407908 697678
rect 407856 697614 407908 697620
rect 407948 697672 408000 697678
rect 407948 697614 408000 697620
rect 404268 696788 404320 696794
rect 404268 696730 404320 696736
rect 407868 695980 407896 697614
rect 412640 696176 412692 696182
rect 412640 696118 412692 696124
rect 412652 695980 412680 696118
rect 417344 695980 417372 699450
rect 431592 699440 431644 699446
rect 431592 699382 431644 699388
rect 422116 697536 422168 697542
rect 422116 697478 422168 697484
rect 422128 695980 422156 697478
rect 431604 695980 431632 699382
rect 577872 699304 577924 699310
rect 530950 699272 531006 699281
rect 445760 699236 445812 699242
rect 577872 699246 577924 699252
rect 530950 699207 531006 699216
rect 445760 699178 445812 699184
rect 432822 698524 433386 698544
rect 432822 698522 432836 698524
rect 432892 698522 432916 698524
rect 432972 698522 432996 698524
rect 433052 698522 433076 698524
rect 433132 698522 433156 698524
rect 433212 698522 433236 698524
rect 433292 698522 433316 698524
rect 433372 698522 433386 698524
rect 433066 698470 433076 698522
rect 433132 698470 433142 698522
rect 432822 698468 432836 698470
rect 432892 698468 432916 698470
rect 432972 698468 432996 698470
rect 433052 698468 433076 698470
rect 433132 698468 433156 698470
rect 433212 698468 433236 698470
rect 433292 698468 433316 698470
rect 433372 698468 433386 698470
rect 432822 698448 433386 698468
rect 436284 697400 436336 697406
rect 436284 697342 436336 697348
rect 436296 695980 436324 697342
rect 445772 695980 445800 699178
rect 450822 699068 451386 699088
rect 450822 699066 450836 699068
rect 450892 699066 450916 699068
rect 450972 699066 450996 699068
rect 451052 699066 451076 699068
rect 451132 699066 451156 699068
rect 451212 699066 451236 699068
rect 451292 699066 451316 699068
rect 451372 699066 451386 699068
rect 451066 699014 451076 699066
rect 451132 699014 451142 699066
rect 450822 699012 450836 699014
rect 450892 699012 450916 699014
rect 450972 699012 450996 699014
rect 451052 699012 451076 699014
rect 451132 699012 451156 699014
rect 451212 699012 451236 699014
rect 451292 699012 451316 699014
rect 451372 699012 451386 699014
rect 450822 698992 451386 699012
rect 486822 699068 487386 699088
rect 486822 699066 486836 699068
rect 486892 699066 486916 699068
rect 486972 699066 486996 699068
rect 487052 699066 487076 699068
rect 487132 699066 487156 699068
rect 487212 699066 487236 699068
rect 487292 699066 487316 699068
rect 487372 699066 487386 699068
rect 487066 699014 487076 699066
rect 487132 699014 487142 699066
rect 486822 699012 486836 699014
rect 486892 699012 486916 699014
rect 486972 699012 486996 699014
rect 487052 699012 487076 699014
rect 487132 699012 487156 699014
rect 487212 699012 487236 699014
rect 487292 699012 487316 699014
rect 487372 699012 487386 699014
rect 486822 698992 487386 699012
rect 522822 699068 523386 699088
rect 522822 699066 522836 699068
rect 522892 699066 522916 699068
rect 522972 699066 522996 699068
rect 523052 699066 523076 699068
rect 523132 699066 523156 699068
rect 523212 699066 523236 699068
rect 523292 699066 523316 699068
rect 523372 699066 523386 699068
rect 523066 699014 523076 699066
rect 523132 699014 523142 699066
rect 522822 699012 522836 699014
rect 522892 699012 522916 699014
rect 522972 699012 522996 699014
rect 523052 699012 523076 699014
rect 523132 699012 523156 699014
rect 523212 699012 523236 699014
rect 523292 699012 523316 699014
rect 523372 699012 523386 699014
rect 522822 698992 523386 699012
rect 526258 698864 526314 698873
rect 474188 698828 474240 698834
rect 526258 698799 526314 698808
rect 474188 698770 474240 698776
rect 468822 698524 469386 698544
rect 468822 698522 468836 698524
rect 468892 698522 468916 698524
rect 468972 698522 468996 698524
rect 469052 698522 469076 698524
rect 469132 698522 469156 698524
rect 469212 698522 469236 698524
rect 469292 698522 469316 698524
rect 469372 698522 469386 698524
rect 469066 698470 469076 698522
rect 469132 698470 469142 698522
rect 468822 698468 468836 698470
rect 468892 698468 468916 698470
rect 468972 698468 468996 698470
rect 469052 698468 469076 698470
rect 469132 698468 469156 698470
rect 469212 698468 469236 698470
rect 469292 698468 469316 698470
rect 469372 698468 469386 698470
rect 468822 698448 469386 698468
rect 455236 697332 455288 697338
rect 455236 697274 455288 697280
rect 450096 695978 450478 695994
rect 455248 695980 455276 697274
rect 464712 697264 464764 697270
rect 464712 697206 464764 697212
rect 464724 695980 464752 697206
rect 474200 695980 474228 698770
rect 516782 698728 516838 698737
rect 488356 698692 488408 698698
rect 516782 698663 516838 698672
rect 488356 698634 488408 698640
rect 488368 695980 488396 698634
rect 504822 698524 505386 698544
rect 504822 698522 504836 698524
rect 504892 698522 504916 698524
rect 504972 698522 504996 698524
rect 505052 698522 505076 698524
rect 505132 698522 505156 698524
rect 505212 698522 505236 698524
rect 505292 698522 505316 698524
rect 505372 698522 505386 698524
rect 505066 698470 505076 698522
rect 505132 698470 505142 698522
rect 504822 698468 504836 698470
rect 504892 698468 504916 698470
rect 504972 698468 504996 698470
rect 505052 698468 505076 698470
rect 505132 698468 505156 698470
rect 505212 698468 505236 698470
rect 505292 698468 505316 698470
rect 505372 698468 505386 698470
rect 504822 698448 505386 698468
rect 493048 697196 493100 697202
rect 493048 697138 493100 697144
rect 493060 695980 493088 697138
rect 516796 695980 516824 698663
rect 526272 695980 526300 698799
rect 530964 695980 530992 699207
rect 558822 699068 559386 699088
rect 558822 699066 558836 699068
rect 558892 699066 558916 699068
rect 558972 699066 558996 699068
rect 559052 699066 559076 699068
rect 559132 699066 559156 699068
rect 559212 699066 559236 699068
rect 559292 699066 559316 699068
rect 559372 699066 559386 699068
rect 559066 699014 559076 699066
rect 559132 699014 559142 699066
rect 558822 699012 558836 699014
rect 558892 699012 558916 699014
rect 558972 699012 558996 699014
rect 559052 699012 559076 699014
rect 559132 699012 559156 699014
rect 559212 699012 559236 699014
rect 559292 699012 559316 699014
rect 559372 699012 559386 699014
rect 558822 698992 559386 699012
rect 576584 698964 576636 698970
rect 576584 698906 576636 698912
rect 576400 698624 576452 698630
rect 576400 698566 576452 698572
rect 540822 698524 541386 698544
rect 540822 698522 540836 698524
rect 540892 698522 540916 698524
rect 540972 698522 540996 698524
rect 541052 698522 541076 698524
rect 541132 698522 541156 698524
rect 541212 698522 541236 698524
rect 541292 698522 541316 698524
rect 541372 698522 541386 698524
rect 541066 698470 541076 698522
rect 541132 698470 541142 698522
rect 540822 698468 540836 698470
rect 540892 698468 540916 698470
rect 540972 698468 540996 698470
rect 541052 698468 541076 698470
rect 541132 698468 541156 698470
rect 541212 698468 541236 698470
rect 541292 698468 541316 698470
rect 541372 698468 541386 698470
rect 540822 698448 541386 698468
rect 576308 698352 576360 698358
rect 576308 698294 576360 698300
rect 574560 698148 574612 698154
rect 574560 698090 574612 698096
rect 535644 697128 535696 697134
rect 535644 697070 535696 697076
rect 540426 697096 540482 697105
rect 535656 695980 535684 697070
rect 540426 697031 540482 697040
rect 540440 695980 540468 697031
rect 450084 695972 450478 695978
rect 450136 695966 450478 695972
rect 450084 695914 450136 695920
rect 459652 695904 459704 695910
rect 509514 695872 509570 695881
rect 459704 695852 459954 695858
rect 459652 695846 459954 695852
rect 459664 695830 459954 695846
rect 478800 695842 478906 695858
rect 478788 695836 478906 695842
rect 478840 695830 478906 695836
rect 509514 695807 509570 695816
rect 518070 695872 518126 695881
rect 518070 695807 518126 695816
rect 478788 695778 478840 695784
rect 483388 695768 483440 695774
rect 502340 695768 502392 695774
rect 483440 695716 483690 695722
rect 483388 695710 483690 695716
rect 502392 695728 502564 695756
rect 502340 695710 502392 695716
rect 483400 695694 483690 695710
rect 502536 695708 502564 695728
rect 506940 695632 506992 695638
rect 509528 695609 509556 695807
rect 518084 695609 518112 695807
rect 545026 695736 545082 695745
rect 545082 695694 545146 695722
rect 545026 695671 545082 695680
rect 509514 695600 509570 695609
rect 506992 695580 507334 695586
rect 506940 695574 507334 695580
rect 506952 695558 507334 695574
rect 509514 695535 509570 695544
rect 518070 695600 518126 695609
rect 518070 695535 518126 695544
rect 355508 695496 355560 695502
rect 355560 695444 355810 695450
rect 355508 695438 355810 695444
rect 355520 695422 355810 695438
rect 369964 695434 370070 695450
rect 369952 695428 370070 695434
rect 370004 695422 370070 695428
rect 369952 695370 370004 695376
rect 383844 695360 383896 695366
rect 185426 695298 185808 695314
rect 199686 695298 199976 695314
rect 426532 695360 426584 695366
rect 383896 695308 384238 695314
rect 383844 695302 384238 695308
rect 440700 695360 440752 695366
rect 426584 695308 426834 695314
rect 426532 695302 426834 695308
rect 469220 695360 469272 695366
rect 440752 695308 441002 695314
rect 440700 695302 441002 695308
rect 497556 695360 497608 695366
rect 469272 695308 469430 695314
rect 469220 695302 469430 695308
rect 511908 695360 511960 695366
rect 497608 695308 497858 695314
rect 497556 695302 497858 695308
rect 521382 695328 521438 695337
rect 511960 695308 512026 695314
rect 511908 695302 512026 695308
rect 176198 695263 176254 695272
rect 179328 695292 179380 695298
rect 157432 695234 157484 695240
rect 185426 695292 185820 695298
rect 185426 695286 185768 695292
rect 179328 695234 179380 695240
rect 199686 695292 199988 695298
rect 199686 695286 199936 695292
rect 185768 695234 185820 695240
rect 383856 695286 384238 695302
rect 426544 695286 426834 695302
rect 440712 695286 441002 695302
rect 469232 695286 469430 695302
rect 497568 695286 497858 695302
rect 511920 695286 512026 695302
rect 521438 695286 521502 695314
rect 521382 695263 521438 695272
rect 199936 695234 199988 695240
rect 569866 694104 569922 694113
rect 569866 694039 569922 694048
rect 569880 693705 569908 694039
rect 569866 693696 569922 693705
rect 569866 693631 569922 693640
rect 574572 674937 574600 698090
rect 574652 697944 574704 697950
rect 574652 697886 574704 697892
rect 574558 674928 574614 674937
rect 574558 674863 574614 674872
rect 574664 628017 574692 697886
rect 575388 697740 575440 697746
rect 575388 697682 575440 697688
rect 574928 697060 574980 697066
rect 574928 697002 574980 697008
rect 574742 696960 574798 696969
rect 574742 696895 574798 696904
rect 574650 628008 574706 628017
rect 574650 627943 574706 627952
rect 7932 165708 7984 165714
rect 7932 165650 7984 165656
rect 7840 136400 7892 136406
rect 7840 136342 7892 136348
rect 7748 122120 7800 122126
rect 7748 122062 7800 122068
rect 7656 79892 7708 79898
rect 7656 79834 7708 79840
rect 7564 35828 7616 35834
rect 7564 35770 7616 35776
rect 574756 17762 574784 696895
rect 574834 694240 574890 694249
rect 574834 694175 574890 694184
rect 574848 41154 574876 694175
rect 574940 111790 574968 697002
rect 575296 694544 575348 694550
rect 575296 694486 575348 694492
rect 575204 694408 575256 694414
rect 575204 694350 575256 694356
rect 575112 694340 575164 694346
rect 575112 694282 575164 694288
rect 575020 694204 575072 694210
rect 575020 694146 575072 694152
rect 575032 182170 575060 694146
rect 575124 205562 575152 694282
rect 575216 252550 575244 694350
rect 575308 299470 575336 694486
rect 575400 580922 575428 697682
rect 576216 696992 576268 696998
rect 576216 696934 576268 696940
rect 576122 695600 576178 695609
rect 576122 695535 576178 695544
rect 576032 695088 576084 695094
rect 576032 695030 576084 695036
rect 575478 674928 575534 674937
rect 575478 674863 575534 674872
rect 575492 674830 575520 674863
rect 575480 674824 575532 674830
rect 575480 674766 575532 674772
rect 575478 628008 575534 628017
rect 575478 627943 575534 627952
rect 575492 627910 575520 627943
rect 575480 627904 575532 627910
rect 575480 627846 575532 627852
rect 575388 580916 575440 580922
rect 575388 580858 575440 580864
rect 576044 510610 576072 695030
rect 576032 510604 576084 510610
rect 576032 510546 576084 510552
rect 575296 299464 575348 299470
rect 575296 299406 575348 299412
rect 575204 252544 575256 252550
rect 575204 252486 575256 252492
rect 575112 205556 575164 205562
rect 575112 205498 575164 205504
rect 575020 182164 575072 182170
rect 575020 182106 575072 182112
rect 574928 111784 574980 111790
rect 574928 111726 574980 111732
rect 575020 41268 575072 41274
rect 575020 41210 575072 41216
rect 575032 41154 575060 41210
rect 574848 41126 575060 41154
rect 576136 30326 576164 695535
rect 576228 64870 576256 696934
rect 576320 171086 576348 698294
rect 576412 264858 576440 698566
rect 576492 694680 576544 694686
rect 576492 694622 576544 694628
rect 576504 346390 576532 694622
rect 576596 416634 576624 698906
rect 577688 698896 577740 698902
rect 577688 698838 577740 698844
rect 577596 698760 577648 698766
rect 577596 698702 577648 698708
rect 576822 698524 577386 698544
rect 576822 698522 576836 698524
rect 576892 698522 576916 698524
rect 576972 698522 576996 698524
rect 577052 698522 577076 698524
rect 577132 698522 577156 698524
rect 577212 698522 577236 698524
rect 577292 698522 577316 698524
rect 577372 698522 577386 698524
rect 577066 698470 577076 698522
rect 577132 698470 577142 698522
rect 576822 698468 576836 698470
rect 576892 698468 576916 698470
rect 576972 698468 576996 698470
rect 577052 698468 577076 698470
rect 577132 698468 577156 698470
rect 577212 698468 577236 698470
rect 577292 698468 577316 698470
rect 577372 698468 577386 698470
rect 576822 698448 577386 698468
rect 576768 697468 576820 697474
rect 576768 697410 576820 697416
rect 576676 694884 576728 694890
rect 576676 694826 576728 694832
rect 576688 440230 576716 694826
rect 576780 487150 576808 697410
rect 577504 695564 577556 695570
rect 577504 695506 577556 695512
rect 577412 695292 577464 695298
rect 577412 695234 577464 695240
rect 577424 651370 577452 695234
rect 577412 651364 577464 651370
rect 577412 651306 577464 651312
rect 576768 487144 576820 487150
rect 576768 487086 576820 487092
rect 576676 440224 576728 440230
rect 576676 440166 576728 440172
rect 576584 416628 576636 416634
rect 576584 416570 576636 416576
rect 576492 346384 576544 346390
rect 576492 346326 576544 346332
rect 576400 264852 576452 264858
rect 576400 264794 576452 264800
rect 576308 171080 576360 171086
rect 576308 171022 576360 171028
rect 577516 158710 577544 695506
rect 577608 311846 577636 698702
rect 577700 358766 577728 698838
rect 577780 696040 577832 696046
rect 577780 695982 577832 695988
rect 577792 463690 577820 695982
rect 577884 499118 577912 699246
rect 579160 699168 579212 699174
rect 579160 699110 579212 699116
rect 578884 698420 578936 698426
rect 578884 698362 578936 698368
rect 577964 697604 578016 697610
rect 577964 697546 578016 697552
rect 577976 534070 578004 697546
rect 578792 696652 578844 696658
rect 578792 696594 578844 696600
rect 578148 695360 578200 695366
rect 578148 695302 578200 695308
rect 578056 695156 578108 695162
rect 578056 695098 578108 695104
rect 578068 557394 578096 695098
rect 578160 604314 578188 695302
rect 578804 687206 578832 696594
rect 578792 687200 578844 687206
rect 578792 687142 578844 687148
rect 578148 604308 578200 604314
rect 578148 604250 578200 604256
rect 578056 557388 578108 557394
rect 578056 557330 578108 557336
rect 577964 534064 578016 534070
rect 577964 534006 578016 534012
rect 577872 499112 577924 499118
rect 577872 499054 577924 499060
rect 577780 463684 577832 463690
rect 577780 463626 577832 463632
rect 577688 358760 577740 358766
rect 577688 358702 577740 358708
rect 577596 311840 577648 311846
rect 577596 311782 577648 311788
rect 578896 217025 578924 698362
rect 579068 694816 579120 694822
rect 579068 694758 579120 694764
rect 578976 694612 579028 694618
rect 578976 694554 579028 694560
rect 578988 322697 579016 694554
rect 579080 393009 579108 694758
rect 579172 404841 579200 699110
rect 580632 698216 580684 698222
rect 580632 698158 580684 698164
rect 579620 698080 579672 698086
rect 579618 698048 579620 698057
rect 579672 698048 579674 698057
rect 579618 697983 579674 697992
rect 579528 696516 579580 696522
rect 579528 696458 579580 696464
rect 579436 696176 579488 696182
rect 579436 696118 579488 696124
rect 579252 696108 579304 696114
rect 579252 696050 579304 696056
rect 579264 451761 579292 696050
rect 579342 694104 579398 694113
rect 579342 694039 579398 694048
rect 579356 545601 579384 694039
rect 579448 592521 579476 696118
rect 579540 639441 579568 696458
rect 580448 696448 580500 696454
rect 580448 696390 580500 696396
rect 580264 696244 580316 696250
rect 580264 696186 580316 696192
rect 579804 674824 579856 674830
rect 579804 674766 579856 674772
rect 579816 674665 579844 674766
rect 579802 674656 579858 674665
rect 579802 674591 579858 674600
rect 579620 651364 579672 651370
rect 579620 651306 579672 651312
rect 579632 651137 579660 651306
rect 579618 651128 579674 651137
rect 579618 651063 579674 651072
rect 579526 639432 579582 639441
rect 579526 639367 579582 639376
rect 579804 627904 579856 627910
rect 579804 627846 579856 627852
rect 579816 627745 579844 627846
rect 579802 627736 579858 627745
rect 579802 627671 579858 627680
rect 579620 604308 579672 604314
rect 579620 604250 579672 604256
rect 579632 604217 579660 604250
rect 579618 604208 579674 604217
rect 579618 604143 579674 604152
rect 579434 592512 579490 592521
rect 579434 592447 579490 592456
rect 580172 580916 580224 580922
rect 580172 580858 580224 580864
rect 580184 580825 580212 580858
rect 580170 580816 580226 580825
rect 580170 580751 580226 580760
rect 579620 557388 579672 557394
rect 579620 557330 579672 557336
rect 579632 557297 579660 557330
rect 579618 557288 579674 557297
rect 579618 557223 579674 557232
rect 579342 545592 579398 545601
rect 579342 545527 579398 545536
rect 579712 534064 579764 534070
rect 579712 534006 579764 534012
rect 579724 533905 579752 534006
rect 579710 533896 579766 533905
rect 579710 533831 579766 533840
rect 580172 510604 580224 510610
rect 580172 510546 580224 510552
rect 580184 510377 580212 510546
rect 580170 510368 580226 510377
rect 580170 510303 580226 510312
rect 580172 499112 580224 499118
rect 580172 499054 580224 499060
rect 580184 498681 580212 499054
rect 580170 498672 580226 498681
rect 580170 498607 580226 498616
rect 579988 487144 580040 487150
rect 579988 487086 580040 487092
rect 580000 486849 580028 487086
rect 579986 486840 580042 486849
rect 579986 486775 580042 486784
rect 579620 463684 579672 463690
rect 579620 463626 579672 463632
rect 579632 463457 579660 463626
rect 579618 463448 579674 463457
rect 579618 463383 579674 463392
rect 579250 451752 579306 451761
rect 579250 451687 579306 451696
rect 579988 440224 580040 440230
rect 579988 440166 580040 440172
rect 580000 439929 580028 440166
rect 579986 439920 580042 439929
rect 579986 439855 580042 439864
rect 580172 416628 580224 416634
rect 580172 416570 580224 416576
rect 580184 416537 580212 416570
rect 580170 416528 580226 416537
rect 580170 416463 580226 416472
rect 579158 404832 579214 404841
rect 579158 404767 579214 404776
rect 579066 393000 579122 393009
rect 579066 392935 579122 392944
rect 579988 346384 580040 346390
rect 579988 346326 580040 346332
rect 580000 346089 580028 346326
rect 579986 346080 580042 346089
rect 579986 346015 580042 346024
rect 578974 322688 579030 322697
rect 578974 322623 579030 322632
rect 579620 299464 579672 299470
rect 579620 299406 579672 299412
rect 579632 299169 579660 299406
rect 579618 299160 579674 299169
rect 579618 299095 579674 299104
rect 580172 264852 580224 264858
rect 580172 264794 580224 264800
rect 580184 263945 580212 264794
rect 580170 263936 580226 263945
rect 580170 263871 580226 263880
rect 580172 252544 580224 252550
rect 580172 252486 580224 252492
rect 580184 252249 580212 252486
rect 580170 252240 580226 252249
rect 580170 252175 580226 252184
rect 578882 217016 578938 217025
rect 578882 216951 578938 216960
rect 580172 205556 580224 205562
rect 580172 205498 580224 205504
rect 580184 205329 580212 205498
rect 580170 205320 580226 205329
rect 580170 205255 580226 205264
rect 580172 182164 580224 182170
rect 580172 182106 580224 182112
rect 580184 181937 580212 182106
rect 580170 181928 580226 181937
rect 580170 181863 580226 181872
rect 579620 171080 579672 171086
rect 579620 171022 579672 171028
rect 579632 170105 579660 171022
rect 579618 170096 579674 170105
rect 579618 170031 579674 170040
rect 577504 158704 577556 158710
rect 577504 158646 577556 158652
rect 579620 111784 579672 111790
rect 579620 111726 579672 111732
rect 579632 111489 579660 111726
rect 579618 111480 579674 111489
rect 579618 111415 579674 111424
rect 580276 76265 580304 696186
rect 580354 693832 580410 693841
rect 580354 693767 580410 693776
rect 580368 87961 580396 693767
rect 580460 123185 580488 696390
rect 580538 693968 580594 693977
rect 580538 693903 580594 693912
rect 580552 134881 580580 693903
rect 580644 228857 580672 698158
rect 580816 697672 580868 697678
rect 580816 697614 580868 697620
rect 580724 696584 580776 696590
rect 580724 696526 580776 696532
rect 580736 275777 580764 696526
rect 580828 369617 580856 697614
rect 580908 687200 580960 687206
rect 580908 687142 580960 687148
rect 580920 686361 580948 687142
rect 580906 686352 580962 686361
rect 580906 686287 580962 686296
rect 580814 369608 580870 369617
rect 580814 369543 580870 369552
rect 580816 358760 580868 358766
rect 580816 358702 580868 358708
rect 580828 357921 580856 358702
rect 580814 357912 580870 357921
rect 580814 357847 580870 357856
rect 580816 311840 580868 311846
rect 580816 311782 580868 311788
rect 580828 310865 580856 311782
rect 580814 310856 580870 310865
rect 580814 310791 580870 310800
rect 580722 275768 580778 275777
rect 580722 275703 580778 275712
rect 580630 228848 580686 228857
rect 580630 228783 580686 228792
rect 580632 158704 580684 158710
rect 580632 158646 580684 158652
rect 580644 158409 580672 158646
rect 580630 158400 580686 158409
rect 580630 158335 580686 158344
rect 580538 134872 580594 134881
rect 580538 134807 580594 134816
rect 580446 123176 580502 123185
rect 580446 123111 580502 123120
rect 580354 87952 580410 87961
rect 580354 87887 580410 87896
rect 580262 76256 580318 76265
rect 580262 76191 580318 76200
rect 576216 64864 576268 64870
rect 576216 64806 576268 64812
rect 579804 64864 579856 64870
rect 579804 64806 579856 64812
rect 579816 64569 579844 64806
rect 579802 64560 579858 64569
rect 579802 64495 579858 64504
rect 580172 41268 580224 41274
rect 580172 41210 580224 41216
rect 580184 41041 580212 41210
rect 580170 41032 580226 41041
rect 580170 40967 580226 40976
rect 576124 30320 576176 30326
rect 576124 30262 576176 30268
rect 580172 30320 580224 30326
rect 580172 30262 580224 30268
rect 580184 29345 580212 30262
rect 580170 29336 580226 29345
rect 580170 29271 580226 29280
rect 575020 17876 575072 17882
rect 575020 17818 575072 17824
rect 580172 17876 580224 17882
rect 580172 17818 580224 17824
rect 575032 17762 575060 17818
rect 574756 17734 575060 17762
rect 580184 17649 580212 17818
rect 580170 17640 580226 17649
rect 580170 17575 580226 17584
rect 3148 7200 3200 7206
rect 3146 7168 3148 7177
rect 6184 7200 6236 7206
rect 3200 7168 3202 7177
rect 6184 7142 6236 7148
rect 3146 7103 3202 7112
rect 5540 6180 5592 6186
rect 5540 6122 5592 6128
rect 572 4072 624 4078
rect 572 4014 624 4020
rect 584 480 612 4014
rect 5264 3732 5316 3738
rect 5264 3674 5316 3680
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 1676 3052 1728 3058
rect 1676 2994 1728 3000
rect 1688 480 1716 2994
rect 2872 2916 2924 2922
rect 2872 2858 2924 2864
rect 2884 480 2912 2858
rect 4080 480 4108 3470
rect 5276 480 5304 3674
rect 5552 2922 5580 6122
rect 8588 4078 8616 8092
rect 9692 5624 9720 8092
rect 10796 6186 10824 8092
rect 10784 6180 10836 6186
rect 10784 6122 10836 6128
rect 9600 5596 9720 5624
rect 8576 4072 8628 4078
rect 8576 4014 8628 4020
rect 6460 3664 6512 3670
rect 6460 3606 6512 3612
rect 5540 2916 5592 2922
rect 5540 2858 5592 2864
rect 6472 480 6500 3606
rect 7656 3460 7708 3466
rect 7656 3402 7708 3408
rect 7668 480 7696 3402
rect 9600 3058 9628 5596
rect 11244 4004 11296 4010
rect 11244 3946 11296 3952
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 8852 2984 8904 2990
rect 8852 2926 8904 2932
rect 8864 480 8892 2926
rect 10048 2916 10100 2922
rect 10048 2858 10100 2864
rect 10060 480 10088 2858
rect 11256 480 11284 3946
rect 11992 3534 12020 8092
rect 12452 8078 13110 8106
rect 13832 8078 14306 8106
rect 12452 5794 12480 8078
rect 12360 5766 12480 5794
rect 13832 5778 13860 8078
rect 12532 5772 12584 5778
rect 12360 3738 12388 5766
rect 12532 5714 12584 5720
rect 13820 5772 13872 5778
rect 13820 5714 13872 5720
rect 12440 5704 12492 5710
rect 12440 5646 12492 5652
rect 12348 3732 12400 3738
rect 12348 3674 12400 3680
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 12452 3466 12480 5646
rect 12544 3670 12572 5714
rect 15396 5710 15424 8092
rect 15384 5704 15436 5710
rect 15384 5646 15436 5652
rect 16592 5642 16620 8092
rect 17592 6180 17644 6186
rect 17592 6122 17644 6128
rect 13820 5636 13872 5642
rect 13820 5578 13872 5584
rect 16580 5636 16632 5642
rect 16580 5578 16632 5584
rect 12532 3664 12584 3670
rect 12532 3606 12584 3612
rect 12440 3460 12492 3466
rect 12440 3402 12492 3408
rect 12440 3120 12492 3126
rect 12440 3062 12492 3068
rect 12452 480 12480 3062
rect 13832 2990 13860 5578
rect 15200 5568 15252 5574
rect 15200 5510 15252 5516
rect 14832 3936 14884 3942
rect 14832 3878 14884 3884
rect 13820 2984 13872 2990
rect 13820 2926 13872 2932
rect 13636 2848 13688 2854
rect 13636 2790 13688 2796
rect 13648 480 13676 2790
rect 14844 480 14872 3878
rect 15212 2922 15240 5510
rect 17604 4010 17632 6122
rect 17696 5574 17724 8092
rect 18892 6186 18920 8092
rect 18880 6180 18932 6186
rect 18880 6122 18932 6128
rect 18822 6012 19386 6032
rect 18822 6010 18836 6012
rect 18892 6010 18916 6012
rect 18972 6010 18996 6012
rect 19052 6010 19076 6012
rect 19132 6010 19156 6012
rect 19212 6010 19236 6012
rect 19292 6010 19316 6012
rect 19372 6010 19386 6012
rect 19066 5958 19076 6010
rect 19132 5958 19142 6010
rect 18822 5956 18836 5958
rect 18892 5956 18916 5958
rect 18972 5956 18996 5958
rect 19052 5956 19076 5958
rect 19132 5956 19156 5958
rect 19212 5956 19236 5958
rect 19292 5956 19316 5958
rect 19372 5956 19386 5958
rect 18822 5936 19386 5956
rect 18696 5704 18748 5710
rect 18696 5646 18748 5652
rect 17684 5568 17736 5574
rect 17684 5510 17736 5516
rect 18328 5568 18380 5574
rect 18328 5510 18380 5516
rect 17592 4004 17644 4010
rect 17592 3946 17644 3952
rect 16028 3664 16080 3670
rect 16028 3606 16080 3612
rect 15200 2916 15252 2922
rect 15200 2858 15252 2864
rect 16040 480 16068 3606
rect 17224 3528 17276 3534
rect 17224 3470 17276 3476
rect 17236 480 17264 3470
rect 18340 3126 18368 5510
rect 18328 3120 18380 3126
rect 18328 3062 18380 3068
rect 18328 2984 18380 2990
rect 18328 2926 18380 2932
rect 18340 480 18368 2926
rect 18708 2854 18736 5646
rect 19432 5636 19484 5642
rect 19432 5578 19484 5584
rect 18822 4924 19386 4944
rect 18822 4922 18836 4924
rect 18892 4922 18916 4924
rect 18972 4922 18996 4924
rect 19052 4922 19076 4924
rect 19132 4922 19156 4924
rect 19212 4922 19236 4924
rect 19292 4922 19316 4924
rect 19372 4922 19386 4924
rect 19066 4870 19076 4922
rect 19132 4870 19142 4922
rect 18822 4868 18836 4870
rect 18892 4868 18916 4870
rect 18972 4868 18996 4870
rect 19052 4868 19076 4870
rect 19132 4868 19156 4870
rect 19212 4868 19236 4870
rect 19292 4868 19316 4870
rect 19372 4868 19386 4870
rect 18822 4848 19386 4868
rect 19444 3942 19472 5578
rect 19996 5574 20024 8092
rect 21100 5710 21128 8092
rect 21088 5704 21140 5710
rect 21088 5646 21140 5652
rect 22100 5704 22152 5710
rect 22100 5646 22152 5652
rect 19984 5568 20036 5574
rect 19984 5510 20036 5516
rect 20812 5568 20864 5574
rect 20812 5510 20864 5516
rect 20720 4072 20772 4078
rect 20720 4014 20772 4020
rect 19432 3936 19484 3942
rect 19432 3878 19484 3884
rect 18822 3836 19386 3856
rect 18822 3834 18836 3836
rect 18892 3834 18916 3836
rect 18972 3834 18996 3836
rect 19052 3834 19076 3836
rect 19132 3834 19156 3836
rect 19212 3834 19236 3836
rect 19292 3834 19316 3836
rect 19372 3834 19386 3836
rect 19066 3782 19076 3834
rect 19132 3782 19142 3834
rect 18822 3780 18836 3782
rect 18892 3780 18916 3782
rect 18972 3780 18996 3782
rect 19052 3780 19076 3782
rect 19132 3780 19156 3782
rect 19212 3780 19236 3782
rect 19292 3780 19316 3782
rect 19372 3780 19386 3782
rect 18822 3760 19386 3780
rect 19524 3052 19576 3058
rect 19524 2994 19576 3000
rect 18696 2848 18748 2854
rect 18696 2790 18748 2796
rect 18822 2748 19386 2768
rect 18822 2746 18836 2748
rect 18892 2746 18916 2748
rect 18972 2746 18996 2748
rect 19052 2746 19076 2748
rect 19132 2746 19156 2748
rect 19212 2746 19236 2748
rect 19292 2746 19316 2748
rect 19372 2746 19386 2748
rect 19066 2694 19076 2746
rect 19132 2694 19142 2746
rect 18822 2692 18836 2694
rect 18892 2692 18916 2694
rect 18972 2692 18996 2694
rect 19052 2692 19076 2694
rect 19132 2692 19156 2694
rect 19212 2692 19236 2694
rect 19292 2692 19316 2694
rect 19372 2692 19386 2694
rect 18822 2672 19386 2692
rect 19536 480 19564 2994
rect 20732 480 20760 4014
rect 20824 3670 20852 5510
rect 20812 3664 20864 3670
rect 20812 3606 20864 3612
rect 22112 3534 22140 5646
rect 22296 5642 22324 8092
rect 22284 5636 22336 5642
rect 22284 5578 22336 5584
rect 23400 5574 23428 8092
rect 24596 5710 24624 8092
rect 24584 5704 24636 5710
rect 24584 5646 24636 5652
rect 25700 5574 25728 8092
rect 26252 8078 26910 8106
rect 27632 8078 28014 8106
rect 26252 6338 26280 8078
rect 26160 6310 26280 6338
rect 23388 5568 23440 5574
rect 23388 5510 23440 5516
rect 23480 5568 23532 5574
rect 23480 5510 23532 5516
rect 25688 5568 25740 5574
rect 25688 5510 25740 5516
rect 22100 3528 22152 3534
rect 22100 3470 22152 3476
rect 23112 3188 23164 3194
rect 23112 3130 23164 3136
rect 21916 2916 21968 2922
rect 21916 2858 21968 2864
rect 21928 480 21956 2858
rect 23124 480 23152 3130
rect 23492 2990 23520 5510
rect 25504 3936 25556 3942
rect 25504 3878 25556 3884
rect 24308 3528 24360 3534
rect 24308 3470 24360 3476
rect 23480 2984 23532 2990
rect 23480 2926 23532 2932
rect 24320 480 24348 3470
rect 25516 480 25544 3878
rect 26160 3058 26188 6310
rect 27632 5658 27660 8078
rect 27540 5630 27660 5658
rect 29000 5704 29052 5710
rect 29000 5646 29052 5652
rect 28264 5636 28316 5642
rect 26608 5568 26660 5574
rect 26608 5510 26660 5516
rect 26148 3052 26200 3058
rect 26148 2994 26200 3000
rect 26620 2922 26648 5510
rect 27540 4078 27568 5630
rect 28264 5578 28316 5584
rect 27528 4072 27580 4078
rect 27528 4014 27580 4020
rect 27896 3596 27948 3602
rect 27896 3538 27948 3544
rect 26700 3460 26752 3466
rect 26700 3402 26752 3408
rect 26608 2916 26660 2922
rect 26608 2858 26660 2864
rect 26712 480 26740 3402
rect 27908 480 27936 3538
rect 28276 3194 28304 5578
rect 29012 3534 29040 5646
rect 29196 5574 29224 8092
rect 30300 5642 30328 8092
rect 31404 5710 31432 8092
rect 31392 5704 31444 5710
rect 31392 5646 31444 5652
rect 30288 5636 30340 5642
rect 30288 5578 30340 5584
rect 31760 5636 31812 5642
rect 31760 5578 31812 5584
rect 29184 5568 29236 5574
rect 29184 5510 29236 5516
rect 30380 5568 30432 5574
rect 30380 5510 30432 5516
rect 30392 3942 30420 5510
rect 31484 4072 31536 4078
rect 31484 4014 31536 4020
rect 30380 3936 30432 3942
rect 30380 3878 30432 3884
rect 29000 3528 29052 3534
rect 29000 3470 29052 3476
rect 28264 3188 28316 3194
rect 28264 3130 28316 3136
rect 29092 2916 29144 2922
rect 29092 2858 29144 2864
rect 29104 480 29132 2858
rect 30288 2848 30340 2854
rect 30288 2790 30340 2796
rect 30300 480 30328 2790
rect 31496 480 31524 4014
rect 31772 3466 31800 5578
rect 32600 5574 32628 8092
rect 33152 8078 33718 8106
rect 34532 8078 34914 8106
rect 35912 8078 36018 8106
rect 33152 5642 33180 8078
rect 34532 5794 34560 8078
rect 34348 5766 34560 5794
rect 33140 5636 33192 5642
rect 33140 5578 33192 5584
rect 32588 5568 32640 5574
rect 32588 5510 32640 5516
rect 34348 3602 34376 5766
rect 35912 5658 35940 8078
rect 34520 5636 34572 5642
rect 34520 5578 34572 5584
rect 35820 5630 35940 5658
rect 37200 5642 37228 8092
rect 37188 5636 37240 5642
rect 34336 3596 34388 3602
rect 34336 3538 34388 3544
rect 31760 3460 31812 3466
rect 31760 3402 31812 3408
rect 33876 3460 33928 3466
rect 33876 3402 33928 3408
rect 32680 3120 32732 3126
rect 32680 3062 32732 3068
rect 32692 480 32720 3062
rect 33888 480 33916 3402
rect 34532 2854 34560 5578
rect 34980 3596 35032 3602
rect 34980 3538 35032 3544
rect 34520 2848 34572 2854
rect 34520 2790 34572 2796
rect 34992 480 35020 3538
rect 35820 2922 35848 5630
rect 37188 5578 37240 5584
rect 37648 5636 37700 5642
rect 37648 5578 37700 5584
rect 36728 5568 36780 5574
rect 36728 5510 36780 5516
rect 36740 4078 36768 5510
rect 36822 5468 37386 5488
rect 36822 5466 36836 5468
rect 36892 5466 36916 5468
rect 36972 5466 36996 5468
rect 37052 5466 37076 5468
rect 37132 5466 37156 5468
rect 37212 5466 37236 5468
rect 37292 5466 37316 5468
rect 37372 5466 37386 5468
rect 37066 5414 37076 5466
rect 37132 5414 37142 5466
rect 36822 5412 36836 5414
rect 36892 5412 36916 5414
rect 36972 5412 36996 5414
rect 37052 5412 37076 5414
rect 37132 5412 37156 5414
rect 37212 5412 37236 5414
rect 37292 5412 37316 5414
rect 37372 5412 37386 5414
rect 36822 5392 37386 5412
rect 36822 4380 37386 4400
rect 36822 4378 36836 4380
rect 36892 4378 36916 4380
rect 36972 4378 36996 4380
rect 37052 4378 37076 4380
rect 37132 4378 37156 4380
rect 37212 4378 37236 4380
rect 37292 4378 37316 4380
rect 37372 4378 37386 4380
rect 37066 4326 37076 4378
rect 37132 4326 37142 4378
rect 36822 4324 36836 4326
rect 36892 4324 36916 4326
rect 36972 4324 36996 4326
rect 37052 4324 37076 4326
rect 37132 4324 37156 4326
rect 37212 4324 37236 4326
rect 37292 4324 37316 4326
rect 37372 4324 37386 4326
rect 36822 4304 37386 4324
rect 36728 4072 36780 4078
rect 36728 4014 36780 4020
rect 36176 3664 36228 3670
rect 36176 3606 36228 3612
rect 35808 2916 35860 2922
rect 35808 2858 35860 2864
rect 36188 480 36216 3606
rect 37464 3528 37516 3534
rect 37464 3470 37516 3476
rect 36822 3292 37386 3312
rect 36822 3290 36836 3292
rect 36892 3290 36916 3292
rect 36972 3290 36996 3292
rect 37052 3290 37076 3292
rect 37132 3290 37156 3292
rect 37212 3290 37236 3292
rect 37292 3290 37316 3292
rect 37372 3290 37386 3292
rect 37066 3238 37076 3290
rect 37132 3238 37142 3290
rect 36822 3236 36836 3238
rect 36892 3236 36916 3238
rect 36972 3236 36996 3238
rect 37052 3236 37076 3238
rect 37132 3236 37156 3238
rect 37212 3236 37236 3238
rect 37292 3236 37316 3238
rect 37372 3236 37386 3238
rect 36822 3216 37386 3236
rect 36822 2204 37386 2224
rect 36822 2202 36836 2204
rect 36892 2202 36916 2204
rect 36972 2202 36996 2204
rect 37052 2202 37076 2204
rect 37132 2202 37156 2204
rect 37212 2202 37236 2204
rect 37292 2202 37316 2204
rect 37372 2202 37386 2204
rect 37066 2150 37076 2202
rect 37132 2150 37142 2202
rect 36822 2148 36836 2150
rect 36892 2148 36916 2150
rect 36972 2148 36996 2150
rect 37052 2148 37076 2150
rect 37132 2148 37156 2150
rect 37212 2148 37236 2150
rect 37292 2148 37316 2150
rect 37372 2148 37386 2150
rect 36822 2128 37386 2148
rect 37476 1986 37504 3470
rect 37660 3126 37688 5578
rect 38304 5574 38332 8092
rect 39500 5642 39528 8092
rect 40052 8078 40618 8106
rect 41432 8078 41722 8106
rect 42812 8078 42918 8106
rect 40052 5658 40080 8078
rect 39488 5636 39540 5642
rect 39488 5578 39540 5584
rect 39868 5630 40080 5658
rect 38292 5568 38344 5574
rect 38292 5510 38344 5516
rect 39868 3466 39896 5630
rect 41432 5574 41460 8078
rect 42812 5658 42840 8078
rect 42628 5630 42840 5658
rect 40040 5568 40092 5574
rect 40040 5510 40092 5516
rect 41420 5568 41472 5574
rect 41420 5510 41472 5516
rect 40052 3602 40080 5510
rect 40960 4072 41012 4078
rect 40960 4014 41012 4020
rect 40040 3596 40092 3602
rect 40040 3538 40092 3544
rect 39856 3460 39908 3466
rect 39856 3402 39908 3408
rect 38568 3392 38620 3398
rect 38568 3334 38620 3340
rect 37648 3120 37700 3126
rect 37648 3062 37700 3068
rect 37384 1958 37504 1986
rect 37384 480 37412 1958
rect 38580 480 38608 3334
rect 39764 2848 39816 2854
rect 39764 2790 39816 2796
rect 39776 480 39804 2790
rect 40972 480 41000 4014
rect 42628 3670 42656 5630
rect 42800 5568 42852 5574
rect 42800 5510 42852 5516
rect 42616 3664 42668 3670
rect 42616 3606 42668 3612
rect 42812 3398 42840 5510
rect 43352 3664 43404 3670
rect 43352 3606 43404 3612
rect 42800 3392 42852 3398
rect 42800 3334 42852 3340
rect 42156 3120 42208 3126
rect 42156 3062 42208 3068
rect 42168 480 42196 3062
rect 43364 480 43392 3606
rect 44008 3534 44036 8092
rect 44180 5636 44232 5642
rect 44180 5578 44232 5584
rect 43996 3528 44048 3534
rect 43996 3470 44048 3476
rect 44192 2854 44220 5578
rect 45204 5574 45232 8092
rect 46308 5642 46336 8092
rect 46952 8078 47518 8106
rect 46296 5636 46348 5642
rect 46296 5578 46348 5584
rect 45192 5568 45244 5574
rect 46952 5556 46980 8078
rect 48608 5658 48636 8092
rect 45192 5510 45244 5516
rect 46860 5528 46980 5556
rect 48240 5630 48636 5658
rect 49712 8078 49818 8106
rect 46860 4078 46888 5528
rect 46848 4072 46900 4078
rect 46848 4014 46900 4020
rect 44548 3732 44600 3738
rect 44548 3674 44600 3680
rect 44180 2848 44232 2854
rect 44180 2790 44232 2796
rect 44560 480 44588 3674
rect 46940 3528 46992 3534
rect 46940 3470 46992 3476
rect 45744 3188 45796 3194
rect 45744 3130 45796 3136
rect 45756 480 45784 3130
rect 46952 480 46980 3470
rect 48136 3460 48188 3466
rect 48136 3402 48188 3408
rect 48148 480 48176 3402
rect 48240 3126 48268 5630
rect 49712 5556 49740 8078
rect 49620 5528 49740 5556
rect 49620 3670 49648 5528
rect 50528 4072 50580 4078
rect 50528 4014 50580 4020
rect 49608 3664 49660 3670
rect 49608 3606 49660 3612
rect 48228 3120 48280 3126
rect 48228 3062 48280 3068
rect 49332 2848 49384 2854
rect 49332 2790 49384 2796
rect 49344 480 49372 2790
rect 50540 480 50568 4014
rect 50908 3738 50936 8092
rect 51632 4140 51684 4146
rect 51632 4082 51684 4088
rect 50896 3732 50948 3738
rect 50896 3674 50948 3680
rect 51644 480 51672 4082
rect 52104 3194 52132 8092
rect 52828 3936 52880 3942
rect 52828 3878 52880 3884
rect 52092 3188 52144 3194
rect 52092 3130 52144 3136
rect 52840 480 52868 3878
rect 53208 3534 53236 8092
rect 53852 8078 54326 8106
rect 53852 5658 53880 8078
rect 54822 6012 55386 6032
rect 54822 6010 54836 6012
rect 54892 6010 54916 6012
rect 54972 6010 54996 6012
rect 55052 6010 55076 6012
rect 55132 6010 55156 6012
rect 55212 6010 55236 6012
rect 55292 6010 55316 6012
rect 55372 6010 55386 6012
rect 55066 5958 55076 6010
rect 55132 5958 55142 6010
rect 54822 5956 54836 5958
rect 54892 5956 54916 5958
rect 54972 5956 54996 5958
rect 55052 5956 55076 5958
rect 55132 5956 55156 5958
rect 55212 5956 55236 5958
rect 55292 5956 55316 5958
rect 55372 5956 55386 5958
rect 54822 5936 55386 5956
rect 53760 5630 53880 5658
rect 53196 3528 53248 3534
rect 53196 3470 53248 3476
rect 53760 3466 53788 5630
rect 55508 5574 55536 8092
rect 56612 5658 56640 8092
rect 56520 5630 56640 5658
rect 53840 5568 53892 5574
rect 53840 5510 53892 5516
rect 55496 5568 55548 5574
rect 55496 5510 55548 5516
rect 53748 3460 53800 3466
rect 53748 3402 53800 3408
rect 53852 2854 53880 5510
rect 54822 4924 55386 4944
rect 54822 4922 54836 4924
rect 54892 4922 54916 4924
rect 54972 4922 54996 4924
rect 55052 4922 55076 4924
rect 55132 4922 55156 4924
rect 55212 4922 55236 4924
rect 55292 4922 55316 4924
rect 55372 4922 55386 4924
rect 55066 4870 55076 4922
rect 55132 4870 55142 4922
rect 54822 4868 54836 4870
rect 54892 4868 54916 4870
rect 54972 4868 54996 4870
rect 55052 4868 55076 4870
rect 55132 4868 55156 4870
rect 55212 4868 55236 4870
rect 55292 4868 55316 4870
rect 55372 4868 55386 4870
rect 54822 4848 55386 4868
rect 56520 4078 56548 5630
rect 57808 4146 57836 8092
rect 57796 4140 57848 4146
rect 57796 4082 57848 4088
rect 56508 4072 56560 4078
rect 56508 4014 56560 4020
rect 55404 4004 55456 4010
rect 55404 3946 55456 3952
rect 54822 3836 55386 3856
rect 54822 3834 54836 3836
rect 54892 3834 54916 3836
rect 54972 3834 54996 3836
rect 55052 3834 55076 3836
rect 55132 3834 55156 3836
rect 55212 3834 55236 3836
rect 55292 3834 55316 3836
rect 55372 3834 55386 3836
rect 55066 3782 55076 3834
rect 55132 3782 55142 3834
rect 54822 3780 54836 3782
rect 54892 3780 54916 3782
rect 54972 3780 54996 3782
rect 55052 3780 55076 3782
rect 55132 3780 55156 3782
rect 55212 3780 55236 3782
rect 55292 3780 55316 3782
rect 55372 3780 55386 3782
rect 54822 3760 55386 3780
rect 54024 3664 54076 3670
rect 54024 3606 54076 3612
rect 53840 2848 53892 2854
rect 53840 2790 53892 2796
rect 54036 480 54064 3606
rect 54822 2748 55386 2768
rect 54822 2746 54836 2748
rect 54892 2746 54916 2748
rect 54972 2746 54996 2748
rect 55052 2746 55076 2748
rect 55132 2746 55156 2748
rect 55212 2746 55236 2748
rect 55292 2746 55316 2748
rect 55372 2746 55386 2748
rect 55066 2694 55076 2746
rect 55132 2694 55142 2746
rect 54822 2692 54836 2694
rect 54892 2692 54916 2694
rect 54972 2692 54996 2694
rect 55052 2692 55076 2694
rect 55132 2692 55156 2694
rect 55212 2692 55236 2694
rect 55292 2692 55316 2694
rect 55372 2692 55386 2694
rect 54822 2672 55386 2692
rect 55416 2530 55444 3946
rect 58912 3942 58940 8092
rect 60004 4072 60056 4078
rect 60004 4014 60056 4020
rect 58900 3936 58952 3942
rect 58900 3878 58952 3884
rect 57612 3596 57664 3602
rect 57612 3538 57664 3544
rect 56416 3528 56468 3534
rect 56416 3470 56468 3476
rect 55232 2502 55444 2530
rect 55232 480 55260 2502
rect 56428 480 56456 3470
rect 57624 480 57652 3538
rect 58808 3460 58860 3466
rect 58808 3402 58860 3408
rect 58820 480 58848 3402
rect 60016 480 60044 4014
rect 60108 3670 60136 8092
rect 61212 4010 61240 8092
rect 62132 8078 62422 8106
rect 62132 5658 62160 8078
rect 61948 5630 62160 5658
rect 61200 4004 61252 4010
rect 61200 3946 61252 3952
rect 61200 3732 61252 3738
rect 61200 3674 61252 3680
rect 60096 3664 60148 3670
rect 60096 3606 60148 3612
rect 61212 480 61240 3674
rect 61948 3534 61976 5630
rect 63512 5574 63540 8092
rect 62120 5568 62172 5574
rect 62120 5510 62172 5516
rect 63500 5568 63552 5574
rect 63500 5510 63552 5516
rect 62132 3602 62160 5510
rect 63592 3936 63644 3942
rect 63592 3878 63644 3884
rect 62120 3596 62172 3602
rect 62120 3538 62172 3544
rect 61936 3528 61988 3534
rect 61936 3470 61988 3476
rect 62396 3528 62448 3534
rect 62396 3470 62448 3476
rect 62408 480 62436 3470
rect 63604 480 63632 3878
rect 64616 3466 64644 8092
rect 65812 4078 65840 8092
rect 65800 4072 65852 4078
rect 65800 4014 65852 4020
rect 66916 3738 66944 8092
rect 66904 3732 66956 3738
rect 66904 3674 66956 3680
rect 67180 3596 67232 3602
rect 67180 3538 67232 3544
rect 64604 3460 64656 3466
rect 64604 3402 64656 3408
rect 64788 3460 64840 3466
rect 64788 3402 64840 3408
rect 64800 480 64828 3402
rect 65984 3188 66036 3194
rect 65984 3130 66036 3136
rect 65996 480 66024 3130
rect 67192 480 67220 3538
rect 68112 3534 68140 8092
rect 69216 3942 69244 8092
rect 70412 5658 70440 8092
rect 70228 5630 70440 5658
rect 69480 4072 69532 4078
rect 69480 4014 69532 4020
rect 69204 3936 69256 3942
rect 69204 3878 69256 3884
rect 68100 3528 68152 3534
rect 68100 3470 68152 3476
rect 68284 3528 68336 3534
rect 68284 3470 68336 3476
rect 68296 480 68324 3470
rect 69492 480 69520 4014
rect 70228 3466 70256 5630
rect 70676 4140 70728 4146
rect 70676 4082 70728 4088
rect 70216 3460 70268 3466
rect 70216 3402 70268 3408
rect 70688 480 70716 4082
rect 71516 3194 71544 8092
rect 72344 8078 72726 8106
rect 71872 5568 71924 5574
rect 71872 5510 71924 5516
rect 71504 3188 71556 3194
rect 71504 3130 71556 3136
rect 71884 480 71912 5510
rect 72344 3602 72372 8078
rect 72822 5468 73386 5488
rect 72822 5466 72836 5468
rect 72892 5466 72916 5468
rect 72972 5466 72996 5468
rect 73052 5466 73076 5468
rect 73132 5466 73156 5468
rect 73212 5466 73236 5468
rect 73292 5466 73316 5468
rect 73372 5466 73386 5468
rect 73066 5414 73076 5466
rect 73132 5414 73142 5466
rect 72822 5412 72836 5414
rect 72892 5412 72916 5414
rect 72972 5412 72996 5414
rect 73052 5412 73076 5414
rect 73132 5412 73156 5414
rect 73212 5412 73236 5414
rect 73292 5412 73316 5414
rect 73372 5412 73386 5414
rect 72822 5392 73386 5412
rect 72822 4380 73386 4400
rect 72822 4378 72836 4380
rect 72892 4378 72916 4380
rect 72972 4378 72996 4380
rect 73052 4378 73076 4380
rect 73132 4378 73156 4380
rect 73212 4378 73236 4380
rect 73292 4378 73316 4380
rect 73372 4378 73386 4380
rect 73066 4326 73076 4378
rect 73132 4326 73142 4378
rect 72822 4324 72836 4326
rect 72892 4324 72916 4326
rect 72972 4324 72996 4326
rect 73052 4324 73076 4326
rect 73132 4324 73156 4326
rect 73212 4324 73236 4326
rect 73292 4324 73316 4326
rect 73372 4324 73386 4326
rect 72822 4304 73386 4324
rect 72332 3596 72384 3602
rect 72332 3538 72384 3544
rect 72700 3596 72752 3602
rect 72700 3538 72752 3544
rect 72712 1850 72740 3538
rect 73816 3534 73844 8092
rect 74920 4078 74948 8092
rect 76116 4146 76144 8092
rect 77220 5574 77248 8092
rect 77208 5568 77260 5574
rect 77208 5510 77260 5516
rect 76104 4140 76156 4146
rect 76104 4082 76156 4088
rect 74908 4072 74960 4078
rect 74908 4014 74960 4020
rect 74264 4004 74316 4010
rect 74264 3946 74316 3952
rect 73804 3528 73856 3534
rect 73804 3470 73856 3476
rect 72822 3292 73386 3312
rect 72822 3290 72836 3292
rect 72892 3290 72916 3292
rect 72972 3290 72996 3292
rect 73052 3290 73076 3292
rect 73132 3290 73156 3292
rect 73212 3290 73236 3292
rect 73292 3290 73316 3292
rect 73372 3290 73386 3292
rect 73066 3238 73076 3290
rect 73132 3238 73142 3290
rect 72822 3236 72836 3238
rect 72892 3236 72916 3238
rect 72972 3236 72996 3238
rect 73052 3236 73076 3238
rect 73132 3236 73156 3238
rect 73212 3236 73236 3238
rect 73292 3236 73316 3238
rect 73372 3236 73386 3238
rect 72822 3216 73386 3236
rect 72822 2204 73386 2224
rect 72822 2202 72836 2204
rect 72892 2202 72916 2204
rect 72972 2202 72996 2204
rect 73052 2202 73076 2204
rect 73132 2202 73156 2204
rect 73212 2202 73236 2204
rect 73292 2202 73316 2204
rect 73372 2202 73386 2204
rect 73066 2150 73076 2202
rect 73132 2150 73142 2202
rect 72822 2148 72836 2150
rect 72892 2148 72916 2150
rect 72972 2148 72996 2150
rect 73052 2148 73076 2150
rect 73132 2148 73156 2150
rect 73212 2148 73236 2150
rect 73292 2148 73316 2150
rect 73372 2148 73386 2150
rect 72822 2128 73386 2148
rect 72712 1822 73108 1850
rect 73080 480 73108 1822
rect 74276 480 74304 3946
rect 78416 3602 78444 8092
rect 79048 5704 79100 5710
rect 79048 5646 79100 5652
rect 78404 3596 78456 3602
rect 78404 3538 78456 3544
rect 76656 3528 76708 3534
rect 76656 3470 76708 3476
rect 75460 3188 75512 3194
rect 75460 3130 75512 3136
rect 75472 480 75500 3130
rect 76668 480 76696 3470
rect 77852 3460 77904 3466
rect 77852 3402 77904 3408
rect 77864 480 77892 3402
rect 79060 480 79088 5646
rect 79520 4010 79548 8092
rect 80244 5568 80296 5574
rect 80244 5510 80296 5516
rect 79508 4004 79560 4010
rect 79508 3946 79560 3952
rect 80256 480 80284 5510
rect 80716 3194 80744 8092
rect 81440 5636 81492 5642
rect 81440 5578 81492 5584
rect 80704 3188 80756 3194
rect 80704 3130 80756 3136
rect 81452 480 81480 5578
rect 81820 3534 81848 8092
rect 82636 3596 82688 3602
rect 82636 3538 82688 3544
rect 81808 3528 81860 3534
rect 81808 3470 81860 3476
rect 82648 480 82676 3538
rect 83016 3466 83044 8092
rect 84120 5710 84148 8092
rect 84108 5704 84160 5710
rect 84108 5646 84160 5652
rect 85224 5574 85252 8092
rect 86132 6180 86184 6186
rect 86132 6122 86184 6128
rect 85212 5568 85264 5574
rect 85212 5510 85264 5516
rect 83832 3528 83884 3534
rect 83832 3470 83884 3476
rect 83004 3460 83056 3466
rect 83004 3402 83056 3408
rect 83844 480 83872 3470
rect 84936 2984 84988 2990
rect 84936 2926 84988 2932
rect 84948 480 84976 2926
rect 86144 480 86172 6122
rect 86420 5642 86448 8092
rect 86408 5636 86460 5642
rect 86408 5578 86460 5584
rect 87328 5636 87380 5642
rect 87328 5578 87380 5584
rect 87340 480 87368 5578
rect 87524 3602 87552 8092
rect 88524 6452 88576 6458
rect 88524 6394 88576 6400
rect 87512 3596 87564 3602
rect 87512 3538 87564 3544
rect 88536 480 88564 6394
rect 88720 3534 88748 8092
rect 89720 5568 89772 5574
rect 89720 5510 89772 5516
rect 88708 3528 88760 3534
rect 88708 3470 88760 3476
rect 89732 480 89760 5510
rect 89824 2990 89852 8092
rect 91020 6186 91048 8092
rect 91008 6180 91060 6186
rect 91008 6122 91060 6128
rect 90822 6012 91386 6032
rect 90822 6010 90836 6012
rect 90892 6010 90916 6012
rect 90972 6010 90996 6012
rect 91052 6010 91076 6012
rect 91132 6010 91156 6012
rect 91212 6010 91236 6012
rect 91292 6010 91316 6012
rect 91372 6010 91386 6012
rect 91066 5958 91076 6010
rect 91132 5958 91142 6010
rect 90822 5956 90836 5958
rect 90892 5956 90916 5958
rect 90972 5956 90996 5958
rect 91052 5956 91076 5958
rect 91132 5956 91156 5958
rect 91212 5956 91236 5958
rect 91292 5956 91316 5958
rect 91372 5956 91386 5958
rect 90822 5936 91386 5956
rect 92124 5642 92152 8092
rect 93320 6458 93348 8092
rect 93308 6452 93360 6458
rect 93308 6394 93360 6400
rect 93308 6316 93360 6322
rect 93308 6258 93360 6264
rect 92112 5636 92164 5642
rect 92112 5578 92164 5584
rect 90822 4924 91386 4944
rect 90822 4922 90836 4924
rect 90892 4922 90916 4924
rect 90972 4922 90996 4924
rect 91052 4922 91076 4924
rect 91132 4922 91156 4924
rect 91212 4922 91236 4924
rect 91292 4922 91316 4924
rect 91372 4922 91386 4924
rect 91066 4870 91076 4922
rect 91132 4870 91142 4922
rect 90822 4868 90836 4870
rect 90892 4868 90916 4870
rect 90972 4868 90996 4870
rect 91052 4868 91076 4870
rect 91132 4868 91156 4870
rect 91212 4868 91236 4870
rect 91292 4868 91316 4870
rect 91372 4868 91386 4870
rect 90822 4848 91386 4868
rect 90732 4072 90784 4078
rect 90732 4014 90784 4020
rect 89812 2984 89864 2990
rect 89812 2926 89864 2932
rect 90744 2122 90772 4014
rect 90822 3836 91386 3856
rect 90822 3834 90836 3836
rect 90892 3834 90916 3836
rect 90972 3834 90996 3836
rect 91052 3834 91076 3836
rect 91132 3834 91156 3836
rect 91212 3834 91236 3836
rect 91292 3834 91316 3836
rect 91372 3834 91386 3836
rect 91066 3782 91076 3834
rect 91132 3782 91142 3834
rect 90822 3780 90836 3782
rect 90892 3780 90916 3782
rect 90972 3780 90996 3782
rect 91052 3780 91076 3782
rect 91132 3780 91156 3782
rect 91212 3780 91236 3782
rect 91292 3780 91316 3782
rect 91372 3780 91386 3782
rect 90822 3760 91386 3780
rect 92112 3528 92164 3534
rect 92112 3470 92164 3476
rect 90822 2748 91386 2768
rect 90822 2746 90836 2748
rect 90892 2746 90916 2748
rect 90972 2746 90996 2748
rect 91052 2746 91076 2748
rect 91132 2746 91156 2748
rect 91212 2746 91236 2748
rect 91292 2746 91316 2748
rect 91372 2746 91386 2748
rect 91066 2694 91076 2746
rect 91132 2694 91142 2746
rect 90822 2692 90836 2694
rect 90892 2692 90916 2694
rect 90972 2692 90996 2694
rect 91052 2692 91076 2694
rect 91132 2692 91156 2694
rect 91212 2692 91236 2694
rect 91292 2692 91316 2694
rect 91372 2692 91386 2694
rect 90822 2672 91386 2692
rect 90744 2094 90956 2122
rect 90928 480 90956 2094
rect 92124 480 92152 3470
rect 93320 480 93348 6258
rect 94424 5574 94452 8092
rect 94504 5772 94556 5778
rect 94504 5714 94556 5720
rect 94412 5568 94464 5574
rect 94412 5510 94464 5516
rect 94516 480 94544 5714
rect 95620 4078 95648 8092
rect 95700 5568 95752 5574
rect 95700 5510 95752 5516
rect 95608 4072 95660 4078
rect 95608 4014 95660 4020
rect 95712 480 95740 5510
rect 96724 3534 96752 8092
rect 97828 6322 97856 8092
rect 97816 6316 97868 6322
rect 97816 6258 97868 6264
rect 99024 5778 99052 8092
rect 99012 5772 99064 5778
rect 99012 5714 99064 5720
rect 96896 5704 96948 5710
rect 96896 5646 96948 5652
rect 96712 3528 96764 3534
rect 96712 3470 96764 3476
rect 96908 480 96936 5646
rect 98092 5636 98144 5642
rect 98092 5578 98144 5584
rect 98104 480 98132 5578
rect 100128 5574 100156 8092
rect 101324 5710 101352 8092
rect 101312 5704 101364 5710
rect 101312 5646 101364 5652
rect 101588 5704 101640 5710
rect 101588 5646 101640 5652
rect 100116 5568 100168 5574
rect 100116 5510 100168 5516
rect 100484 5568 100536 5574
rect 100484 5510 100536 5516
rect 99288 4072 99340 4078
rect 99288 4014 99340 4020
rect 99300 480 99328 4014
rect 100496 480 100524 5510
rect 101600 480 101628 5646
rect 102428 5642 102456 8092
rect 102784 6452 102836 6458
rect 102784 6394 102836 6400
rect 102416 5636 102468 5642
rect 102416 5578 102468 5584
rect 102796 480 102824 6394
rect 103624 4078 103652 8092
rect 103980 5636 104032 5642
rect 103980 5578 104032 5584
rect 103612 4072 103664 4078
rect 103612 4014 103664 4020
rect 103992 480 104020 5578
rect 104728 5574 104756 8092
rect 105176 5840 105228 5846
rect 105176 5782 105228 5788
rect 104716 5568 104768 5574
rect 104716 5510 104768 5516
rect 105188 480 105216 5782
rect 105924 5710 105952 8092
rect 107028 6458 107056 8092
rect 107016 6452 107068 6458
rect 107016 6394 107068 6400
rect 107568 5772 107620 5778
rect 107568 5714 107620 5720
rect 105912 5704 105964 5710
rect 105912 5646 105964 5652
rect 106372 5568 106424 5574
rect 106372 5510 106424 5516
rect 106384 480 106412 5510
rect 107580 480 107608 5714
rect 108132 5642 108160 8092
rect 109328 5846 109356 8092
rect 109316 5840 109368 5846
rect 109316 5782 109368 5788
rect 109960 5704 110012 5710
rect 109960 5646 110012 5652
rect 108120 5636 108172 5642
rect 108120 5578 108172 5584
rect 108672 5636 108724 5642
rect 108672 5578 108724 5584
rect 108684 1986 108712 5578
rect 108822 5468 109386 5488
rect 108822 5466 108836 5468
rect 108892 5466 108916 5468
rect 108972 5466 108996 5468
rect 109052 5466 109076 5468
rect 109132 5466 109156 5468
rect 109212 5466 109236 5468
rect 109292 5466 109316 5468
rect 109372 5466 109386 5468
rect 109066 5414 109076 5466
rect 109132 5414 109142 5466
rect 108822 5412 108836 5414
rect 108892 5412 108916 5414
rect 108972 5412 108996 5414
rect 109052 5412 109076 5414
rect 109132 5412 109156 5414
rect 109212 5412 109236 5414
rect 109292 5412 109316 5414
rect 109372 5412 109386 5414
rect 108822 5392 109386 5412
rect 108822 4380 109386 4400
rect 108822 4378 108836 4380
rect 108892 4378 108916 4380
rect 108972 4378 108996 4380
rect 109052 4378 109076 4380
rect 109132 4378 109156 4380
rect 109212 4378 109236 4380
rect 109292 4378 109316 4380
rect 109372 4378 109386 4380
rect 109066 4326 109076 4378
rect 109132 4326 109142 4378
rect 108822 4324 108836 4326
rect 108892 4324 108916 4326
rect 108972 4324 108996 4326
rect 109052 4324 109076 4326
rect 109132 4324 109156 4326
rect 109212 4324 109236 4326
rect 109292 4324 109316 4326
rect 109372 4324 109386 4326
rect 108822 4304 109386 4324
rect 108822 3292 109386 3312
rect 108822 3290 108836 3292
rect 108892 3290 108916 3292
rect 108972 3290 108996 3292
rect 109052 3290 109076 3292
rect 109132 3290 109156 3292
rect 109212 3290 109236 3292
rect 109292 3290 109316 3292
rect 109372 3290 109386 3292
rect 109066 3238 109076 3290
rect 109132 3238 109142 3290
rect 108822 3236 108836 3238
rect 108892 3236 108916 3238
rect 108972 3236 108996 3238
rect 109052 3236 109076 3238
rect 109132 3236 109156 3238
rect 109212 3236 109236 3238
rect 109292 3236 109316 3238
rect 109372 3236 109386 3238
rect 108822 3216 109386 3236
rect 108822 2204 109386 2224
rect 108822 2202 108836 2204
rect 108892 2202 108916 2204
rect 108972 2202 108996 2204
rect 109052 2202 109076 2204
rect 109132 2202 109156 2204
rect 109212 2202 109236 2204
rect 109292 2202 109316 2204
rect 109372 2202 109386 2204
rect 109066 2150 109076 2202
rect 109132 2150 109142 2202
rect 108822 2148 108836 2150
rect 108892 2148 108916 2150
rect 108972 2148 108996 2150
rect 109052 2148 109076 2150
rect 109132 2148 109156 2150
rect 109212 2148 109236 2150
rect 109292 2148 109316 2150
rect 109372 2148 109386 2150
rect 108822 2128 109386 2148
rect 108684 1958 108804 1986
rect 108776 480 108804 1958
rect 109972 480 110000 5646
rect 110432 5574 110460 8092
rect 111628 5778 111656 8092
rect 112352 6180 112404 6186
rect 112352 6122 112404 6128
rect 111616 5772 111668 5778
rect 111616 5714 111668 5720
rect 110420 5568 110472 5574
rect 110420 5510 110472 5516
rect 111156 5568 111208 5574
rect 111156 5510 111208 5516
rect 111168 480 111196 5510
rect 112364 480 112392 6122
rect 112732 5642 112760 8092
rect 113548 5772 113600 5778
rect 113548 5714 113600 5720
rect 112720 5636 112772 5642
rect 112720 5578 112772 5584
rect 113560 480 113588 5714
rect 113928 5710 113956 8092
rect 113916 5704 113968 5710
rect 113916 5646 113968 5652
rect 114744 5704 114796 5710
rect 114744 5646 114796 5652
rect 114756 480 114784 5646
rect 115032 5574 115060 8092
rect 116228 6186 116256 8092
rect 116216 6180 116268 6186
rect 116216 6122 116268 6128
rect 117332 5778 117360 8092
rect 117320 5772 117372 5778
rect 117320 5714 117372 5720
rect 118240 5772 118292 5778
rect 118240 5714 118292 5720
rect 115940 5636 115992 5642
rect 115940 5578 115992 5584
rect 115020 5568 115072 5574
rect 115020 5510 115072 5516
rect 115952 480 115980 5578
rect 117136 5568 117188 5574
rect 117136 5510 117188 5516
rect 117148 480 117176 5510
rect 118252 480 118280 5714
rect 118436 5710 118464 8092
rect 119436 6520 119488 6526
rect 119436 6462 119488 6468
rect 118424 5704 118476 5710
rect 118424 5646 118476 5652
rect 119448 480 119476 6462
rect 119632 5642 119660 8092
rect 120632 6452 120684 6458
rect 120632 6394 120684 6400
rect 119620 5636 119672 5642
rect 119620 5578 119672 5584
rect 120644 480 120672 6394
rect 120736 5574 120764 8092
rect 121932 5778 121960 8092
rect 123036 6526 123064 8092
rect 123024 6520 123076 6526
rect 123024 6462 123076 6468
rect 124232 6458 124260 8092
rect 124220 6452 124272 6458
rect 124220 6394 124272 6400
rect 121920 5772 121972 5778
rect 121920 5714 121972 5720
rect 123024 5772 123076 5778
rect 123024 5714 123076 5720
rect 120724 5568 120776 5574
rect 120724 5510 120776 5516
rect 121828 5568 121880 5574
rect 121828 5510 121880 5516
rect 121840 480 121868 5510
rect 123036 480 123064 5714
rect 124220 5636 124272 5642
rect 124220 5578 124272 5584
rect 124232 480 124260 5578
rect 125336 5574 125364 8092
rect 126532 5778 126560 8092
rect 126822 6012 127386 6032
rect 126822 6010 126836 6012
rect 126892 6010 126916 6012
rect 126972 6010 126996 6012
rect 127052 6010 127076 6012
rect 127132 6010 127156 6012
rect 127212 6010 127236 6012
rect 127292 6010 127316 6012
rect 127372 6010 127386 6012
rect 127066 5958 127076 6010
rect 127132 5958 127142 6010
rect 126822 5956 126836 5958
rect 126892 5956 126916 5958
rect 126972 5956 126996 5958
rect 127052 5956 127076 5958
rect 127132 5956 127156 5958
rect 127212 5956 127236 5958
rect 127292 5956 127316 5958
rect 127372 5956 127386 5958
rect 126822 5936 127386 5956
rect 126520 5772 126572 5778
rect 126520 5714 126572 5720
rect 125416 5704 125468 5710
rect 125416 5646 125468 5652
rect 125324 5568 125376 5574
rect 125324 5510 125376 5516
rect 125428 480 125456 5646
rect 127636 5642 127664 8092
rect 128740 5710 128768 8092
rect 128728 5704 128780 5710
rect 128728 5646 128780 5652
rect 129004 5704 129056 5710
rect 129004 5646 129056 5652
rect 127624 5636 127676 5642
rect 127624 5578 127676 5584
rect 127808 5636 127860 5642
rect 127808 5578 127860 5584
rect 126612 5568 126664 5574
rect 126612 5510 126664 5516
rect 126624 480 126652 5510
rect 126822 4924 127386 4944
rect 126822 4922 126836 4924
rect 126892 4922 126916 4924
rect 126972 4922 126996 4924
rect 127052 4922 127076 4924
rect 127132 4922 127156 4924
rect 127212 4922 127236 4924
rect 127292 4922 127316 4924
rect 127372 4922 127386 4924
rect 127066 4870 127076 4922
rect 127132 4870 127142 4922
rect 126822 4868 126836 4870
rect 126892 4868 126916 4870
rect 126972 4868 126996 4870
rect 127052 4868 127076 4870
rect 127132 4868 127156 4870
rect 127212 4868 127236 4870
rect 127292 4868 127316 4870
rect 127372 4868 127386 4870
rect 126822 4848 127386 4868
rect 126822 3836 127386 3856
rect 126822 3834 126836 3836
rect 126892 3834 126916 3836
rect 126972 3834 126996 3836
rect 127052 3834 127076 3836
rect 127132 3834 127156 3836
rect 127212 3834 127236 3836
rect 127292 3834 127316 3836
rect 127372 3834 127386 3836
rect 127066 3782 127076 3834
rect 127132 3782 127142 3834
rect 126822 3780 126836 3782
rect 126892 3780 126916 3782
rect 126972 3780 126996 3782
rect 127052 3780 127076 3782
rect 127132 3780 127156 3782
rect 127212 3780 127236 3782
rect 127292 3780 127316 3782
rect 127372 3780 127386 3782
rect 126822 3760 127386 3780
rect 126822 2748 127386 2768
rect 126822 2746 126836 2748
rect 126892 2746 126916 2748
rect 126972 2746 126996 2748
rect 127052 2746 127076 2748
rect 127132 2746 127156 2748
rect 127212 2746 127236 2748
rect 127292 2746 127316 2748
rect 127372 2746 127386 2748
rect 127066 2694 127076 2746
rect 127132 2694 127142 2746
rect 126822 2692 126836 2694
rect 126892 2692 126916 2694
rect 126972 2692 126996 2694
rect 127052 2692 127076 2694
rect 127132 2692 127156 2694
rect 127212 2692 127236 2694
rect 127292 2692 127316 2694
rect 127372 2692 127386 2694
rect 126822 2672 127386 2692
rect 127820 480 127848 5578
rect 129016 480 129044 5646
rect 129936 5574 129964 8092
rect 131040 5642 131068 8092
rect 132236 5710 132264 8092
rect 132224 5704 132276 5710
rect 132224 5646 132276 5652
rect 132592 5704 132644 5710
rect 132592 5646 132644 5652
rect 131028 5636 131080 5642
rect 131028 5578 131080 5584
rect 131396 5636 131448 5642
rect 131396 5578 131448 5584
rect 129924 5568 129976 5574
rect 129924 5510 129976 5516
rect 130200 5568 130252 5574
rect 130200 5510 130252 5516
rect 130212 480 130240 5510
rect 131408 480 131436 5578
rect 132604 480 132632 5646
rect 133340 5574 133368 8092
rect 134536 5642 134564 8092
rect 135640 5710 135668 8092
rect 135628 5704 135680 5710
rect 135628 5646 135680 5652
rect 136088 5704 136140 5710
rect 136088 5646 136140 5652
rect 134524 5636 134576 5642
rect 134524 5578 134576 5584
rect 134892 5636 134944 5642
rect 134892 5578 134944 5584
rect 133328 5568 133380 5574
rect 133328 5510 133380 5516
rect 133788 5568 133840 5574
rect 133788 5510 133840 5516
rect 133800 480 133828 5510
rect 134904 480 134932 5578
rect 136100 480 136128 5646
rect 136836 5574 136864 8092
rect 137940 5642 137968 8092
rect 139136 5710 139164 8092
rect 139124 5704 139176 5710
rect 139124 5646 139176 5652
rect 139676 5704 139728 5710
rect 139676 5646 139728 5652
rect 137928 5636 137980 5642
rect 137928 5578 137980 5584
rect 138480 5636 138532 5642
rect 138480 5578 138532 5584
rect 136824 5568 136876 5574
rect 136824 5510 136876 5516
rect 137284 5568 137336 5574
rect 137284 5510 137336 5516
rect 137296 480 137324 5510
rect 138492 480 138520 5578
rect 139688 480 139716 5646
rect 140240 5574 140268 8092
rect 141344 5642 141372 8092
rect 142540 5710 142568 8092
rect 143264 5772 143316 5778
rect 143264 5714 143316 5720
rect 142528 5704 142580 5710
rect 142528 5646 142580 5652
rect 141332 5636 141384 5642
rect 141332 5578 141384 5584
rect 142068 5636 142120 5642
rect 142068 5578 142120 5584
rect 140228 5568 140280 5574
rect 140228 5510 140280 5516
rect 140872 5568 140924 5574
rect 140872 5510 140924 5516
rect 140884 480 140912 5510
rect 142080 480 142108 5578
rect 143276 480 143304 5714
rect 143644 5574 143672 8092
rect 144460 5704 144512 5710
rect 144460 5646 144512 5652
rect 143632 5568 143684 5574
rect 143632 5510 143684 5516
rect 144472 480 144500 5646
rect 144840 5642 144868 8092
rect 145944 5778 145972 8092
rect 145932 5772 145984 5778
rect 145932 5714 145984 5720
rect 147140 5710 147168 8092
rect 147128 5704 147180 5710
rect 147128 5646 147180 5652
rect 148048 5704 148100 5710
rect 148048 5646 148100 5652
rect 144828 5636 144880 5642
rect 144828 5578 144880 5584
rect 146852 5636 146904 5642
rect 146852 5578 146904 5584
rect 145656 5568 145708 5574
rect 145656 5510 145708 5516
rect 144822 5468 145386 5488
rect 144822 5466 144836 5468
rect 144892 5466 144916 5468
rect 144972 5466 144996 5468
rect 145052 5466 145076 5468
rect 145132 5466 145156 5468
rect 145212 5466 145236 5468
rect 145292 5466 145316 5468
rect 145372 5466 145386 5468
rect 145066 5414 145076 5466
rect 145132 5414 145142 5466
rect 144822 5412 144836 5414
rect 144892 5412 144916 5414
rect 144972 5412 144996 5414
rect 145052 5412 145076 5414
rect 145132 5412 145156 5414
rect 145212 5412 145236 5414
rect 145292 5412 145316 5414
rect 145372 5412 145386 5414
rect 144822 5392 145386 5412
rect 144822 4380 145386 4400
rect 144822 4378 144836 4380
rect 144892 4378 144916 4380
rect 144972 4378 144996 4380
rect 145052 4378 145076 4380
rect 145132 4378 145156 4380
rect 145212 4378 145236 4380
rect 145292 4378 145316 4380
rect 145372 4378 145386 4380
rect 145066 4326 145076 4378
rect 145132 4326 145142 4378
rect 144822 4324 144836 4326
rect 144892 4324 144916 4326
rect 144972 4324 144996 4326
rect 145052 4324 145076 4326
rect 145132 4324 145156 4326
rect 145212 4324 145236 4326
rect 145292 4324 145316 4326
rect 145372 4324 145386 4326
rect 144822 4304 145386 4324
rect 144822 3292 145386 3312
rect 144822 3290 144836 3292
rect 144892 3290 144916 3292
rect 144972 3290 144996 3292
rect 145052 3290 145076 3292
rect 145132 3290 145156 3292
rect 145212 3290 145236 3292
rect 145292 3290 145316 3292
rect 145372 3290 145386 3292
rect 145066 3238 145076 3290
rect 145132 3238 145142 3290
rect 144822 3236 144836 3238
rect 144892 3236 144916 3238
rect 144972 3236 144996 3238
rect 145052 3236 145076 3238
rect 145132 3236 145156 3238
rect 145212 3236 145236 3238
rect 145292 3236 145316 3238
rect 145372 3236 145386 3238
rect 144822 3216 145386 3236
rect 144822 2204 145386 2224
rect 144822 2202 144836 2204
rect 144892 2202 144916 2204
rect 144972 2202 144996 2204
rect 145052 2202 145076 2204
rect 145132 2202 145156 2204
rect 145212 2202 145236 2204
rect 145292 2202 145316 2204
rect 145372 2202 145386 2204
rect 145066 2150 145076 2202
rect 145132 2150 145142 2202
rect 144822 2148 144836 2150
rect 144892 2148 144916 2150
rect 144972 2148 144996 2150
rect 145052 2148 145076 2150
rect 145132 2148 145156 2150
rect 145212 2148 145236 2150
rect 145292 2148 145316 2150
rect 145372 2148 145386 2150
rect 144822 2128 145386 2148
rect 145668 480 145696 5510
rect 146864 480 146892 5578
rect 148060 480 148088 5646
rect 148244 5574 148272 8092
rect 149440 5642 149468 8092
rect 150544 5710 150572 8092
rect 151544 6384 151596 6390
rect 151544 6326 151596 6332
rect 150532 5704 150584 5710
rect 150532 5646 150584 5652
rect 149428 5636 149480 5642
rect 149428 5578 149480 5584
rect 150440 5636 150492 5642
rect 150440 5578 150492 5584
rect 148232 5568 148284 5574
rect 148232 5510 148284 5516
rect 149244 5568 149296 5574
rect 149244 5510 149296 5516
rect 149256 480 149284 5510
rect 150452 480 150480 5578
rect 151556 480 151584 6326
rect 151648 5574 151676 8092
rect 152740 5772 152792 5778
rect 152740 5714 152792 5720
rect 151636 5568 151688 5574
rect 151636 5510 151688 5516
rect 152752 480 152780 5714
rect 152844 5642 152872 8092
rect 153948 6390 153976 8092
rect 153936 6384 153988 6390
rect 153936 6326 153988 6332
rect 155144 5778 155172 8092
rect 155132 5772 155184 5778
rect 155132 5714 155184 5720
rect 152832 5636 152884 5642
rect 152832 5578 152884 5584
rect 155132 5636 155184 5642
rect 155132 5578 155184 5584
rect 153936 5568 153988 5574
rect 153936 5510 153988 5516
rect 153948 480 153976 5510
rect 155144 480 155172 5578
rect 156248 5574 156276 8092
rect 157444 5642 157472 8092
rect 157524 5704 157576 5710
rect 157524 5646 157576 5652
rect 157432 5636 157484 5642
rect 157432 5578 157484 5584
rect 156236 5568 156288 5574
rect 156236 5510 156288 5516
rect 156328 5568 156380 5574
rect 156328 5510 156380 5516
rect 156340 480 156368 5510
rect 157536 480 157564 5646
rect 158548 5574 158576 8092
rect 159744 5710 159772 8092
rect 159732 5704 159784 5710
rect 159732 5646 159784 5652
rect 160848 5642 160876 8092
rect 161112 6248 161164 6254
rect 161112 6190 161164 6196
rect 158720 5636 158772 5642
rect 158720 5578 158772 5584
rect 160836 5636 160888 5642
rect 160836 5578 160888 5584
rect 158536 5568 158588 5574
rect 158536 5510 158588 5516
rect 158732 480 158760 5578
rect 159916 5568 159968 5574
rect 159916 5510 159968 5516
rect 159928 480 159956 5510
rect 161124 480 161152 6190
rect 161952 5574 161980 8092
rect 163148 6254 163176 8092
rect 163136 6248 163188 6254
rect 163136 6190 163188 6196
rect 162822 6012 163386 6032
rect 162822 6010 162836 6012
rect 162892 6010 162916 6012
rect 162972 6010 162996 6012
rect 163052 6010 163076 6012
rect 163132 6010 163156 6012
rect 163212 6010 163236 6012
rect 163292 6010 163316 6012
rect 163372 6010 163386 6012
rect 163066 5958 163076 6010
rect 163132 5958 163142 6010
rect 162822 5956 162836 5958
rect 162892 5956 162916 5958
rect 162972 5956 162996 5958
rect 163052 5956 163076 5958
rect 163132 5956 163156 5958
rect 163212 5956 163236 5958
rect 163292 5956 163316 5958
rect 163372 5956 163386 5958
rect 162822 5936 163386 5956
rect 163504 5636 163556 5642
rect 163504 5578 163556 5584
rect 161940 5568 161992 5574
rect 161940 5510 161992 5516
rect 162308 5568 162360 5574
rect 162308 5510 162360 5516
rect 162320 480 162348 5510
rect 162822 4924 163386 4944
rect 162822 4922 162836 4924
rect 162892 4922 162916 4924
rect 162972 4922 162996 4924
rect 163052 4922 163076 4924
rect 163132 4922 163156 4924
rect 163212 4922 163236 4924
rect 163292 4922 163316 4924
rect 163372 4922 163386 4924
rect 163066 4870 163076 4922
rect 163132 4870 163142 4922
rect 162822 4868 162836 4870
rect 162892 4868 162916 4870
rect 162972 4868 162996 4870
rect 163052 4868 163076 4870
rect 163132 4868 163156 4870
rect 163212 4868 163236 4870
rect 163292 4868 163316 4870
rect 163372 4868 163386 4870
rect 162822 4848 163386 4868
rect 162822 3836 163386 3856
rect 162822 3834 162836 3836
rect 162892 3834 162916 3836
rect 162972 3834 162996 3836
rect 163052 3834 163076 3836
rect 163132 3834 163156 3836
rect 163212 3834 163236 3836
rect 163292 3834 163316 3836
rect 163372 3834 163386 3836
rect 163066 3782 163076 3834
rect 163132 3782 163142 3834
rect 162822 3780 162836 3782
rect 162892 3780 162916 3782
rect 162972 3780 162996 3782
rect 163052 3780 163076 3782
rect 163132 3780 163156 3782
rect 163212 3780 163236 3782
rect 163292 3780 163316 3782
rect 163372 3780 163386 3782
rect 162822 3760 163386 3780
rect 162822 2748 163386 2768
rect 162822 2746 162836 2748
rect 162892 2746 162916 2748
rect 162972 2746 162996 2748
rect 163052 2746 163076 2748
rect 163132 2746 163156 2748
rect 163212 2746 163236 2748
rect 163292 2746 163316 2748
rect 163372 2746 163386 2748
rect 163066 2694 163076 2746
rect 163132 2694 163142 2746
rect 162822 2692 162836 2694
rect 162892 2692 162916 2694
rect 162972 2692 162996 2694
rect 163052 2692 163076 2694
rect 163132 2692 163156 2694
rect 163212 2692 163236 2694
rect 163292 2692 163316 2694
rect 163372 2692 163386 2694
rect 162822 2672 163386 2692
rect 163516 480 163544 5578
rect 164252 5574 164280 8092
rect 165448 5642 165476 8092
rect 165436 5636 165488 5642
rect 165436 5578 165488 5584
rect 165896 5636 165948 5642
rect 165896 5578 165948 5584
rect 164240 5568 164292 5574
rect 164240 5510 164292 5516
rect 164700 5568 164752 5574
rect 164700 5510 164752 5516
rect 164712 480 164740 5510
rect 165908 480 165936 5578
rect 166552 5574 166580 8092
rect 167748 5642 167776 8092
rect 167736 5636 167788 5642
rect 167736 5578 167788 5584
rect 168196 5636 168248 5642
rect 168196 5578 168248 5584
rect 166540 5568 166592 5574
rect 166540 5510 166592 5516
rect 167092 5568 167144 5574
rect 167092 5510 167144 5516
rect 167104 480 167132 5510
rect 168208 480 168236 5578
rect 168852 5574 168880 8092
rect 170048 5642 170076 8092
rect 170036 5636 170088 5642
rect 170036 5578 170088 5584
rect 170588 5636 170640 5642
rect 170588 5578 170640 5584
rect 168840 5568 168892 5574
rect 168840 5510 168892 5516
rect 169392 5568 169444 5574
rect 169392 5510 169444 5516
rect 169404 480 169432 5510
rect 170600 480 170628 5578
rect 171152 5574 171180 8092
rect 171784 5704 171836 5710
rect 171784 5646 171836 5652
rect 171140 5568 171192 5574
rect 171140 5510 171192 5516
rect 171796 480 171824 5646
rect 172348 5642 172376 8092
rect 173452 5710 173480 8092
rect 173440 5704 173492 5710
rect 173440 5646 173492 5652
rect 172336 5636 172388 5642
rect 172336 5578 172388 5584
rect 174176 5636 174228 5642
rect 174176 5578 174228 5584
rect 172980 5568 173032 5574
rect 172980 5510 173032 5516
rect 172992 480 173020 5510
rect 174188 480 174216 5578
rect 174556 5574 174584 8092
rect 175752 5642 175780 8092
rect 175740 5636 175792 5642
rect 175740 5578 175792 5584
rect 176568 5636 176620 5642
rect 176568 5578 176620 5584
rect 174544 5568 174596 5574
rect 174544 5510 174596 5516
rect 175372 5568 175424 5574
rect 175372 5510 175424 5516
rect 175384 480 175412 5510
rect 176580 480 176608 5578
rect 176856 5574 176884 8092
rect 178052 5642 178080 8092
rect 178040 5636 178092 5642
rect 178040 5578 178092 5584
rect 178960 5636 179012 5642
rect 178960 5578 179012 5584
rect 176844 5568 176896 5574
rect 176844 5510 176896 5516
rect 177764 5568 177816 5574
rect 177764 5510 177816 5516
rect 177776 480 177804 5510
rect 178972 480 179000 5578
rect 179156 5574 179184 8092
rect 180352 5642 180380 8092
rect 180340 5636 180392 5642
rect 180340 5578 180392 5584
rect 181456 5574 181484 8092
rect 182652 5642 182680 8092
rect 181536 5636 181588 5642
rect 181536 5578 181588 5584
rect 182640 5636 182692 5642
rect 182640 5578 182692 5584
rect 179144 5568 179196 5574
rect 179144 5510 179196 5516
rect 180156 5568 180208 5574
rect 180156 5510 180208 5516
rect 181444 5568 181496 5574
rect 181444 5510 181496 5516
rect 180168 480 180196 5510
rect 180822 5468 181386 5488
rect 180822 5466 180836 5468
rect 180892 5466 180916 5468
rect 180972 5466 180996 5468
rect 181052 5466 181076 5468
rect 181132 5466 181156 5468
rect 181212 5466 181236 5468
rect 181292 5466 181316 5468
rect 181372 5466 181386 5468
rect 181066 5414 181076 5466
rect 181132 5414 181142 5466
rect 180822 5412 180836 5414
rect 180892 5412 180916 5414
rect 180972 5412 180996 5414
rect 181052 5412 181076 5414
rect 181132 5412 181156 5414
rect 181212 5412 181236 5414
rect 181292 5412 181316 5414
rect 181372 5412 181386 5414
rect 180822 5392 181386 5412
rect 180822 4380 181386 4400
rect 180822 4378 180836 4380
rect 180892 4378 180916 4380
rect 180972 4378 180996 4380
rect 181052 4378 181076 4380
rect 181132 4378 181156 4380
rect 181212 4378 181236 4380
rect 181292 4378 181316 4380
rect 181372 4378 181386 4380
rect 181066 4326 181076 4378
rect 181132 4326 181142 4378
rect 180822 4324 180836 4326
rect 180892 4324 180916 4326
rect 180972 4324 180996 4326
rect 181052 4324 181076 4326
rect 181132 4324 181156 4326
rect 181212 4324 181236 4326
rect 181292 4324 181316 4326
rect 181372 4324 181386 4326
rect 180822 4304 181386 4324
rect 180822 3292 181386 3312
rect 180822 3290 180836 3292
rect 180892 3290 180916 3292
rect 180972 3290 180996 3292
rect 181052 3290 181076 3292
rect 181132 3290 181156 3292
rect 181212 3290 181236 3292
rect 181292 3290 181316 3292
rect 181372 3290 181386 3292
rect 181066 3238 181076 3290
rect 181132 3238 181142 3290
rect 180822 3236 180836 3238
rect 180892 3236 180916 3238
rect 180972 3236 180996 3238
rect 181052 3236 181076 3238
rect 181132 3236 181156 3238
rect 181212 3236 181236 3238
rect 181292 3236 181316 3238
rect 181372 3236 181386 3238
rect 180822 3216 181386 3236
rect 180822 2204 181386 2224
rect 180822 2202 180836 2204
rect 180892 2202 180916 2204
rect 180972 2202 180996 2204
rect 181052 2202 181076 2204
rect 181132 2202 181156 2204
rect 181212 2202 181236 2204
rect 181292 2202 181316 2204
rect 181372 2202 181386 2204
rect 181066 2150 181076 2202
rect 181132 2150 181142 2202
rect 180822 2148 180836 2150
rect 180892 2148 180916 2150
rect 180972 2148 180996 2150
rect 181052 2148 181076 2150
rect 181132 2148 181156 2150
rect 181212 2148 181236 2150
rect 181292 2148 181316 2150
rect 181372 2148 181386 2150
rect 180822 2128 181386 2148
rect 181548 1986 181576 5578
rect 183756 5574 183784 8092
rect 184756 5704 184808 5710
rect 184756 5646 184808 5652
rect 182548 5568 182600 5574
rect 182548 5510 182600 5516
rect 183744 5568 183796 5574
rect 183744 5510 183796 5516
rect 181364 1958 181576 1986
rect 181364 480 181392 1958
rect 182560 480 182588 5510
rect 183744 3528 183796 3534
rect 183744 3470 183796 3476
rect 183756 480 183784 3470
rect 184768 3346 184796 5646
rect 184860 3534 184888 8092
rect 186056 5710 186084 8092
rect 186044 5704 186096 5710
rect 186044 5646 186096 5652
rect 187160 5574 187188 8092
rect 188356 5574 188384 8092
rect 189460 5574 189488 8092
rect 190656 5574 190684 8092
rect 186044 5568 186096 5574
rect 186044 5510 186096 5516
rect 187148 5568 187200 5574
rect 187148 5510 187200 5516
rect 187240 5568 187292 5574
rect 187240 5510 187292 5516
rect 188344 5568 188396 5574
rect 188344 5510 188396 5516
rect 188436 5568 188488 5574
rect 188436 5510 188488 5516
rect 189448 5568 189500 5574
rect 189448 5510 189500 5516
rect 189632 5568 189684 5574
rect 189632 5510 189684 5516
rect 190644 5568 190696 5574
rect 190644 5510 190696 5516
rect 184848 3528 184900 3534
rect 184848 3470 184900 3476
rect 184768 3318 184888 3346
rect 184860 480 184888 3318
rect 186056 480 186084 5510
rect 187252 480 187280 5510
rect 188448 480 188476 5510
rect 189644 480 189672 5510
rect 191760 3534 191788 8092
rect 192956 3534 192984 8092
rect 194060 3534 194088 8092
rect 195164 5574 195192 8092
rect 195992 8078 196374 8106
rect 195992 5658 196020 8078
rect 195716 5630 196020 5658
rect 194416 5568 194468 5574
rect 194416 5510 194468 5516
rect 195152 5568 195204 5574
rect 195152 5510 195204 5516
rect 190828 3528 190880 3534
rect 190828 3470 190880 3476
rect 191748 3528 191800 3534
rect 191748 3470 191800 3476
rect 192024 3528 192076 3534
rect 192024 3470 192076 3476
rect 192944 3528 192996 3534
rect 192944 3470 192996 3476
rect 193220 3528 193272 3534
rect 193220 3470 193272 3476
rect 194048 3528 194100 3534
rect 194048 3470 194100 3476
rect 190840 480 190868 3470
rect 192036 480 192064 3470
rect 193232 480 193260 3470
rect 194428 480 194456 5510
rect 195716 626 195744 5630
rect 197464 5574 197492 8092
rect 198016 8078 198674 8106
rect 199488 8078 199778 8106
rect 200408 8078 200974 8106
rect 201512 8078 202078 8106
rect 196808 5568 196860 5574
rect 196808 5510 196860 5516
rect 197452 5568 197504 5574
rect 197452 5510 197504 5516
rect 195624 598 195744 626
rect 195624 480 195652 598
rect 196820 480 196848 5510
rect 198016 480 198044 8078
rect 198822 6012 199386 6032
rect 198822 6010 198836 6012
rect 198892 6010 198916 6012
rect 198972 6010 198996 6012
rect 199052 6010 199076 6012
rect 199132 6010 199156 6012
rect 199212 6010 199236 6012
rect 199292 6010 199316 6012
rect 199372 6010 199386 6012
rect 199066 5958 199076 6010
rect 199132 5958 199142 6010
rect 198822 5956 198836 5958
rect 198892 5956 198916 5958
rect 198972 5956 198996 5958
rect 199052 5956 199076 5958
rect 199132 5956 199156 5958
rect 199212 5956 199236 5958
rect 199292 5956 199316 5958
rect 199372 5956 199386 5958
rect 198822 5936 199386 5956
rect 198822 4924 199386 4944
rect 198822 4922 198836 4924
rect 198892 4922 198916 4924
rect 198972 4922 198996 4924
rect 199052 4922 199076 4924
rect 199132 4922 199156 4924
rect 199212 4922 199236 4924
rect 199292 4922 199316 4924
rect 199372 4922 199386 4924
rect 199066 4870 199076 4922
rect 199132 4870 199142 4922
rect 198822 4868 198836 4870
rect 198892 4868 198916 4870
rect 198972 4868 198996 4870
rect 199052 4868 199076 4870
rect 199132 4868 199156 4870
rect 199212 4868 199236 4870
rect 199292 4868 199316 4870
rect 199372 4868 199386 4870
rect 198822 4848 199386 4868
rect 198822 3836 199386 3856
rect 198822 3834 198836 3836
rect 198892 3834 198916 3836
rect 198972 3834 198996 3836
rect 199052 3834 199076 3836
rect 199132 3834 199156 3836
rect 199212 3834 199236 3836
rect 199292 3834 199316 3836
rect 199372 3834 199386 3836
rect 199066 3782 199076 3834
rect 199132 3782 199142 3834
rect 198822 3780 198836 3782
rect 198892 3780 198916 3782
rect 198972 3780 198996 3782
rect 199052 3780 199076 3782
rect 199132 3780 199156 3782
rect 199212 3780 199236 3782
rect 199292 3780 199316 3782
rect 199372 3780 199386 3782
rect 198822 3760 199386 3780
rect 198822 2748 199386 2768
rect 198822 2746 198836 2748
rect 198892 2746 198916 2748
rect 198972 2746 198996 2748
rect 199052 2746 199076 2748
rect 199132 2746 199156 2748
rect 199212 2746 199236 2748
rect 199292 2746 199316 2748
rect 199372 2746 199386 2748
rect 199066 2694 199076 2746
rect 199132 2694 199142 2746
rect 198822 2692 198836 2694
rect 198892 2692 198916 2694
rect 198972 2692 198996 2694
rect 199052 2692 199076 2694
rect 199132 2692 199156 2694
rect 199212 2692 199236 2694
rect 199292 2692 199316 2694
rect 199372 2692 199386 2694
rect 198822 2672 199386 2692
rect 199488 2530 199516 8078
rect 199212 2502 199516 2530
rect 199212 480 199240 2502
rect 200408 480 200436 8078
rect 201512 480 201540 8078
rect 203260 5574 203288 8092
rect 204272 8078 204378 8106
rect 205100 8078 205482 8106
rect 206296 8078 206678 8106
rect 207492 8078 207782 8106
rect 208688 8078 208978 8106
rect 209884 8078 210082 8106
rect 211172 8078 211278 8106
rect 212276 8078 212382 8106
rect 213472 8078 213578 8106
rect 204272 5658 204300 8078
rect 203996 5630 204300 5658
rect 202696 5568 202748 5574
rect 202696 5510 202748 5516
rect 203248 5568 203300 5574
rect 203248 5510 203300 5516
rect 202708 480 202736 5510
rect 203996 626 204024 5630
rect 203904 598 204024 626
rect 203904 480 203932 598
rect 205100 480 205128 8078
rect 206296 480 206324 8078
rect 207492 480 207520 8078
rect 208688 480 208716 8078
rect 209884 480 209912 8078
rect 211172 5658 211200 8078
rect 210988 5630 211200 5658
rect 210988 626 211016 5630
rect 210988 598 211108 626
rect 211080 480 211108 598
rect 212276 480 212304 8078
rect 213472 480 213500 8078
rect 214668 480 214696 8092
rect 215864 480 215892 8092
rect 216692 8078 216982 8106
rect 218086 8078 218192 8106
rect 219282 8078 219388 8106
rect 220386 8078 220584 8106
rect 221582 8078 221780 8106
rect 222686 8078 222976 8106
rect 223882 8078 224172 8106
rect 224986 8078 225368 8106
rect 226182 8078 226288 8106
rect 227286 8078 227668 8106
rect 228390 8078 228956 8106
rect 229586 8078 230152 8106
rect 230690 8078 231348 8106
rect 231886 8078 232544 8106
rect 216692 1986 216720 8078
rect 216822 5468 217386 5488
rect 216822 5466 216836 5468
rect 216892 5466 216916 5468
rect 216972 5466 216996 5468
rect 217052 5466 217076 5468
rect 217132 5466 217156 5468
rect 217212 5466 217236 5468
rect 217292 5466 217316 5468
rect 217372 5466 217386 5468
rect 217066 5414 217076 5466
rect 217132 5414 217142 5466
rect 216822 5412 216836 5414
rect 216892 5412 216916 5414
rect 216972 5412 216996 5414
rect 217052 5412 217076 5414
rect 217132 5412 217156 5414
rect 217212 5412 217236 5414
rect 217292 5412 217316 5414
rect 217372 5412 217386 5414
rect 216822 5392 217386 5412
rect 216822 4380 217386 4400
rect 216822 4378 216836 4380
rect 216892 4378 216916 4380
rect 216972 4378 216996 4380
rect 217052 4378 217076 4380
rect 217132 4378 217156 4380
rect 217212 4378 217236 4380
rect 217292 4378 217316 4380
rect 217372 4378 217386 4380
rect 217066 4326 217076 4378
rect 217132 4326 217142 4378
rect 216822 4324 216836 4326
rect 216892 4324 216916 4326
rect 216972 4324 216996 4326
rect 217052 4324 217076 4326
rect 217132 4324 217156 4326
rect 217212 4324 217236 4326
rect 217292 4324 217316 4326
rect 217372 4324 217386 4326
rect 216822 4304 217386 4324
rect 216822 3292 217386 3312
rect 216822 3290 216836 3292
rect 216892 3290 216916 3292
rect 216972 3290 216996 3292
rect 217052 3290 217076 3292
rect 217132 3290 217156 3292
rect 217212 3290 217236 3292
rect 217292 3290 217316 3292
rect 217372 3290 217386 3292
rect 217066 3238 217076 3290
rect 217132 3238 217142 3290
rect 216822 3236 216836 3238
rect 216892 3236 216916 3238
rect 216972 3236 216996 3238
rect 217052 3236 217076 3238
rect 217132 3236 217156 3238
rect 217212 3236 217236 3238
rect 217292 3236 217316 3238
rect 217372 3236 217386 3238
rect 216822 3216 217386 3236
rect 216822 2204 217386 2224
rect 216822 2202 216836 2204
rect 216892 2202 216916 2204
rect 216972 2202 216996 2204
rect 217052 2202 217076 2204
rect 217132 2202 217156 2204
rect 217212 2202 217236 2204
rect 217292 2202 217316 2204
rect 217372 2202 217386 2204
rect 217066 2150 217076 2202
rect 217132 2150 217142 2202
rect 216822 2148 216836 2150
rect 216892 2148 216916 2150
rect 216972 2148 216996 2150
rect 217052 2148 217076 2150
rect 217132 2148 217156 2150
rect 217212 2148 217236 2150
rect 217292 2148 217316 2150
rect 217372 2148 217386 2150
rect 216822 2128 217386 2148
rect 216692 1958 217088 1986
rect 217060 480 217088 1958
rect 218164 480 218192 8078
rect 219360 480 219388 8078
rect 220556 480 220584 8078
rect 221752 480 221780 8078
rect 222948 480 222976 8078
rect 224144 480 224172 8078
rect 225340 480 225368 8078
rect 226260 5658 226288 8078
rect 227640 5658 227668 8078
rect 226260 5630 226380 5658
rect 227640 5630 227852 5658
rect 226352 610 226380 5630
rect 227824 626 227852 5630
rect 226340 604 226392 610
rect 226340 546 226392 552
rect 226524 604 226576 610
rect 226524 546 226576 552
rect 227732 598 227852 626
rect 226536 480 226564 546
rect 227732 480 227760 598
rect 228928 480 228956 8078
rect 230124 480 230152 8078
rect 231320 480 231348 8078
rect 232516 480 232544 8078
rect 232976 5574 233004 8092
rect 234186 8078 234568 8106
rect 235290 8078 235948 8106
rect 234540 5658 234568 8078
rect 234822 6012 235386 6032
rect 234822 6010 234836 6012
rect 234892 6010 234916 6012
rect 234972 6010 234996 6012
rect 235052 6010 235076 6012
rect 235132 6010 235156 6012
rect 235212 6010 235236 6012
rect 235292 6010 235316 6012
rect 235372 6010 235386 6012
rect 235066 5958 235076 6010
rect 235132 5958 235142 6010
rect 234822 5956 234836 5958
rect 234892 5956 234916 5958
rect 234972 5956 234996 5958
rect 235052 5956 235076 5958
rect 235132 5956 235156 5958
rect 235212 5956 235236 5958
rect 235292 5956 235316 5958
rect 235372 5956 235386 5958
rect 234822 5936 235386 5956
rect 235920 5658 235948 8078
rect 234540 5630 234660 5658
rect 235920 5630 236132 5658
rect 232964 5568 233016 5574
rect 232964 5510 233016 5516
rect 233700 5568 233752 5574
rect 233700 5510 233752 5516
rect 233712 480 233740 5510
rect 234632 2394 234660 5630
rect 234822 4924 235386 4944
rect 234822 4922 234836 4924
rect 234892 4922 234916 4924
rect 234972 4922 234996 4924
rect 235052 4922 235076 4924
rect 235132 4922 235156 4924
rect 235212 4922 235236 4924
rect 235292 4922 235316 4924
rect 235372 4922 235386 4924
rect 235066 4870 235076 4922
rect 235132 4870 235142 4922
rect 234822 4868 234836 4870
rect 234892 4868 234916 4870
rect 234972 4868 234996 4870
rect 235052 4868 235076 4870
rect 235132 4868 235156 4870
rect 235212 4868 235236 4870
rect 235292 4868 235316 4870
rect 235372 4868 235386 4870
rect 234822 4848 235386 4868
rect 234822 3836 235386 3856
rect 234822 3834 234836 3836
rect 234892 3834 234916 3836
rect 234972 3834 234996 3836
rect 235052 3834 235076 3836
rect 235132 3834 235156 3836
rect 235212 3834 235236 3836
rect 235292 3834 235316 3836
rect 235372 3834 235386 3836
rect 235066 3782 235076 3834
rect 235132 3782 235142 3834
rect 234822 3780 234836 3782
rect 234892 3780 234916 3782
rect 234972 3780 234996 3782
rect 235052 3780 235076 3782
rect 235132 3780 235156 3782
rect 235212 3780 235236 3782
rect 235292 3780 235316 3782
rect 235372 3780 235386 3782
rect 234822 3760 235386 3780
rect 234822 2748 235386 2768
rect 234822 2746 234836 2748
rect 234892 2746 234916 2748
rect 234972 2746 234996 2748
rect 235052 2746 235076 2748
rect 235132 2746 235156 2748
rect 235212 2746 235236 2748
rect 235292 2746 235316 2748
rect 235372 2746 235386 2748
rect 235066 2694 235076 2746
rect 235132 2694 235142 2746
rect 234822 2692 234836 2694
rect 234892 2692 234916 2694
rect 234972 2692 234996 2694
rect 235052 2692 235076 2694
rect 235132 2692 235156 2694
rect 235212 2692 235236 2694
rect 235292 2692 235316 2694
rect 235372 2692 235386 2694
rect 234822 2672 235386 2692
rect 234632 2366 234844 2394
rect 234816 480 234844 2366
rect 236104 626 236132 5630
rect 236472 3534 236500 8092
rect 237576 3534 237604 8092
rect 238680 5574 238708 8092
rect 239876 5574 239904 8092
rect 240980 5574 241008 8092
rect 242176 5574 242204 8092
rect 243280 5574 243308 8092
rect 238668 5568 238720 5574
rect 238668 5510 238720 5516
rect 239588 5568 239640 5574
rect 239588 5510 239640 5516
rect 239864 5568 239916 5574
rect 239864 5510 239916 5516
rect 240784 5568 240836 5574
rect 240784 5510 240836 5516
rect 240968 5568 241020 5574
rect 240968 5510 241020 5516
rect 241980 5568 242032 5574
rect 241980 5510 242032 5516
rect 242164 5568 242216 5574
rect 242164 5510 242216 5516
rect 243176 5568 243228 5574
rect 243176 5510 243228 5516
rect 243268 5568 243320 5574
rect 243268 5510 243320 5516
rect 244372 5568 244424 5574
rect 244372 5510 244424 5516
rect 236460 3528 236512 3534
rect 236460 3470 236512 3476
rect 237196 3528 237248 3534
rect 237196 3470 237248 3476
rect 237564 3528 237616 3534
rect 237564 3470 237616 3476
rect 238392 3528 238444 3534
rect 238392 3470 238444 3476
rect 236012 598 236132 626
rect 236012 480 236040 598
rect 237208 480 237236 3470
rect 238404 480 238432 3470
rect 239600 480 239628 5510
rect 240796 480 240824 5510
rect 241992 480 242020 5510
rect 243188 480 243216 5510
rect 244384 480 244412 5510
rect 244476 3534 244504 8092
rect 245580 5574 245608 8092
rect 246776 5574 246804 8092
rect 247880 5642 247908 8092
rect 248984 5710 249012 8092
rect 248972 5704 249024 5710
rect 248972 5646 249024 5652
rect 247868 5636 247920 5642
rect 247868 5578 247920 5584
rect 249156 5636 249208 5642
rect 249156 5578 249208 5584
rect 245568 5568 245620 5574
rect 245568 5510 245620 5516
rect 246672 5568 246724 5574
rect 246672 5510 246724 5516
rect 246764 5568 246816 5574
rect 246764 5510 246816 5516
rect 247960 5568 248012 5574
rect 247960 5510 248012 5516
rect 244464 3528 244516 3534
rect 244464 3470 244516 3476
rect 245568 3528 245620 3534
rect 245568 3470 245620 3476
rect 246684 3482 246712 5510
rect 245580 480 245608 3470
rect 246684 3454 246804 3482
rect 246776 480 246804 3454
rect 247972 480 248000 5510
rect 249168 480 249196 5578
rect 250180 5574 250208 8092
rect 250352 5704 250404 5710
rect 250352 5646 250404 5652
rect 250168 5568 250220 5574
rect 250168 5510 250220 5516
rect 250364 480 250392 5646
rect 251284 5642 251312 8092
rect 251272 5636 251324 5642
rect 251272 5578 251324 5584
rect 252480 5574 252508 8092
rect 253584 5642 253612 8092
rect 252652 5636 252704 5642
rect 252652 5578 252704 5584
rect 253572 5636 253624 5642
rect 253572 5578 253624 5584
rect 251456 5568 251508 5574
rect 251456 5510 251508 5516
rect 252468 5568 252520 5574
rect 252468 5510 252520 5516
rect 251468 480 251496 5510
rect 252664 480 252692 5578
rect 254780 5574 254808 8092
rect 255884 5642 255912 8092
rect 255044 5636 255096 5642
rect 255044 5578 255096 5584
rect 255872 5636 255924 5642
rect 255872 5578 255924 5584
rect 253848 5568 253900 5574
rect 253848 5510 253900 5516
rect 254768 5568 254820 5574
rect 254768 5510 254820 5516
rect 252822 5468 253386 5488
rect 252822 5466 252836 5468
rect 252892 5466 252916 5468
rect 252972 5466 252996 5468
rect 253052 5466 253076 5468
rect 253132 5466 253156 5468
rect 253212 5466 253236 5468
rect 253292 5466 253316 5468
rect 253372 5466 253386 5468
rect 253066 5414 253076 5466
rect 253132 5414 253142 5466
rect 252822 5412 252836 5414
rect 252892 5412 252916 5414
rect 252972 5412 252996 5414
rect 253052 5412 253076 5414
rect 253132 5412 253156 5414
rect 253212 5412 253236 5414
rect 253292 5412 253316 5414
rect 253372 5412 253386 5414
rect 252822 5392 253386 5412
rect 252822 4380 253386 4400
rect 252822 4378 252836 4380
rect 252892 4378 252916 4380
rect 252972 4378 252996 4380
rect 253052 4378 253076 4380
rect 253132 4378 253156 4380
rect 253212 4378 253236 4380
rect 253292 4378 253316 4380
rect 253372 4378 253386 4380
rect 253066 4326 253076 4378
rect 253132 4326 253142 4378
rect 252822 4324 252836 4326
rect 252892 4324 252916 4326
rect 252972 4324 252996 4326
rect 253052 4324 253076 4326
rect 253132 4324 253156 4326
rect 253212 4324 253236 4326
rect 253292 4324 253316 4326
rect 253372 4324 253386 4326
rect 252822 4304 253386 4324
rect 252822 3292 253386 3312
rect 252822 3290 252836 3292
rect 252892 3290 252916 3292
rect 252972 3290 252996 3292
rect 253052 3290 253076 3292
rect 253132 3290 253156 3292
rect 253212 3290 253236 3292
rect 253292 3290 253316 3292
rect 253372 3290 253386 3292
rect 253066 3238 253076 3290
rect 253132 3238 253142 3290
rect 252822 3236 252836 3238
rect 252892 3236 252916 3238
rect 252972 3236 252996 3238
rect 253052 3236 253076 3238
rect 253132 3236 253156 3238
rect 253212 3236 253236 3238
rect 253292 3236 253316 3238
rect 253372 3236 253386 3238
rect 252822 3216 253386 3236
rect 252822 2204 253386 2224
rect 252822 2202 252836 2204
rect 252892 2202 252916 2204
rect 252972 2202 252996 2204
rect 253052 2202 253076 2204
rect 253132 2202 253156 2204
rect 253212 2202 253236 2204
rect 253292 2202 253316 2204
rect 253372 2202 253386 2204
rect 253066 2150 253076 2202
rect 253132 2150 253142 2202
rect 252822 2148 252836 2150
rect 252892 2148 252916 2150
rect 252972 2148 252996 2150
rect 253052 2148 253076 2150
rect 253132 2148 253156 2150
rect 253212 2148 253236 2150
rect 253292 2148 253316 2150
rect 253372 2148 253386 2150
rect 252822 2128 253386 2148
rect 253860 480 253888 5510
rect 255056 480 255084 5578
rect 257080 5574 257108 8092
rect 258184 5642 258212 8092
rect 257436 5636 257488 5642
rect 257436 5578 257488 5584
rect 258172 5636 258224 5642
rect 258172 5578 258224 5584
rect 256240 5568 256292 5574
rect 256240 5510 256292 5516
rect 257068 5568 257120 5574
rect 257068 5510 257120 5516
rect 256252 480 256280 5510
rect 257448 480 257476 5578
rect 259380 5574 259408 8092
rect 260484 5642 260512 8092
rect 259828 5636 259880 5642
rect 259828 5578 259880 5584
rect 260472 5636 260524 5642
rect 260472 5578 260524 5584
rect 258632 5568 258684 5574
rect 258632 5510 258684 5516
rect 259368 5568 259420 5574
rect 259368 5510 259420 5516
rect 258644 480 258672 5510
rect 259840 480 259868 5578
rect 261588 5574 261616 8092
rect 262784 5642 262812 8092
rect 262220 5636 262272 5642
rect 262220 5578 262272 5584
rect 262772 5636 262824 5642
rect 262772 5578 262824 5584
rect 261024 5568 261076 5574
rect 261024 5510 261076 5516
rect 261576 5568 261628 5574
rect 261576 5510 261628 5516
rect 261036 480 261064 5510
rect 262232 480 262260 5578
rect 263888 5574 263916 8092
rect 265084 5642 265112 8092
rect 266188 5710 266216 8092
rect 266176 5704 266228 5710
rect 266176 5646 266228 5652
rect 264612 5636 264664 5642
rect 264612 5578 264664 5584
rect 265072 5636 265124 5642
rect 265072 5578 265124 5584
rect 267004 5636 267056 5642
rect 267004 5578 267056 5584
rect 263416 5568 263468 5574
rect 263416 5510 263468 5516
rect 263876 5568 263928 5574
rect 263876 5510 263928 5516
rect 263428 480 263456 5510
rect 264624 480 264652 5578
rect 265808 5568 265860 5574
rect 265808 5510 265860 5516
rect 265820 480 265848 5510
rect 267016 480 267044 5578
rect 267384 5574 267412 8092
rect 268108 5704 268160 5710
rect 268108 5646 268160 5652
rect 267372 5568 267424 5574
rect 267372 5510 267424 5516
rect 268120 480 268148 5646
rect 268488 5642 268516 8092
rect 268476 5636 268528 5642
rect 268476 5578 268528 5584
rect 269684 5574 269712 8092
rect 270788 6186 270816 8092
rect 270776 6180 270828 6186
rect 270776 6122 270828 6128
rect 270822 6012 271386 6032
rect 270822 6010 270836 6012
rect 270892 6010 270916 6012
rect 270972 6010 270996 6012
rect 271052 6010 271076 6012
rect 271132 6010 271156 6012
rect 271212 6010 271236 6012
rect 271292 6010 271316 6012
rect 271372 6010 271386 6012
rect 271066 5958 271076 6010
rect 271132 5958 271142 6010
rect 270822 5956 270836 5958
rect 270892 5956 270916 5958
rect 270972 5956 270996 5958
rect 271052 5956 271076 5958
rect 271132 5956 271156 5958
rect 271212 5956 271236 5958
rect 271292 5956 271316 5958
rect 271372 5956 271386 5958
rect 270822 5936 271386 5956
rect 270500 5636 270552 5642
rect 270500 5578 270552 5584
rect 269304 5568 269356 5574
rect 269304 5510 269356 5516
rect 269672 5568 269724 5574
rect 269672 5510 269724 5516
rect 269316 480 269344 5510
rect 270512 480 270540 5578
rect 271892 5574 271920 8092
rect 272892 6180 272944 6186
rect 272892 6122 272944 6128
rect 271696 5568 271748 5574
rect 271696 5510 271748 5516
rect 271880 5568 271932 5574
rect 271880 5510 271932 5516
rect 270822 4924 271386 4944
rect 270822 4922 270836 4924
rect 270892 4922 270916 4924
rect 270972 4922 270996 4924
rect 271052 4922 271076 4924
rect 271132 4922 271156 4924
rect 271212 4922 271236 4924
rect 271292 4922 271316 4924
rect 271372 4922 271386 4924
rect 271066 4870 271076 4922
rect 271132 4870 271142 4922
rect 270822 4868 270836 4870
rect 270892 4868 270916 4870
rect 270972 4868 270996 4870
rect 271052 4868 271076 4870
rect 271132 4868 271156 4870
rect 271212 4868 271236 4870
rect 271292 4868 271316 4870
rect 271372 4868 271386 4870
rect 270822 4848 271386 4868
rect 270822 3836 271386 3856
rect 270822 3834 270836 3836
rect 270892 3834 270916 3836
rect 270972 3834 270996 3836
rect 271052 3834 271076 3836
rect 271132 3834 271156 3836
rect 271212 3834 271236 3836
rect 271292 3834 271316 3836
rect 271372 3834 271386 3836
rect 271066 3782 271076 3834
rect 271132 3782 271142 3834
rect 270822 3780 270836 3782
rect 270892 3780 270916 3782
rect 270972 3780 270996 3782
rect 271052 3780 271076 3782
rect 271132 3780 271156 3782
rect 271212 3780 271236 3782
rect 271292 3780 271316 3782
rect 271372 3780 271386 3782
rect 270822 3760 271386 3780
rect 270822 2748 271386 2768
rect 270822 2746 270836 2748
rect 270892 2746 270916 2748
rect 270972 2746 270996 2748
rect 271052 2746 271076 2748
rect 271132 2746 271156 2748
rect 271212 2746 271236 2748
rect 271292 2746 271316 2748
rect 271372 2746 271386 2748
rect 271066 2694 271076 2746
rect 271132 2694 271142 2746
rect 270822 2692 270836 2694
rect 270892 2692 270916 2694
rect 270972 2692 270996 2694
rect 271052 2692 271076 2694
rect 271132 2692 271156 2694
rect 271212 2692 271236 2694
rect 271292 2692 271316 2694
rect 271372 2692 271386 2694
rect 270822 2672 271386 2692
rect 271708 480 271736 5510
rect 272904 480 272932 6122
rect 273088 5642 273116 8092
rect 273076 5636 273128 5642
rect 273076 5578 273128 5584
rect 274192 5574 274220 8092
rect 275388 5642 275416 8092
rect 276492 5710 276520 8092
rect 277688 5778 277716 8092
rect 277676 5772 277728 5778
rect 277676 5714 277728 5720
rect 276480 5704 276532 5710
rect 276480 5646 276532 5652
rect 275284 5636 275336 5642
rect 275284 5578 275336 5584
rect 275376 5636 275428 5642
rect 275376 5578 275428 5584
rect 277676 5636 277728 5642
rect 277676 5578 277728 5584
rect 274088 5568 274140 5574
rect 274088 5510 274140 5516
rect 274180 5568 274232 5574
rect 274180 5510 274232 5516
rect 274100 480 274128 5510
rect 275296 480 275324 5578
rect 276480 5568 276532 5574
rect 276480 5510 276532 5516
rect 276492 480 276520 5510
rect 277688 480 277716 5578
rect 278792 5574 278820 8092
rect 278872 5704 278924 5710
rect 278872 5646 278924 5652
rect 278780 5568 278832 5574
rect 278780 5510 278832 5516
rect 278884 480 278912 5646
rect 279988 5642 280016 8092
rect 280068 5772 280120 5778
rect 280068 5714 280120 5720
rect 279976 5636 280028 5642
rect 279976 5578 280028 5584
rect 280080 480 280108 5714
rect 281092 5710 281120 8092
rect 282196 5778 282224 8092
rect 283392 5846 283420 8092
rect 283380 5840 283432 5846
rect 283380 5782 283432 5788
rect 282184 5772 282236 5778
rect 282184 5714 282236 5720
rect 281080 5704 281132 5710
rect 281080 5646 281132 5652
rect 283656 5704 283708 5710
rect 283656 5646 283708 5652
rect 282460 5636 282512 5642
rect 282460 5578 282512 5584
rect 281264 5568 281316 5574
rect 281264 5510 281316 5516
rect 281276 480 281304 5510
rect 282472 480 282500 5578
rect 283668 480 283696 5646
rect 284496 5574 284524 8092
rect 284760 5772 284812 5778
rect 284760 5714 284812 5720
rect 284484 5568 284536 5574
rect 284484 5510 284536 5516
rect 284772 480 284800 5714
rect 285692 5642 285720 8092
rect 285956 5840 286008 5846
rect 285956 5782 286008 5788
rect 285680 5636 285732 5642
rect 285680 5578 285732 5584
rect 285968 480 285996 5782
rect 286796 5710 286824 8092
rect 286784 5704 286836 5710
rect 286784 5646 286836 5652
rect 287992 5574 288020 8092
rect 289096 5642 289124 8092
rect 290292 5710 290320 8092
rect 291396 5778 291424 8092
rect 292592 5846 292620 8092
rect 292580 5840 292632 5846
rect 292580 5782 292632 5788
rect 291384 5772 291436 5778
rect 291384 5714 291436 5720
rect 289544 5704 289596 5710
rect 289544 5646 289596 5652
rect 290280 5704 290332 5710
rect 290280 5646 290332 5652
rect 293132 5704 293184 5710
rect 293132 5646 293184 5652
rect 288348 5636 288400 5642
rect 288348 5578 288400 5584
rect 289084 5636 289136 5642
rect 289084 5578 289136 5584
rect 287152 5568 287204 5574
rect 287152 5510 287204 5516
rect 287980 5568 288032 5574
rect 287980 5510 288032 5516
rect 287164 480 287192 5510
rect 288360 480 288388 5578
rect 288822 5468 289386 5488
rect 288822 5466 288836 5468
rect 288892 5466 288916 5468
rect 288972 5466 288996 5468
rect 289052 5466 289076 5468
rect 289132 5466 289156 5468
rect 289212 5466 289236 5468
rect 289292 5466 289316 5468
rect 289372 5466 289386 5468
rect 289066 5414 289076 5466
rect 289132 5414 289142 5466
rect 288822 5412 288836 5414
rect 288892 5412 288916 5414
rect 288972 5412 288996 5414
rect 289052 5412 289076 5414
rect 289132 5412 289156 5414
rect 289212 5412 289236 5414
rect 289292 5412 289316 5414
rect 289372 5412 289386 5414
rect 288822 5392 289386 5412
rect 288822 4380 289386 4400
rect 288822 4378 288836 4380
rect 288892 4378 288916 4380
rect 288972 4378 288996 4380
rect 289052 4378 289076 4380
rect 289132 4378 289156 4380
rect 289212 4378 289236 4380
rect 289292 4378 289316 4380
rect 289372 4378 289386 4380
rect 289066 4326 289076 4378
rect 289132 4326 289142 4378
rect 288822 4324 288836 4326
rect 288892 4324 288916 4326
rect 288972 4324 288996 4326
rect 289052 4324 289076 4326
rect 289132 4324 289156 4326
rect 289212 4324 289236 4326
rect 289292 4324 289316 4326
rect 289372 4324 289386 4326
rect 288822 4304 289386 4324
rect 288822 3292 289386 3312
rect 288822 3290 288836 3292
rect 288892 3290 288916 3292
rect 288972 3290 288996 3292
rect 289052 3290 289076 3292
rect 289132 3290 289156 3292
rect 289212 3290 289236 3292
rect 289292 3290 289316 3292
rect 289372 3290 289386 3292
rect 289066 3238 289076 3290
rect 289132 3238 289142 3290
rect 288822 3236 288836 3238
rect 288892 3236 288916 3238
rect 288972 3236 288996 3238
rect 289052 3236 289076 3238
rect 289132 3236 289156 3238
rect 289212 3236 289236 3238
rect 289292 3236 289316 3238
rect 289372 3236 289386 3238
rect 288822 3216 289386 3236
rect 288822 2204 289386 2224
rect 288822 2202 288836 2204
rect 288892 2202 288916 2204
rect 288972 2202 288996 2204
rect 289052 2202 289076 2204
rect 289132 2202 289156 2204
rect 289212 2202 289236 2204
rect 289292 2202 289316 2204
rect 289372 2202 289386 2204
rect 289066 2150 289076 2202
rect 289132 2150 289142 2202
rect 288822 2148 288836 2150
rect 288892 2148 288916 2150
rect 288972 2148 288996 2150
rect 289052 2148 289076 2150
rect 289132 2148 289156 2150
rect 289212 2148 289236 2150
rect 289292 2148 289316 2150
rect 289372 2148 289386 2150
rect 288822 2128 289386 2148
rect 289556 480 289584 5646
rect 291936 5636 291988 5642
rect 291936 5578 291988 5584
rect 290740 5568 290792 5574
rect 290740 5510 290792 5516
rect 290752 480 290780 5510
rect 291948 480 291976 5578
rect 293144 480 293172 5646
rect 293696 5574 293724 8092
rect 294328 5772 294380 5778
rect 294328 5714 294380 5720
rect 293684 5568 293736 5574
rect 293684 5510 293736 5516
rect 294340 480 294368 5714
rect 294800 5642 294828 8092
rect 295524 5840 295576 5846
rect 295524 5782 295576 5788
rect 294788 5636 294840 5642
rect 294788 5578 294840 5584
rect 295536 480 295564 5782
rect 295996 5710 296024 8092
rect 297100 5778 297128 8092
rect 297088 5772 297140 5778
rect 297088 5714 297140 5720
rect 295984 5704 296036 5710
rect 295984 5646 296036 5652
rect 297916 5636 297968 5642
rect 297916 5578 297968 5584
rect 296628 5568 296680 5574
rect 296628 5510 296680 5516
rect 296640 4026 296668 5510
rect 296640 3998 296760 4026
rect 296732 480 296760 3998
rect 297928 480 297956 5578
rect 298296 5574 298324 8092
rect 299112 5704 299164 5710
rect 299112 5646 299164 5652
rect 298284 5568 298336 5574
rect 298284 5510 298336 5516
rect 299124 480 299152 5646
rect 299400 5642 299428 8092
rect 300308 5772 300360 5778
rect 300308 5714 300360 5720
rect 299388 5636 299440 5642
rect 299388 5578 299440 5584
rect 300320 480 300348 5714
rect 300596 5710 300624 8092
rect 300584 5704 300636 5710
rect 300584 5646 300636 5652
rect 301700 5642 301728 8092
rect 302896 5778 302924 8092
rect 302884 5772 302936 5778
rect 302884 5714 302936 5720
rect 303528 5704 303580 5710
rect 303528 5646 303580 5652
rect 301044 5636 301096 5642
rect 301044 5578 301096 5584
rect 301688 5636 301740 5642
rect 301688 5578 301740 5584
rect 301056 3534 301084 5578
rect 301412 5568 301464 5574
rect 301412 5510 301464 5516
rect 301044 3528 301096 3534
rect 301044 3470 301096 3476
rect 301424 480 301452 5510
rect 302608 3528 302660 3534
rect 302608 3470 302660 3476
rect 303540 3482 303568 5646
rect 304000 5574 304028 8092
rect 305104 5642 305132 8092
rect 306300 5846 306328 8092
rect 307404 6186 307432 8092
rect 307392 6180 307444 6186
rect 307392 6122 307444 6128
rect 306822 6012 307386 6032
rect 306822 6010 306836 6012
rect 306892 6010 306916 6012
rect 306972 6010 306996 6012
rect 307052 6010 307076 6012
rect 307132 6010 307156 6012
rect 307212 6010 307236 6012
rect 307292 6010 307316 6012
rect 307372 6010 307386 6012
rect 307066 5958 307076 6010
rect 307132 5958 307142 6010
rect 306822 5956 306836 5958
rect 306892 5956 306916 5958
rect 306972 5956 306996 5958
rect 307052 5956 307076 5958
rect 307132 5956 307156 5958
rect 307212 5956 307236 5958
rect 307292 5956 307316 5958
rect 307372 5956 307386 5958
rect 306822 5936 307386 5956
rect 306288 5840 306340 5846
rect 306288 5782 306340 5788
rect 307944 5840 307996 5846
rect 307944 5782 307996 5788
rect 306196 5772 306248 5778
rect 306196 5714 306248 5720
rect 304908 5636 304960 5642
rect 304908 5578 304960 5584
rect 305092 5636 305144 5642
rect 305092 5578 305144 5584
rect 303988 5568 304040 5574
rect 303988 5510 304040 5516
rect 304920 3482 304948 5578
rect 302620 480 302648 3470
rect 303540 3454 303844 3482
rect 304920 3454 305040 3482
rect 303816 480 303844 3454
rect 305012 480 305040 3454
rect 306208 480 306236 5714
rect 307484 5568 307536 5574
rect 307484 5510 307536 5516
rect 306822 4924 307386 4944
rect 306822 4922 306836 4924
rect 306892 4922 306916 4924
rect 306972 4922 306996 4924
rect 307052 4922 307076 4924
rect 307132 4922 307156 4924
rect 307212 4922 307236 4924
rect 307292 4922 307316 4924
rect 307372 4922 307386 4924
rect 307066 4870 307076 4922
rect 307132 4870 307142 4922
rect 306822 4868 306836 4870
rect 306892 4868 306916 4870
rect 306972 4868 306996 4870
rect 307052 4868 307076 4870
rect 307132 4868 307156 4870
rect 307212 4868 307236 4870
rect 307292 4868 307316 4870
rect 307372 4868 307386 4870
rect 306822 4848 307386 4868
rect 306822 3836 307386 3856
rect 306822 3834 306836 3836
rect 306892 3834 306916 3836
rect 306972 3834 306996 3836
rect 307052 3834 307076 3836
rect 307132 3834 307156 3836
rect 307212 3834 307236 3836
rect 307292 3834 307316 3836
rect 307372 3834 307386 3836
rect 307066 3782 307076 3834
rect 307132 3782 307142 3834
rect 306822 3780 306836 3782
rect 306892 3780 306916 3782
rect 306972 3780 306996 3782
rect 307052 3780 307076 3782
rect 307132 3780 307156 3782
rect 307212 3780 307236 3782
rect 307292 3780 307316 3782
rect 307372 3780 307386 3782
rect 306822 3760 307386 3780
rect 306822 2748 307386 2768
rect 306822 2746 306836 2748
rect 306892 2746 306916 2748
rect 306972 2746 306996 2748
rect 307052 2746 307076 2748
rect 307132 2746 307156 2748
rect 307212 2746 307236 2748
rect 307292 2746 307316 2748
rect 307372 2746 307386 2748
rect 307066 2694 307076 2746
rect 307132 2694 307142 2746
rect 306822 2692 306836 2694
rect 306892 2692 306916 2694
rect 306972 2692 306996 2694
rect 307052 2692 307076 2694
rect 307132 2692 307156 2694
rect 307212 2692 307236 2694
rect 307292 2692 307316 2694
rect 307372 2692 307386 2694
rect 306822 2672 307386 2692
rect 307496 2530 307524 5510
rect 307956 4078 307984 5782
rect 308600 5778 308628 8092
rect 309140 6180 309192 6186
rect 309140 6122 309192 6128
rect 308588 5772 308640 5778
rect 308588 5714 308640 5720
rect 308588 5636 308640 5642
rect 308588 5578 308640 5584
rect 307944 4072 307996 4078
rect 307944 4014 307996 4020
rect 307404 2502 307524 2530
rect 307404 480 307432 2502
rect 308600 480 308628 5578
rect 309152 3194 309180 6122
rect 309704 5574 309732 8092
rect 310900 5642 310928 8092
rect 311808 5772 311860 5778
rect 311808 5714 311860 5720
rect 310888 5636 310940 5642
rect 310888 5578 310940 5584
rect 309692 5568 309744 5574
rect 309692 5510 309744 5516
rect 309784 4072 309836 4078
rect 309784 4014 309836 4020
rect 309140 3188 309192 3194
rect 309140 3130 309192 3136
rect 309796 480 309824 4014
rect 311820 3482 311848 5714
rect 312004 5710 312032 8092
rect 313200 6390 313228 8092
rect 313188 6384 313240 6390
rect 313188 6326 313240 6332
rect 311992 5704 312044 5710
rect 311992 5646 312044 5652
rect 314304 5574 314332 8092
rect 314660 6384 314712 6390
rect 314660 6326 314712 6332
rect 314568 5636 314620 5642
rect 314568 5578 314620 5584
rect 313188 5568 313240 5574
rect 313188 5510 313240 5516
rect 314292 5568 314344 5574
rect 314292 5510 314344 5516
rect 313200 3482 313228 5510
rect 311820 3454 312216 3482
rect 313200 3454 313412 3482
rect 310980 3188 311032 3194
rect 310980 3130 311032 3136
rect 310992 480 311020 3130
rect 312188 480 312216 3454
rect 313384 480 313412 3454
rect 314580 480 314608 5578
rect 314672 4010 314700 6326
rect 315408 5642 315436 8092
rect 315764 5704 315816 5710
rect 315764 5646 315816 5652
rect 315396 5636 315448 5642
rect 315396 5578 315448 5584
rect 314660 4004 314712 4010
rect 314660 3946 314712 3952
rect 315776 480 315804 5646
rect 316604 5574 316632 8092
rect 317708 5778 317736 8092
rect 317696 5772 317748 5778
rect 317696 5714 317748 5720
rect 318904 5642 318932 8092
rect 320008 5710 320036 8092
rect 321204 5846 321232 8092
rect 322308 6186 322336 8092
rect 322296 6180 322348 6186
rect 322296 6122 322348 6128
rect 321192 5840 321244 5846
rect 321192 5782 321244 5788
rect 321468 5772 321520 5778
rect 321468 5714 321520 5720
rect 319996 5704 320048 5710
rect 319996 5646 320048 5652
rect 317696 5636 317748 5642
rect 317696 5578 317748 5584
rect 318892 5636 318944 5642
rect 318892 5578 318944 5584
rect 316500 5568 316552 5574
rect 316500 5510 316552 5516
rect 316592 5568 316644 5574
rect 316592 5510 316644 5516
rect 316512 3942 316540 5510
rect 316960 4004 317012 4010
rect 316960 3946 317012 3952
rect 316500 3936 316552 3942
rect 316500 3878 316552 3884
rect 316972 480 317000 3946
rect 317708 2854 317736 5578
rect 320088 5568 320140 5574
rect 320088 5510 320140 5516
rect 318064 3936 318116 3942
rect 318064 3878 318116 3884
rect 317696 2848 317748 2854
rect 317696 2790 317748 2796
rect 318076 480 318104 3878
rect 320100 3482 320128 5510
rect 321480 3482 321508 5714
rect 322020 5704 322072 5710
rect 322020 5646 322072 5652
rect 322032 3534 322060 5646
rect 322848 5636 322900 5642
rect 322848 5578 322900 5584
rect 322020 3528 322072 3534
rect 320100 3454 320496 3482
rect 321480 3454 321692 3482
rect 322020 3470 322072 3476
rect 319260 2848 319312 2854
rect 319260 2790 319312 2796
rect 319272 480 319300 2790
rect 320468 480 320496 3454
rect 321664 480 321692 3454
rect 322860 480 322888 5578
rect 323504 5574 323532 8092
rect 324320 6180 324372 6186
rect 324320 6122 324372 6128
rect 324136 5840 324188 5846
rect 324136 5782 324188 5788
rect 323492 5568 323544 5574
rect 323492 5510 323544 5516
rect 324148 3534 324176 5782
rect 324332 4078 324360 6122
rect 324608 5846 324636 8092
rect 324596 5840 324648 5846
rect 324596 5782 324648 5788
rect 325712 5642 325740 8092
rect 325700 5636 325752 5642
rect 325700 5578 325752 5584
rect 326908 5574 326936 8092
rect 327172 5840 327224 5846
rect 327172 5782 327224 5788
rect 326528 5568 326580 5574
rect 326528 5510 326580 5516
rect 326896 5568 326948 5574
rect 326896 5510 326948 5516
rect 324822 5468 325386 5488
rect 324822 5466 324836 5468
rect 324892 5466 324916 5468
rect 324972 5466 324996 5468
rect 325052 5466 325076 5468
rect 325132 5466 325156 5468
rect 325212 5466 325236 5468
rect 325292 5466 325316 5468
rect 325372 5466 325386 5468
rect 325066 5414 325076 5466
rect 325132 5414 325142 5466
rect 324822 5412 324836 5414
rect 324892 5412 324916 5414
rect 324972 5412 324996 5414
rect 325052 5412 325076 5414
rect 325132 5412 325156 5414
rect 325212 5412 325236 5414
rect 325292 5412 325316 5414
rect 325372 5412 325386 5414
rect 324822 5392 325386 5412
rect 324822 4380 325386 4400
rect 324822 4378 324836 4380
rect 324892 4378 324916 4380
rect 324972 4378 324996 4380
rect 325052 4378 325076 4380
rect 325132 4378 325156 4380
rect 325212 4378 325236 4380
rect 325292 4378 325316 4380
rect 325372 4378 325386 4380
rect 325066 4326 325076 4378
rect 325132 4326 325142 4378
rect 324822 4324 324836 4326
rect 324892 4324 324916 4326
rect 324972 4324 324996 4326
rect 325052 4324 325076 4326
rect 325132 4324 325156 4326
rect 325212 4324 325236 4326
rect 325292 4324 325316 4326
rect 325372 4324 325386 4326
rect 324822 4304 325386 4324
rect 324320 4072 324372 4078
rect 324320 4014 324372 4020
rect 326436 4072 326488 4078
rect 326436 4014 326488 4020
rect 324044 3528 324096 3534
rect 324044 3470 324096 3476
rect 324136 3528 324188 3534
rect 324136 3470 324188 3476
rect 325424 3528 325476 3534
rect 325424 3470 325476 3476
rect 324056 480 324084 3470
rect 324822 3292 325386 3312
rect 324822 3290 324836 3292
rect 324892 3290 324916 3292
rect 324972 3290 324996 3292
rect 325052 3290 325076 3292
rect 325132 3290 325156 3292
rect 325212 3290 325236 3292
rect 325292 3290 325316 3292
rect 325372 3290 325386 3292
rect 325066 3238 325076 3290
rect 325132 3238 325142 3290
rect 324822 3236 324836 3238
rect 324892 3236 324916 3238
rect 324972 3236 324996 3238
rect 325052 3236 325076 3238
rect 325132 3236 325156 3238
rect 325212 3236 325236 3238
rect 325292 3236 325316 3238
rect 325372 3236 325386 3238
rect 324822 3216 325386 3236
rect 324822 2204 325386 2224
rect 324822 2202 324836 2204
rect 324892 2202 324916 2204
rect 324972 2202 324996 2204
rect 325052 2202 325076 2204
rect 325132 2202 325156 2204
rect 325212 2202 325236 2204
rect 325292 2202 325316 2204
rect 325372 2202 325386 2204
rect 325066 2150 325076 2202
rect 325132 2150 325142 2202
rect 324822 2148 324836 2150
rect 324892 2148 324916 2150
rect 324972 2148 324996 2150
rect 325052 2148 325076 2150
rect 325132 2148 325156 2150
rect 325212 2148 325236 2150
rect 325292 2148 325316 2150
rect 325372 2148 325386 2150
rect 324822 2128 325386 2148
rect 325436 1986 325464 3470
rect 325252 1958 325464 1986
rect 325252 480 325280 1958
rect 326448 480 326476 4014
rect 326540 3058 326568 5510
rect 326528 3052 326580 3058
rect 326528 2994 326580 3000
rect 327184 2922 327212 5782
rect 328012 5710 328040 8092
rect 328000 5704 328052 5710
rect 328000 5646 328052 5652
rect 329208 5574 329236 8092
rect 330116 5704 330168 5710
rect 330116 5646 330168 5652
rect 329748 5636 329800 5642
rect 329748 5578 329800 5584
rect 329012 5568 329064 5574
rect 329012 5510 329064 5516
rect 329196 5568 329248 5574
rect 329196 5510 329248 5516
rect 329024 3466 329052 5510
rect 329760 3482 329788 5578
rect 329012 3460 329064 3466
rect 329760 3454 330064 3482
rect 329012 3402 329064 3408
rect 327632 3052 327684 3058
rect 327632 2994 327684 3000
rect 327172 2916 327224 2922
rect 327172 2858 327224 2864
rect 327644 480 327672 2994
rect 328828 2916 328880 2922
rect 328828 2858 328880 2864
rect 328840 480 328868 2858
rect 330036 480 330064 3454
rect 330128 3194 330156 5646
rect 330312 5642 330340 8092
rect 331508 5914 331536 8092
rect 331496 5908 331548 5914
rect 331496 5850 331548 5856
rect 332612 5778 332640 8092
rect 333808 5846 333836 8092
rect 333980 5908 334032 5914
rect 333980 5850 334032 5856
rect 333796 5840 333848 5846
rect 333796 5782 333848 5788
rect 332600 5772 332652 5778
rect 332600 5714 332652 5720
rect 330300 5636 330352 5642
rect 330300 5578 330352 5584
rect 332600 5636 332652 5642
rect 332600 5578 332652 5584
rect 331312 5568 331364 5574
rect 331312 5510 331364 5516
rect 331324 3534 331352 5510
rect 331312 3528 331364 3534
rect 331312 3470 331364 3476
rect 331220 3460 331272 3466
rect 331220 3402 331272 3408
rect 330116 3188 330168 3194
rect 330116 3130 330168 3136
rect 331232 480 331260 3402
rect 332612 3398 332640 5578
rect 333612 3528 333664 3534
rect 333612 3470 333664 3476
rect 332600 3392 332652 3398
rect 332600 3334 332652 3340
rect 332416 3188 332468 3194
rect 332416 3130 332468 3136
rect 332428 480 332456 3130
rect 333624 480 333652 3470
rect 333992 3466 334020 5850
rect 334912 5642 334940 8092
rect 335820 5772 335872 5778
rect 335820 5714 335872 5720
rect 334900 5636 334952 5642
rect 334900 5578 334952 5584
rect 335832 3942 335860 5714
rect 336108 5574 336136 8092
rect 336648 5840 336700 5846
rect 336648 5782 336700 5788
rect 336096 5568 336148 5574
rect 336096 5510 336148 5516
rect 335820 3936 335872 3942
rect 335820 3878 335872 3884
rect 333980 3460 334032 3466
rect 333980 3402 334032 3408
rect 335912 3460 335964 3466
rect 335912 3402 335964 3408
rect 334716 3392 334768 3398
rect 334716 3334 334768 3340
rect 334728 480 334756 3334
rect 335924 480 335952 3402
rect 336660 2990 336688 5782
rect 337212 5710 337240 8092
rect 338316 5778 338344 8092
rect 339512 5846 339540 8092
rect 340616 6390 340644 8092
rect 340604 6384 340656 6390
rect 340604 6326 340656 6332
rect 341812 6118 341840 8092
rect 342720 6384 342772 6390
rect 342720 6326 342772 6332
rect 341800 6112 341852 6118
rect 341800 6054 341852 6060
rect 339500 5840 339552 5846
rect 339500 5782 339552 5788
rect 342260 5840 342312 5846
rect 342260 5782 342312 5788
rect 338304 5772 338356 5778
rect 338304 5714 338356 5720
rect 340880 5772 340932 5778
rect 340880 5714 340932 5720
rect 337200 5704 337252 5710
rect 337200 5646 337252 5652
rect 339500 5704 339552 5710
rect 339500 5646 339552 5652
rect 337292 5636 337344 5642
rect 337292 5578 337344 5584
rect 337108 3936 337160 3942
rect 337108 3878 337160 3884
rect 336648 2984 336700 2990
rect 336648 2926 336700 2932
rect 337120 480 337148 3878
rect 337304 2922 337332 5578
rect 338304 5568 338356 5574
rect 338304 5510 338356 5516
rect 338316 3534 338344 5510
rect 338304 3528 338356 3534
rect 338304 3470 338356 3476
rect 339512 3398 339540 5646
rect 340696 3528 340748 3534
rect 340696 3470 340748 3476
rect 339500 3392 339552 3398
rect 339500 3334 339552 3340
rect 338304 2984 338356 2990
rect 338304 2926 338356 2932
rect 337292 2916 337344 2922
rect 337292 2858 337344 2864
rect 338316 480 338344 2926
rect 339500 2916 339552 2922
rect 339500 2858 339552 2864
rect 339512 480 339540 2858
rect 340708 480 340736 3470
rect 340892 3466 340920 5714
rect 342272 3534 342300 5782
rect 342732 3602 342760 6326
rect 342916 6186 342944 8092
rect 342904 6180 342956 6186
rect 342904 6122 342956 6128
rect 343640 6112 343692 6118
rect 343640 6054 343692 6060
rect 342822 6012 343386 6032
rect 342822 6010 342836 6012
rect 342892 6010 342916 6012
rect 342972 6010 342996 6012
rect 343052 6010 343076 6012
rect 343132 6010 343156 6012
rect 343212 6010 343236 6012
rect 343292 6010 343316 6012
rect 343372 6010 343386 6012
rect 343066 5958 343076 6010
rect 343132 5958 343142 6010
rect 342822 5956 342836 5958
rect 342892 5956 342916 5958
rect 342972 5956 342996 5958
rect 343052 5956 343076 5958
rect 343132 5956 343156 5958
rect 343212 5956 343236 5958
rect 343292 5956 343316 5958
rect 343372 5956 343386 5958
rect 342822 5936 343386 5956
rect 342822 4924 343386 4944
rect 342822 4922 342836 4924
rect 342892 4922 342916 4924
rect 342972 4922 342996 4924
rect 343052 4922 343076 4924
rect 343132 4922 343156 4924
rect 343212 4922 343236 4924
rect 343292 4922 343316 4924
rect 343372 4922 343386 4924
rect 343066 4870 343076 4922
rect 343132 4870 343142 4922
rect 342822 4868 342836 4870
rect 342892 4868 342916 4870
rect 342972 4868 342996 4870
rect 343052 4868 343076 4870
rect 343132 4868 343156 4870
rect 343212 4868 343236 4870
rect 343292 4868 343316 4870
rect 343372 4868 343386 4870
rect 342822 4848 343386 4868
rect 343652 4078 343680 6054
rect 344112 5574 344140 8092
rect 345216 5710 345244 8092
rect 346124 6180 346176 6186
rect 346124 6122 346176 6128
rect 345204 5704 345256 5710
rect 345204 5646 345256 5652
rect 344100 5568 344152 5574
rect 344100 5510 344152 5516
rect 343640 4072 343692 4078
rect 343640 4014 343692 4020
rect 342822 3836 343386 3856
rect 342822 3834 342836 3836
rect 342892 3834 342916 3836
rect 342972 3834 342996 3836
rect 343052 3834 343076 3836
rect 343132 3834 343156 3836
rect 343212 3834 343236 3836
rect 343292 3834 343316 3836
rect 343372 3834 343386 3836
rect 343066 3782 343076 3834
rect 343132 3782 343142 3834
rect 342822 3780 342836 3782
rect 342892 3780 342916 3782
rect 342972 3780 342996 3782
rect 343052 3780 343076 3782
rect 343132 3780 343156 3782
rect 343212 3780 343236 3782
rect 343292 3780 343316 3782
rect 343372 3780 343386 3782
rect 342822 3760 343386 3780
rect 342720 3596 342772 3602
rect 342720 3538 342772 3544
rect 345480 3596 345532 3602
rect 345480 3538 345532 3544
rect 342260 3528 342312 3534
rect 342260 3470 342312 3476
rect 344284 3528 344336 3534
rect 344284 3470 344336 3476
rect 340880 3460 340932 3466
rect 340880 3402 340932 3408
rect 342720 3460 342772 3466
rect 342720 3402 342772 3408
rect 341892 3392 341944 3398
rect 341892 3334 341944 3340
rect 341904 480 341932 3334
rect 342732 2530 342760 3402
rect 342822 2748 343386 2768
rect 342822 2746 342836 2748
rect 342892 2746 342916 2748
rect 342972 2746 342996 2748
rect 343052 2746 343076 2748
rect 343132 2746 343156 2748
rect 343212 2746 343236 2748
rect 343292 2746 343316 2748
rect 343372 2746 343386 2748
rect 343066 2694 343076 2746
rect 343132 2694 343142 2746
rect 342822 2692 342836 2694
rect 342892 2692 342916 2694
rect 342972 2692 342996 2694
rect 343052 2692 343076 2694
rect 343132 2692 343156 2694
rect 343212 2692 343236 2694
rect 343292 2692 343316 2694
rect 343372 2692 343386 2694
rect 342822 2672 343386 2692
rect 342732 2502 343128 2530
rect 343100 480 343128 2502
rect 344296 480 344324 3470
rect 345492 480 345520 3538
rect 346136 3126 346164 6122
rect 346412 5642 346440 8092
rect 346400 5636 346452 5642
rect 346400 5578 346452 5584
rect 347516 5574 347544 8092
rect 348620 5710 348648 8092
rect 349816 5846 349844 8092
rect 350920 6118 350948 8092
rect 350908 6112 350960 6118
rect 350908 6054 350960 6060
rect 349804 5840 349856 5846
rect 349804 5782 349856 5788
rect 347780 5704 347832 5710
rect 347780 5646 347832 5652
rect 348608 5704 348660 5710
rect 348608 5646 348660 5652
rect 351092 5704 351144 5710
rect 351092 5646 351144 5652
rect 346860 5568 346912 5574
rect 346860 5510 346912 5516
rect 347504 5568 347556 5574
rect 347504 5510 347556 5516
rect 346676 4072 346728 4078
rect 346676 4014 346728 4020
rect 346124 3120 346176 3126
rect 346124 3062 346176 3068
rect 346688 480 346716 4014
rect 346872 2854 346900 5510
rect 347792 3602 347820 5646
rect 349160 5636 349212 5642
rect 349160 5578 349212 5584
rect 347780 3596 347832 3602
rect 347780 3538 347832 3544
rect 349172 3534 349200 5578
rect 349988 5568 350040 5574
rect 349988 5510 350040 5516
rect 349160 3528 349212 3534
rect 349160 3470 349212 3476
rect 350000 3194 350028 5510
rect 350264 3596 350316 3602
rect 350264 3538 350316 3544
rect 349988 3188 350040 3194
rect 349988 3130 350040 3136
rect 347872 3120 347924 3126
rect 347872 3062 347924 3068
rect 346860 2848 346912 2854
rect 346860 2790 346912 2796
rect 347884 480 347912 3062
rect 349068 2848 349120 2854
rect 349068 2790 349120 2796
rect 349080 480 349108 2790
rect 350276 480 350304 3538
rect 351104 3126 351132 5646
rect 352116 5642 352144 8092
rect 353220 5846 353248 8092
rect 353300 6112 353352 6118
rect 353300 6054 353352 6060
rect 352288 5840 352340 5846
rect 352288 5782 352340 5788
rect 353208 5840 353260 5846
rect 353208 5782 353260 5788
rect 352104 5636 352156 5642
rect 352104 5578 352156 5584
rect 352300 4078 352328 5782
rect 352288 4072 352340 4078
rect 352288 4014 352340 4020
rect 353312 3738 353340 6054
rect 354416 5710 354444 8092
rect 355520 6118 355548 8092
rect 355508 6112 355560 6118
rect 355508 6054 355560 6060
rect 355508 5840 355560 5846
rect 355508 5782 355560 5788
rect 354404 5704 354456 5710
rect 354404 5646 354456 5652
rect 355520 4146 355548 5782
rect 355600 5636 355652 5642
rect 355600 5578 355652 5584
rect 355508 4140 355560 4146
rect 355508 4082 355560 4088
rect 354956 4072 355008 4078
rect 354956 4014 355008 4020
rect 353300 3732 353352 3738
rect 353300 3674 353352 3680
rect 351368 3528 351420 3534
rect 351368 3470 351420 3476
rect 351092 3120 351144 3126
rect 351092 3062 351144 3068
rect 351380 480 351408 3470
rect 352564 3188 352616 3194
rect 352564 3130 352616 3136
rect 352576 480 352604 3130
rect 353760 3120 353812 3126
rect 353760 3062 353812 3068
rect 353772 480 353800 3062
rect 354968 480 354996 4014
rect 355612 2854 355640 5578
rect 356716 5574 356744 8092
rect 357256 5704 357308 5710
rect 357256 5646 357308 5652
rect 356704 5568 356756 5574
rect 356704 5510 356756 5516
rect 356152 3732 356204 3738
rect 356152 3674 356204 3680
rect 355600 2848 355652 2854
rect 355600 2790 355652 2796
rect 356164 480 356192 3674
rect 357268 2922 357296 5646
rect 357820 5642 357848 8092
rect 358176 6112 358228 6118
rect 358176 6054 358228 6060
rect 357808 5636 357860 5642
rect 357808 5578 357860 5584
rect 358188 3602 358216 6054
rect 358924 5710 358952 8092
rect 360120 6118 360148 8092
rect 361224 6254 361252 8092
rect 361212 6248 361264 6254
rect 361212 6190 361264 6196
rect 360108 6112 360160 6118
rect 360108 6054 360160 6060
rect 362224 6112 362276 6118
rect 362224 6054 362276 6060
rect 358912 5704 358964 5710
rect 358912 5646 358964 5652
rect 361580 5704 361632 5710
rect 361580 5646 361632 5652
rect 360568 5636 360620 5642
rect 360568 5578 360620 5584
rect 359372 5568 359424 5574
rect 359372 5510 359424 5516
rect 358544 4140 358596 4146
rect 358544 4082 358596 4088
rect 358176 3596 358228 3602
rect 358176 3538 358228 3544
rect 357256 2916 357308 2922
rect 357256 2858 357308 2864
rect 357348 2848 357400 2854
rect 357348 2790 357400 2796
rect 357360 480 357388 2790
rect 358556 480 358584 4082
rect 359384 3534 359412 5510
rect 359372 3528 359424 3534
rect 359372 3470 359424 3476
rect 360580 3466 360608 5578
rect 360822 5468 361386 5488
rect 360822 5466 360836 5468
rect 360892 5466 360916 5468
rect 360972 5466 360996 5468
rect 361052 5466 361076 5468
rect 361132 5466 361156 5468
rect 361212 5466 361236 5468
rect 361292 5466 361316 5468
rect 361372 5466 361386 5468
rect 361066 5414 361076 5466
rect 361132 5414 361142 5466
rect 360822 5412 360836 5414
rect 360892 5412 360916 5414
rect 360972 5412 360996 5414
rect 361052 5412 361076 5414
rect 361132 5412 361156 5414
rect 361212 5412 361236 5414
rect 361292 5412 361316 5414
rect 361372 5412 361386 5414
rect 360822 5392 361386 5412
rect 360822 4380 361386 4400
rect 360822 4378 360836 4380
rect 360892 4378 360916 4380
rect 360972 4378 360996 4380
rect 361052 4378 361076 4380
rect 361132 4378 361156 4380
rect 361212 4378 361236 4380
rect 361292 4378 361316 4380
rect 361372 4378 361386 4380
rect 361066 4326 361076 4378
rect 361132 4326 361142 4378
rect 360822 4324 360836 4326
rect 360892 4324 360916 4326
rect 360972 4324 360996 4326
rect 361052 4324 361076 4326
rect 361132 4324 361156 4326
rect 361212 4324 361236 4326
rect 361292 4324 361316 4326
rect 361372 4324 361386 4326
rect 360822 4304 361386 4324
rect 361592 3942 361620 5646
rect 361580 3936 361632 3942
rect 361580 3878 361632 3884
rect 362236 3602 362264 6054
rect 362420 5574 362448 8092
rect 362960 6248 363012 6254
rect 362960 6190 363012 6196
rect 362408 5568 362460 5574
rect 362408 5510 362460 5516
rect 362972 4078 363000 6190
rect 363524 5710 363552 8092
rect 363512 5704 363564 5710
rect 363512 5646 363564 5652
rect 364720 5642 364748 8092
rect 365824 5778 365852 8092
rect 365812 5772 365864 5778
rect 365812 5714 365864 5720
rect 366548 5704 366600 5710
rect 366548 5646 366600 5652
rect 364708 5636 364760 5642
rect 364708 5578 364760 5584
rect 365628 5568 365680 5574
rect 365628 5510 365680 5516
rect 362960 4072 363012 4078
rect 362960 4014 363012 4020
rect 364524 3936 364576 3942
rect 364524 3878 364576 3884
rect 360752 3596 360804 3602
rect 360752 3538 360804 3544
rect 362224 3596 362276 3602
rect 362224 3538 362276 3544
rect 360568 3460 360620 3466
rect 360568 3402 360620 3408
rect 359740 2916 359792 2922
rect 359740 2858 359792 2864
rect 359752 480 359780 2858
rect 360764 1986 360792 3538
rect 362132 3528 362184 3534
rect 362132 3470 362184 3476
rect 360822 3292 361386 3312
rect 360822 3290 360836 3292
rect 360892 3290 360916 3292
rect 360972 3290 360996 3292
rect 361052 3290 361076 3292
rect 361132 3290 361156 3292
rect 361212 3290 361236 3292
rect 361292 3290 361316 3292
rect 361372 3290 361386 3292
rect 361066 3238 361076 3290
rect 361132 3238 361142 3290
rect 360822 3236 360836 3238
rect 360892 3236 360916 3238
rect 360972 3236 360996 3238
rect 361052 3236 361076 3238
rect 361132 3236 361156 3238
rect 361212 3236 361236 3238
rect 361292 3236 361316 3238
rect 361372 3236 361386 3238
rect 360822 3216 361386 3236
rect 360822 2204 361386 2224
rect 360822 2202 360836 2204
rect 360892 2202 360916 2204
rect 360972 2202 360996 2204
rect 361052 2202 361076 2204
rect 361132 2202 361156 2204
rect 361212 2202 361236 2204
rect 361292 2202 361316 2204
rect 361372 2202 361386 2204
rect 361066 2150 361076 2202
rect 361132 2150 361142 2202
rect 360822 2148 360836 2150
rect 360892 2148 360916 2150
rect 360972 2148 360996 2150
rect 361052 2148 361076 2150
rect 361132 2148 361156 2150
rect 361212 2148 361236 2150
rect 361292 2148 361316 2150
rect 361372 2148 361386 2150
rect 360822 2128 361386 2148
rect 360764 1958 360976 1986
rect 360948 480 360976 1958
rect 362144 480 362172 3470
rect 363328 3460 363380 3466
rect 363328 3402 363380 3408
rect 363340 480 363368 3402
rect 364536 480 364564 3878
rect 365640 3058 365668 5510
rect 366560 4146 366588 5646
rect 367020 5574 367048 8092
rect 368124 5846 368152 8092
rect 369228 6118 369256 8092
rect 370424 6390 370452 8092
rect 370412 6384 370464 6390
rect 370412 6326 370464 6332
rect 369216 6112 369268 6118
rect 369216 6054 369268 6060
rect 368112 5840 368164 5846
rect 368112 5782 368164 5788
rect 371056 5840 371108 5846
rect 371056 5782 371108 5788
rect 368664 5772 368716 5778
rect 368664 5714 368716 5720
rect 367468 5636 367520 5642
rect 367468 5578 367520 5584
rect 367008 5568 367060 5574
rect 367008 5510 367060 5516
rect 366548 4140 366600 4146
rect 366548 4082 366600 4088
rect 366916 4072 366968 4078
rect 366916 4014 366968 4020
rect 365720 3596 365772 3602
rect 365720 3538 365772 3544
rect 365628 3052 365680 3058
rect 365628 2994 365680 3000
rect 365732 480 365760 3538
rect 366928 480 366956 4014
rect 367480 3534 367508 5578
rect 367468 3528 367520 3534
rect 367468 3470 367520 3476
rect 368676 3194 368704 5714
rect 369768 5568 369820 5574
rect 369768 5510 369820 5516
rect 369216 4140 369268 4146
rect 369216 4082 369268 4088
rect 368664 3188 368716 3194
rect 368664 3130 368716 3136
rect 368020 3052 368072 3058
rect 368020 2994 368072 3000
rect 368032 480 368060 2994
rect 369228 480 369256 4082
rect 369780 3602 369808 5510
rect 371068 4078 371096 5782
rect 371528 5574 371556 8092
rect 372620 6384 372672 6390
rect 372620 6326 372672 6332
rect 371608 6112 371660 6118
rect 371608 6054 371660 6060
rect 371516 5568 371568 5574
rect 371516 5510 371568 5516
rect 371620 4146 371648 6054
rect 371608 4140 371660 4146
rect 371608 4082 371660 4088
rect 371056 4072 371108 4078
rect 371056 4014 371108 4020
rect 369768 3596 369820 3602
rect 369768 3538 369820 3544
rect 370412 3528 370464 3534
rect 370412 3470 370464 3476
rect 370424 480 370452 3470
rect 372632 3466 372660 6326
rect 372724 5710 372752 8092
rect 373828 5846 373856 8092
rect 373816 5840 373868 5846
rect 373816 5782 373868 5788
rect 372712 5704 372764 5710
rect 372712 5646 372764 5652
rect 375024 5574 375052 8092
rect 376128 5710 376156 8092
rect 376668 5840 376720 5846
rect 376668 5782 376720 5788
rect 375840 5704 375892 5710
rect 375840 5646 375892 5652
rect 376116 5704 376168 5710
rect 376116 5646 376168 5652
rect 374736 5568 374788 5574
rect 374736 5510 374788 5516
rect 375012 5568 375064 5574
rect 375012 5510 375064 5516
rect 374000 4072 374052 4078
rect 374000 4014 374052 4020
rect 372804 3596 372856 3602
rect 372804 3538 372856 3544
rect 372620 3460 372672 3466
rect 372620 3402 372672 3408
rect 371608 3188 371660 3194
rect 371608 3130 371660 3136
rect 371620 480 371648 3130
rect 372816 480 372844 3538
rect 374012 480 374040 4014
rect 374748 3738 374776 5510
rect 375852 4146 375880 5646
rect 375196 4140 375248 4146
rect 375196 4082 375248 4088
rect 375840 4140 375892 4146
rect 375840 4082 375892 4088
rect 374736 3732 374788 3738
rect 374736 3674 374788 3680
rect 375208 480 375236 4082
rect 376392 3460 376444 3466
rect 376392 3402 376444 3408
rect 376404 480 376432 3402
rect 376680 3194 376708 5782
rect 377324 5642 377352 8092
rect 377312 5636 377364 5642
rect 377312 5578 377364 5584
rect 378428 5574 378456 8092
rect 379624 6390 379652 8092
rect 379612 6384 379664 6390
rect 379612 6326 379664 6332
rect 378822 6012 379386 6032
rect 378822 6010 378836 6012
rect 378892 6010 378916 6012
rect 378972 6010 378996 6012
rect 379052 6010 379076 6012
rect 379132 6010 379156 6012
rect 379212 6010 379236 6012
rect 379292 6010 379316 6012
rect 379372 6010 379386 6012
rect 379066 5958 379076 6010
rect 379132 5958 379142 6010
rect 378822 5956 378836 5958
rect 378892 5956 378916 5958
rect 378972 5956 378996 5958
rect 379052 5956 379076 5958
rect 379132 5956 379156 5958
rect 379212 5956 379236 5958
rect 379292 5956 379316 5958
rect 379372 5956 379386 5958
rect 378822 5936 379386 5956
rect 380728 5846 380756 8092
rect 380716 5840 380768 5846
rect 380716 5782 380768 5788
rect 379428 5704 379480 5710
rect 379428 5646 379480 5652
rect 378048 5568 378100 5574
rect 378048 5510 378100 5516
rect 378416 5568 378468 5574
rect 378416 5510 378468 5516
rect 377588 3732 377640 3738
rect 377588 3674 377640 3680
rect 376668 3188 376720 3194
rect 376668 3130 376720 3136
rect 377600 480 377628 3674
rect 378060 3534 378088 5510
rect 378822 4924 379386 4944
rect 378822 4922 378836 4924
rect 378892 4922 378916 4924
rect 378972 4922 378996 4924
rect 379052 4922 379076 4924
rect 379132 4922 379156 4924
rect 379212 4922 379236 4924
rect 379292 4922 379316 4924
rect 379372 4922 379386 4924
rect 379066 4870 379076 4922
rect 379132 4870 379142 4922
rect 378822 4868 378836 4870
rect 378892 4868 378916 4870
rect 378972 4868 378996 4870
rect 379052 4868 379076 4870
rect 379132 4868 379156 4870
rect 379212 4868 379236 4870
rect 379292 4868 379316 4870
rect 379372 4868 379386 4870
rect 378822 4848 379386 4868
rect 378692 4140 378744 4146
rect 378692 4082 378744 4088
rect 378048 3528 378100 3534
rect 378048 3470 378100 3476
rect 378704 2530 378732 4082
rect 378822 3836 379386 3856
rect 378822 3834 378836 3836
rect 378892 3834 378916 3836
rect 378972 3834 378996 3836
rect 379052 3834 379076 3836
rect 379132 3834 379156 3836
rect 379212 3834 379236 3836
rect 379292 3834 379316 3836
rect 379372 3834 379386 3836
rect 379066 3782 379076 3834
rect 379132 3782 379142 3834
rect 378822 3780 378836 3782
rect 378892 3780 378916 3782
rect 378972 3780 378996 3782
rect 379052 3780 379076 3782
rect 379132 3780 379156 3782
rect 379212 3780 379236 3782
rect 379292 3780 379316 3782
rect 379372 3780 379386 3782
rect 378822 3760 379386 3780
rect 379440 3602 379468 5646
rect 380440 5636 380492 5642
rect 380440 5578 380492 5584
rect 379428 3596 379480 3602
rect 379428 3538 379480 3544
rect 380452 3466 380480 5578
rect 381832 5574 381860 8092
rect 382372 6384 382424 6390
rect 382372 6326 382424 6332
rect 382280 5840 382332 5846
rect 382280 5782 382332 5788
rect 380900 5568 380952 5574
rect 380900 5510 380952 5516
rect 381820 5568 381872 5574
rect 381820 5510 381872 5516
rect 380912 4146 380940 5510
rect 380900 4140 380952 4146
rect 380900 4082 380952 4088
rect 382292 3534 382320 5782
rect 382384 4078 382412 6326
rect 383028 5846 383056 8092
rect 383016 5840 383068 5846
rect 383016 5782 383068 5788
rect 384132 5642 384160 8092
rect 384120 5636 384172 5642
rect 384120 5578 384172 5584
rect 385328 5574 385356 8092
rect 386144 5840 386196 5846
rect 386144 5782 386196 5788
rect 384948 5568 385000 5574
rect 384948 5510 385000 5516
rect 385316 5568 385368 5574
rect 385316 5510 385368 5516
rect 384672 4140 384724 4146
rect 384672 4082 384724 4088
rect 382372 4072 382424 4078
rect 382372 4014 382424 4020
rect 382372 3596 382424 3602
rect 382372 3538 382424 3544
rect 381176 3528 381228 3534
rect 381176 3470 381228 3476
rect 382280 3528 382332 3534
rect 382280 3470 382332 3476
rect 380440 3460 380492 3466
rect 380440 3402 380492 3408
rect 379980 3188 380032 3194
rect 379980 3130 380032 3136
rect 378822 2748 379386 2768
rect 378822 2746 378836 2748
rect 378892 2746 378916 2748
rect 378972 2746 378996 2748
rect 379052 2746 379076 2748
rect 379132 2746 379156 2748
rect 379212 2746 379236 2748
rect 379292 2746 379316 2748
rect 379372 2746 379386 2748
rect 379066 2694 379076 2746
rect 379132 2694 379142 2746
rect 378822 2692 378836 2694
rect 378892 2692 378916 2694
rect 378972 2692 378996 2694
rect 379052 2692 379076 2694
rect 379132 2692 379156 2694
rect 379212 2692 379236 2694
rect 379292 2692 379316 2694
rect 379372 2692 379386 2694
rect 378822 2672 379386 2692
rect 378704 2502 378824 2530
rect 378796 480 378824 2502
rect 379992 480 380020 3130
rect 381188 480 381216 3470
rect 382384 480 382412 3538
rect 383568 3460 383620 3466
rect 383568 3402 383620 3408
rect 383580 480 383608 3402
rect 384684 480 384712 4082
rect 384960 3738 384988 5510
rect 385868 4072 385920 4078
rect 385868 4014 385920 4020
rect 384948 3732 385000 3738
rect 384948 3674 385000 3680
rect 385880 480 385908 4014
rect 386156 3058 386184 5782
rect 386432 5710 386460 8092
rect 387628 5846 387656 8092
rect 388732 6118 388760 8092
rect 388720 6112 388772 6118
rect 388720 6054 388772 6060
rect 387616 5840 387668 5846
rect 387616 5782 387668 5788
rect 389180 5840 389232 5846
rect 389180 5782 389232 5788
rect 386420 5704 386472 5710
rect 386420 5646 386472 5652
rect 387340 5636 387392 5642
rect 387340 5578 387392 5584
rect 387352 3534 387380 5578
rect 388536 5568 388588 5574
rect 388536 5510 388588 5516
rect 388260 3732 388312 3738
rect 388260 3674 388312 3680
rect 387064 3528 387116 3534
rect 387064 3470 387116 3476
rect 387340 3528 387392 3534
rect 387340 3470 387392 3476
rect 386144 3052 386196 3058
rect 386144 2994 386196 3000
rect 387076 480 387104 3470
rect 388272 480 388300 3674
rect 388548 3466 388576 5510
rect 389192 3602 389220 5782
rect 389640 5704 389692 5710
rect 389640 5646 389692 5652
rect 389180 3596 389232 3602
rect 389180 3538 389232 3544
rect 388536 3460 388588 3466
rect 388536 3402 388588 3408
rect 389652 3398 389680 5646
rect 389928 5642 389956 8092
rect 389916 5636 389968 5642
rect 389916 5578 389968 5584
rect 391032 5574 391060 8092
rect 391112 6112 391164 6118
rect 391112 6054 391164 6060
rect 391020 5568 391072 5574
rect 391020 5510 391072 5516
rect 391124 4146 391152 6054
rect 392136 5846 392164 8092
rect 392124 5840 392176 5846
rect 392124 5782 392176 5788
rect 393332 5642 393360 8092
rect 391940 5636 391992 5642
rect 391940 5578 391992 5584
rect 393320 5636 393372 5642
rect 393320 5578 393372 5584
rect 391112 4140 391164 4146
rect 391112 4082 391164 4088
rect 391952 3534 391980 5578
rect 394436 5574 394464 8092
rect 395344 5840 395396 5846
rect 395344 5782 395396 5788
rect 393596 5568 393648 5574
rect 393596 5510 393648 5516
rect 394424 5568 394476 5574
rect 394424 5510 394476 5516
rect 393608 4078 393636 5510
rect 393596 4072 393648 4078
rect 393596 4014 393648 4020
rect 394240 3596 394292 3602
rect 394240 3538 394292 3544
rect 390652 3528 390704 3534
rect 390652 3470 390704 3476
rect 391940 3528 391992 3534
rect 391940 3470 391992 3476
rect 389640 3392 389692 3398
rect 389640 3334 389692 3340
rect 389456 3052 389508 3058
rect 389456 2994 389508 3000
rect 389468 480 389496 2994
rect 390664 480 390692 3470
rect 391848 3460 391900 3466
rect 391848 3402 391900 3408
rect 391860 480 391888 3402
rect 393044 3392 393096 3398
rect 393044 3334 393096 3340
rect 393056 480 393084 3334
rect 394252 480 394280 3538
rect 395356 2922 395384 5782
rect 395632 5710 395660 8092
rect 396736 5846 396764 8092
rect 396724 5840 396776 5846
rect 396724 5782 396776 5788
rect 395620 5704 395672 5710
rect 395620 5646 395672 5652
rect 397932 5642 397960 8092
rect 399036 5778 399064 8092
rect 399852 5840 399904 5846
rect 399852 5782 399904 5788
rect 399024 5772 399076 5778
rect 399024 5714 399076 5720
rect 398748 5704 398800 5710
rect 398748 5646 398800 5652
rect 396540 5636 396592 5642
rect 396540 5578 396592 5584
rect 397920 5636 397972 5642
rect 397920 5578 397972 5584
rect 395436 4140 395488 4146
rect 395436 4082 395488 4088
rect 395344 2916 395396 2922
rect 395344 2858 395396 2864
rect 395448 480 395476 4082
rect 396552 3602 396580 5578
rect 396724 5568 396776 5574
rect 396724 5510 396776 5516
rect 396540 3596 396592 3602
rect 396540 3538 396592 3544
rect 396632 3528 396684 3534
rect 396632 3470 396684 3476
rect 396644 480 396672 3470
rect 396736 3466 396764 5510
rect 396822 5468 397386 5488
rect 396822 5466 396836 5468
rect 396892 5466 396916 5468
rect 396972 5466 396996 5468
rect 397052 5466 397076 5468
rect 397132 5466 397156 5468
rect 397212 5466 397236 5468
rect 397292 5466 397316 5468
rect 397372 5466 397386 5468
rect 397066 5414 397076 5466
rect 397132 5414 397142 5466
rect 396822 5412 396836 5414
rect 396892 5412 396916 5414
rect 396972 5412 396996 5414
rect 397052 5412 397076 5414
rect 397132 5412 397156 5414
rect 397212 5412 397236 5414
rect 397292 5412 397316 5414
rect 397372 5412 397386 5414
rect 396822 5392 397386 5412
rect 396822 4380 397386 4400
rect 396822 4378 396836 4380
rect 396892 4378 396916 4380
rect 396972 4378 396996 4380
rect 397052 4378 397076 4380
rect 397132 4378 397156 4380
rect 397212 4378 397236 4380
rect 397292 4378 397316 4380
rect 397372 4378 397386 4380
rect 397066 4326 397076 4378
rect 397132 4326 397142 4378
rect 396822 4324 396836 4326
rect 396892 4324 396916 4326
rect 396972 4324 396996 4326
rect 397052 4324 397076 4326
rect 397132 4324 397156 4326
rect 397212 4324 397236 4326
rect 397292 4324 397316 4326
rect 397372 4324 397386 4326
rect 396822 4304 397386 4324
rect 397828 4072 397880 4078
rect 397828 4014 397880 4020
rect 396724 3460 396776 3466
rect 396724 3402 396776 3408
rect 396822 3292 397386 3312
rect 396822 3290 396836 3292
rect 396892 3290 396916 3292
rect 396972 3290 396996 3292
rect 397052 3290 397076 3292
rect 397132 3290 397156 3292
rect 397212 3290 397236 3292
rect 397292 3290 397316 3292
rect 397372 3290 397386 3292
rect 397066 3238 397076 3290
rect 397132 3238 397142 3290
rect 396822 3236 396836 3238
rect 396892 3236 396916 3238
rect 396972 3236 396996 3238
rect 397052 3236 397076 3238
rect 397132 3236 397156 3238
rect 397212 3236 397236 3238
rect 397292 3236 397316 3238
rect 397372 3236 397386 3238
rect 396822 3216 397386 3236
rect 396822 2204 397386 2224
rect 396822 2202 396836 2204
rect 396892 2202 396916 2204
rect 396972 2202 396996 2204
rect 397052 2202 397076 2204
rect 397132 2202 397156 2204
rect 397212 2202 397236 2204
rect 397292 2202 397316 2204
rect 397372 2202 397386 2204
rect 397066 2150 397076 2202
rect 397132 2150 397142 2202
rect 396822 2148 396836 2150
rect 396892 2148 396916 2150
rect 396972 2148 396996 2150
rect 397052 2148 397076 2150
rect 397132 2148 397156 2150
rect 397212 2148 397236 2150
rect 397292 2148 397316 2150
rect 397372 2148 397386 2150
rect 396822 2128 397386 2148
rect 397840 480 397868 4014
rect 398760 3534 398788 5646
rect 399864 4010 399892 5782
rect 400232 5574 400260 8092
rect 401336 5846 401364 8092
rect 402440 5914 402468 8092
rect 402428 5908 402480 5914
rect 402428 5850 402480 5856
rect 401324 5840 401376 5846
rect 401324 5782 401376 5788
rect 401600 5772 401652 5778
rect 401600 5714 401652 5720
rect 400496 5636 400548 5642
rect 400496 5578 400548 5584
rect 400220 5568 400272 5574
rect 400220 5510 400272 5516
rect 400508 4078 400536 5578
rect 400496 4072 400548 4078
rect 400496 4014 400548 4020
rect 399852 4004 399904 4010
rect 399852 3946 399904 3952
rect 401612 3670 401640 5714
rect 403636 5642 403664 8092
rect 403900 5840 403952 5846
rect 403900 5782 403952 5788
rect 403624 5636 403676 5642
rect 403624 5578 403676 5584
rect 403716 4004 403768 4010
rect 403716 3946 403768 3952
rect 401600 3664 401652 3670
rect 401600 3606 401652 3612
rect 400220 3596 400272 3602
rect 400220 3538 400272 3544
rect 398748 3528 398800 3534
rect 398748 3470 398800 3476
rect 399024 2916 399076 2922
rect 399024 2858 399076 2864
rect 399036 480 399064 2858
rect 400232 480 400260 3538
rect 402520 3528 402572 3534
rect 402520 3470 402572 3476
rect 401324 3460 401376 3466
rect 401324 3402 401376 3408
rect 401336 480 401364 3402
rect 402532 480 402560 3470
rect 403728 480 403756 3946
rect 403912 3738 403940 5782
rect 404740 5574 404768 8092
rect 405648 5908 405700 5914
rect 405648 5850 405700 5856
rect 404084 5568 404136 5574
rect 404084 5510 404136 5516
rect 404728 5568 404780 5574
rect 404728 5510 404780 5516
rect 404096 4146 404124 5510
rect 404084 4140 404136 4146
rect 404084 4082 404136 4088
rect 404912 4072 404964 4078
rect 404912 4014 404964 4020
rect 403900 3732 403952 3738
rect 403900 3674 403952 3680
rect 404924 480 404952 4014
rect 405660 3194 405688 5850
rect 405936 5710 405964 8092
rect 407040 6526 407068 8092
rect 407028 6520 407080 6526
rect 407028 6462 407080 6468
rect 408236 5846 408264 8092
rect 408500 6520 408552 6526
rect 408500 6462 408552 6468
rect 408224 5840 408276 5846
rect 408224 5782 408276 5788
rect 405924 5704 405976 5710
rect 405924 5646 405976 5652
rect 407028 5636 407080 5642
rect 407028 5578 407080 5584
rect 406108 3664 406160 3670
rect 406108 3606 406160 3612
rect 405648 3188 405700 3194
rect 405648 3130 405700 3136
rect 406120 480 406148 3606
rect 407040 3466 407068 5578
rect 408408 5568 408460 5574
rect 408408 5510 408460 5516
rect 407304 4140 407356 4146
rect 407304 4082 407356 4088
rect 407028 3460 407080 3466
rect 407028 3402 407080 3408
rect 407316 480 407344 4082
rect 408420 3602 408448 5510
rect 408512 4146 408540 6462
rect 409340 5642 409368 8092
rect 410536 5914 410564 8092
rect 410524 5908 410576 5914
rect 410524 5850 410576 5856
rect 410432 5840 410484 5846
rect 410432 5782 410484 5788
rect 409420 5704 409472 5710
rect 409420 5646 409472 5652
rect 409328 5636 409380 5642
rect 409328 5578 409380 5584
rect 408500 4140 408552 4146
rect 408500 4082 408552 4088
rect 409432 4078 409460 5646
rect 409420 4072 409472 4078
rect 409420 4014 409472 4020
rect 408500 3732 408552 3738
rect 408500 3674 408552 3680
rect 408408 3596 408460 3602
rect 408408 3538 408460 3544
rect 408512 480 408540 3674
rect 410444 3534 410472 5782
rect 411260 5636 411312 5642
rect 411260 5578 411312 5584
rect 410432 3528 410484 3534
rect 410432 3470 410484 3476
rect 411272 3466 411300 5578
rect 411640 5574 411668 8092
rect 412744 5642 412772 8092
rect 413744 5908 413796 5914
rect 413744 5850 413796 5856
rect 412732 5636 412784 5642
rect 412732 5578 412784 5584
rect 411628 5568 411680 5574
rect 411628 5510 411680 5516
rect 413284 4072 413336 4078
rect 413284 4014 413336 4020
rect 412088 3596 412140 3602
rect 412088 3538 412140 3544
rect 410892 3460 410944 3466
rect 410892 3402 410944 3408
rect 411260 3460 411312 3466
rect 411260 3402 411312 3408
rect 409696 3188 409748 3194
rect 409696 3130 409748 3136
rect 409708 480 409736 3130
rect 410904 480 410932 3402
rect 412100 480 412128 3538
rect 413296 480 413324 4014
rect 413756 3058 413784 5850
rect 413940 5710 413968 8092
rect 415044 6254 415072 8092
rect 416240 6390 416268 8092
rect 416228 6384 416280 6390
rect 416228 6326 416280 6332
rect 415032 6248 415084 6254
rect 415032 6190 415084 6196
rect 416964 6248 417016 6254
rect 416964 6190 417016 6196
rect 414822 6012 415386 6032
rect 414822 6010 414836 6012
rect 414892 6010 414916 6012
rect 414972 6010 414996 6012
rect 415052 6010 415076 6012
rect 415132 6010 415156 6012
rect 415212 6010 415236 6012
rect 415292 6010 415316 6012
rect 415372 6010 415386 6012
rect 415066 5958 415076 6010
rect 415132 5958 415142 6010
rect 414822 5956 414836 5958
rect 414892 5956 414916 5958
rect 414972 5956 414996 5958
rect 415052 5956 415076 5958
rect 415132 5956 415156 5958
rect 415212 5956 415236 5958
rect 415292 5956 415316 5958
rect 415372 5956 415386 5958
rect 414822 5936 415386 5956
rect 413928 5704 413980 5710
rect 413928 5646 413980 5652
rect 416688 5704 416740 5710
rect 416688 5646 416740 5652
rect 416504 5636 416556 5642
rect 416504 5578 416556 5584
rect 414664 5568 414716 5574
rect 414664 5510 414716 5516
rect 414480 4140 414532 4146
rect 414480 4082 414532 4088
rect 413744 3052 413796 3058
rect 413744 2994 413796 3000
rect 414492 480 414520 4082
rect 414676 2854 414704 5510
rect 414822 4924 415386 4944
rect 414822 4922 414836 4924
rect 414892 4922 414916 4924
rect 414972 4922 414996 4924
rect 415052 4922 415076 4924
rect 415132 4922 415156 4924
rect 415212 4922 415236 4924
rect 415292 4922 415316 4924
rect 415372 4922 415386 4924
rect 415066 4870 415076 4922
rect 415132 4870 415142 4922
rect 414822 4868 414836 4870
rect 414892 4868 414916 4870
rect 414972 4868 414996 4870
rect 415052 4868 415076 4870
rect 415132 4868 415156 4870
rect 415212 4868 415236 4870
rect 415292 4868 415316 4870
rect 415372 4868 415386 4870
rect 414822 4848 415386 4868
rect 414822 3836 415386 3856
rect 414822 3834 414836 3836
rect 414892 3834 414916 3836
rect 414972 3834 414996 3836
rect 415052 3834 415076 3836
rect 415132 3834 415156 3836
rect 415212 3834 415236 3836
rect 415292 3834 415316 3836
rect 415372 3834 415386 3836
rect 415066 3782 415076 3834
rect 415132 3782 415142 3834
rect 414822 3780 414836 3782
rect 414892 3780 414916 3782
rect 414972 3780 414996 3782
rect 415052 3780 415076 3782
rect 415132 3780 415156 3782
rect 415212 3780 415236 3782
rect 415292 3780 415316 3782
rect 415372 3780 415386 3782
rect 414822 3760 415386 3780
rect 416516 3602 416544 5578
rect 416504 3596 416556 3602
rect 416504 3538 416556 3544
rect 415676 3528 415728 3534
rect 415676 3470 415728 3476
rect 414664 2848 414716 2854
rect 414664 2790 414716 2796
rect 414822 2748 415386 2768
rect 414822 2746 414836 2748
rect 414892 2746 414916 2748
rect 414972 2746 414996 2748
rect 415052 2746 415076 2748
rect 415132 2746 415156 2748
rect 415212 2746 415236 2748
rect 415292 2746 415316 2748
rect 415372 2746 415386 2748
rect 415066 2694 415076 2746
rect 415132 2694 415142 2746
rect 414822 2692 414836 2694
rect 414892 2692 414916 2694
rect 414972 2692 414996 2694
rect 415052 2692 415076 2694
rect 415132 2692 415156 2694
rect 415212 2692 415236 2694
rect 415292 2692 415316 2694
rect 415372 2692 415386 2694
rect 414822 2672 415386 2692
rect 415688 480 415716 3470
rect 416700 3398 416728 5646
rect 416976 3466 417004 6190
rect 417344 5574 417372 8092
rect 418160 6384 418212 6390
rect 418160 6326 418212 6332
rect 417332 5568 417384 5574
rect 417332 5510 417384 5516
rect 418172 4078 418200 6326
rect 418540 6322 418568 8092
rect 418528 6316 418580 6322
rect 418528 6258 418580 6264
rect 419644 6118 419672 8092
rect 419632 6112 419684 6118
rect 419632 6054 419684 6060
rect 420840 5846 420868 8092
rect 420920 6316 420972 6322
rect 420920 6258 420972 6264
rect 420828 5840 420880 5846
rect 420828 5782 420880 5788
rect 419816 5568 419868 5574
rect 419816 5510 419868 5516
rect 418160 4072 418212 4078
rect 418160 4014 418212 4020
rect 419828 3534 419856 5510
rect 420932 3738 420960 6258
rect 421944 5914 421972 8092
rect 421932 5908 421984 5914
rect 421932 5850 421984 5856
rect 423140 5642 423168 8092
rect 423588 6112 423640 6118
rect 423588 6054 423640 6060
rect 423312 5840 423364 5846
rect 423312 5782 423364 5788
rect 423128 5636 423180 5642
rect 423128 5578 423180 5584
rect 420920 3732 420972 3738
rect 420920 3674 420972 3680
rect 420368 3596 420420 3602
rect 420368 3538 420420 3544
rect 419816 3528 419868 3534
rect 419816 3470 419868 3476
rect 416872 3460 416924 3466
rect 416872 3402 416924 3408
rect 416964 3460 417016 3466
rect 416964 3402 417016 3408
rect 416688 3392 416740 3398
rect 416688 3334 416740 3340
rect 416884 480 416912 3402
rect 417976 3052 418028 3058
rect 417976 2994 418028 3000
rect 417988 480 418016 2994
rect 419172 2848 419224 2854
rect 419172 2790 419224 2796
rect 419184 480 419212 2790
rect 420380 480 420408 3538
rect 422760 3460 422812 3466
rect 422760 3402 422812 3408
rect 421564 3392 421616 3398
rect 421564 3334 421616 3340
rect 421576 480 421604 3334
rect 422772 480 422800 3402
rect 423324 2922 423352 5782
rect 423600 3194 423628 6054
rect 424244 5574 424272 8092
rect 424508 5908 424560 5914
rect 424508 5850 424560 5856
rect 424232 5568 424284 5574
rect 424232 5510 424284 5516
rect 423956 4072 424008 4078
rect 423956 4014 424008 4020
rect 423588 3188 423640 3194
rect 423588 3130 423640 3136
rect 423312 2916 423364 2922
rect 423312 2858 423364 2864
rect 423968 480 423996 4014
rect 424520 2990 424548 5850
rect 425348 5846 425376 8092
rect 425336 5840 425388 5846
rect 425336 5782 425388 5788
rect 426256 5636 426308 5642
rect 426256 5578 426308 5584
rect 426268 3534 426296 5578
rect 426544 5574 426572 8092
rect 427648 6254 427676 8092
rect 427636 6248 427688 6254
rect 427636 6190 427688 6196
rect 427820 5840 427872 5846
rect 427820 5782 427872 5788
rect 426440 5568 426492 5574
rect 426440 5510 426492 5516
rect 426532 5568 426584 5574
rect 426532 5510 426584 5516
rect 426348 3732 426400 3738
rect 426348 3674 426400 3680
rect 425152 3528 425204 3534
rect 425152 3470 425204 3476
rect 426256 3528 426308 3534
rect 426256 3470 426308 3476
rect 424508 2984 424560 2990
rect 424508 2926 424560 2932
rect 425164 480 425192 3470
rect 426360 480 426388 3674
rect 426452 3126 426480 5510
rect 427832 3466 427860 5782
rect 428844 5710 428872 8092
rect 429844 6248 429896 6254
rect 429844 6190 429896 6196
rect 428832 5704 428884 5710
rect 428832 5646 428884 5652
rect 429200 5568 429252 5574
rect 429200 5510 429252 5516
rect 429212 4078 429240 5510
rect 429200 4072 429252 4078
rect 429200 4014 429252 4020
rect 429856 3670 429884 6190
rect 429948 5574 429976 8092
rect 431144 5914 431172 8092
rect 431132 5908 431184 5914
rect 431132 5850 431184 5856
rect 430580 5704 430632 5710
rect 430580 5646 430632 5652
rect 429936 5568 429988 5574
rect 429936 5510 429988 5516
rect 429844 3664 429896 3670
rect 429844 3606 429896 3612
rect 430592 3602 430620 5646
rect 432248 5642 432276 8092
rect 433444 6254 433472 8092
rect 433432 6248 433484 6254
rect 433432 6190 433484 6196
rect 434548 6186 434576 8092
rect 434536 6180 434588 6186
rect 434536 6122 434588 6128
rect 434168 5908 434220 5914
rect 434168 5850 434220 5856
rect 432236 5636 432288 5642
rect 432236 5578 432288 5584
rect 432696 5568 432748 5574
rect 432696 5510 432748 5516
rect 430580 3596 430632 3602
rect 430580 3538 430632 3544
rect 431132 3528 431184 3534
rect 431132 3470 431184 3476
rect 427820 3460 427872 3466
rect 427820 3402 427872 3408
rect 427544 3188 427596 3194
rect 427544 3130 427596 3136
rect 426440 3120 426492 3126
rect 426440 3062 426492 3068
rect 427556 480 427584 3130
rect 429936 2984 429988 2990
rect 429936 2926 429988 2932
rect 428740 2916 428792 2922
rect 428740 2858 428792 2864
rect 428752 480 428780 2858
rect 429948 480 429976 2926
rect 431144 480 431172 3470
rect 432328 3120 432380 3126
rect 432328 3062 432380 3068
rect 432340 480 432368 3062
rect 432708 2922 432736 5510
rect 432822 5468 433386 5488
rect 432822 5466 432836 5468
rect 432892 5466 432916 5468
rect 432972 5466 432996 5468
rect 433052 5466 433076 5468
rect 433132 5466 433156 5468
rect 433212 5466 433236 5468
rect 433292 5466 433316 5468
rect 433372 5466 433386 5468
rect 433066 5414 433076 5466
rect 433132 5414 433142 5466
rect 432822 5412 432836 5414
rect 432892 5412 432916 5414
rect 432972 5412 432996 5414
rect 433052 5412 433076 5414
rect 433132 5412 433156 5414
rect 433212 5412 433236 5414
rect 433292 5412 433316 5414
rect 433372 5412 433386 5414
rect 432822 5392 433386 5412
rect 432822 4380 433386 4400
rect 432822 4378 432836 4380
rect 432892 4378 432916 4380
rect 432972 4378 432996 4380
rect 433052 4378 433076 4380
rect 433132 4378 433156 4380
rect 433212 4378 433236 4380
rect 433292 4378 433316 4380
rect 433372 4378 433386 4380
rect 433066 4326 433076 4378
rect 433132 4326 433142 4378
rect 432822 4324 432836 4326
rect 432892 4324 432916 4326
rect 432972 4324 432996 4326
rect 433052 4324 433076 4326
rect 433132 4324 433156 4326
rect 433212 4324 433236 4326
rect 433292 4324 433316 4326
rect 433372 4324 433386 4326
rect 432822 4304 433386 4324
rect 433524 3460 433576 3466
rect 433524 3402 433576 3408
rect 432822 3292 433386 3312
rect 432822 3290 432836 3292
rect 432892 3290 432916 3292
rect 432972 3290 432996 3292
rect 433052 3290 433076 3292
rect 433132 3290 433156 3292
rect 433212 3290 433236 3292
rect 433292 3290 433316 3292
rect 433372 3290 433386 3292
rect 433066 3238 433076 3290
rect 433132 3238 433142 3290
rect 432822 3236 432836 3238
rect 432892 3236 432916 3238
rect 432972 3236 432996 3238
rect 433052 3236 433076 3238
rect 433132 3236 433156 3238
rect 433212 3236 433236 3238
rect 433292 3236 433316 3238
rect 433372 3236 433386 3238
rect 432822 3216 433386 3236
rect 432696 2916 432748 2922
rect 432696 2858 432748 2864
rect 432822 2204 433386 2224
rect 432822 2202 432836 2204
rect 432892 2202 432916 2204
rect 432972 2202 432996 2204
rect 433052 2202 433076 2204
rect 433132 2202 433156 2204
rect 433212 2202 433236 2204
rect 433292 2202 433316 2204
rect 433372 2202 433386 2204
rect 433066 2150 433076 2202
rect 433132 2150 433142 2202
rect 432822 2148 432836 2150
rect 432892 2148 432916 2150
rect 432972 2148 432996 2150
rect 433052 2148 433076 2150
rect 433132 2148 433156 2150
rect 433212 2148 433236 2150
rect 433292 2148 433316 2150
rect 433372 2148 433386 2150
rect 432822 2128 433386 2148
rect 433536 480 433564 3402
rect 434180 3058 434208 5850
rect 435652 5574 435680 8092
rect 436100 6248 436152 6254
rect 436100 6190 436152 6196
rect 436008 5636 436060 5642
rect 436008 5578 436060 5584
rect 435640 5568 435692 5574
rect 435640 5510 435692 5516
rect 434628 4072 434680 4078
rect 434628 4014 434680 4020
rect 434168 3052 434220 3058
rect 434168 2994 434220 3000
rect 434640 480 434668 4014
rect 435824 3664 435876 3670
rect 435824 3606 435876 3612
rect 435836 480 435864 3606
rect 436020 3534 436048 5578
rect 436008 3528 436060 3534
rect 436008 3470 436060 3476
rect 436112 3398 436140 6190
rect 436848 6118 436876 8092
rect 437952 6254 437980 8092
rect 437940 6248 437992 6254
rect 437940 6190 437992 6196
rect 436836 6112 436888 6118
rect 436836 6054 436888 6060
rect 439148 5574 439176 8092
rect 439228 6112 439280 6118
rect 439228 6054 439280 6060
rect 438584 5568 438636 5574
rect 438584 5510 438636 5516
rect 439136 5568 439188 5574
rect 439136 5510 439188 5516
rect 438596 4078 438624 5510
rect 438584 4072 438636 4078
rect 438584 4014 438636 4020
rect 437020 3596 437072 3602
rect 437020 3538 437072 3544
rect 436100 3392 436152 3398
rect 436100 3334 436152 3340
rect 437032 480 437060 3538
rect 439240 3466 439268 6054
rect 440252 5914 440280 8092
rect 440332 6248 440384 6254
rect 440332 6190 440384 6196
rect 440240 5908 440292 5914
rect 440240 5850 440292 5856
rect 440344 3670 440372 6190
rect 441448 5846 441476 8092
rect 442552 6390 442580 8092
rect 442540 6384 442592 6390
rect 442540 6326 442592 6332
rect 443000 6180 443052 6186
rect 443000 6122 443052 6128
rect 441436 5840 441488 5846
rect 441436 5782 441488 5788
rect 442080 5568 442132 5574
rect 442080 5510 442132 5516
rect 442092 3942 442120 5510
rect 442080 3936 442132 3942
rect 442080 3878 442132 3884
rect 440332 3664 440384 3670
rect 440332 3606 440384 3612
rect 440608 3528 440660 3534
rect 440608 3470 440660 3476
rect 439228 3460 439280 3466
rect 439228 3402 439280 3408
rect 439412 3052 439464 3058
rect 439412 2994 439464 3000
rect 438216 2916 438268 2922
rect 438216 2858 438268 2864
rect 438228 480 438256 2858
rect 439424 480 439452 2994
rect 440620 480 440648 3470
rect 441804 3392 441856 3398
rect 441804 3334 441856 3340
rect 441816 480 441844 3334
rect 443012 480 443040 6122
rect 443748 5846 443776 8092
rect 443828 5908 443880 5914
rect 443828 5850 443880 5856
rect 443460 5840 443512 5846
rect 443460 5782 443512 5788
rect 443736 5840 443788 5846
rect 443736 5782 443788 5788
rect 443472 2922 443500 5782
rect 443840 2990 443868 5850
rect 444852 5710 444880 8092
rect 445484 6384 445536 6390
rect 445484 6326 445536 6332
rect 444840 5704 444892 5710
rect 444840 5646 444892 5652
rect 444196 4072 444248 4078
rect 444196 4014 444248 4020
rect 443828 2984 443880 2990
rect 443828 2926 443880 2932
rect 443460 2916 443512 2922
rect 443460 2858 443512 2864
rect 444208 480 444236 4014
rect 445496 3466 445524 6326
rect 445956 5846 445984 8092
rect 447152 6118 447180 8092
rect 448256 6254 448284 8092
rect 449452 6390 449480 8092
rect 450556 6798 450584 8092
rect 450544 6792 450596 6798
rect 450544 6734 450596 6740
rect 449440 6384 449492 6390
rect 449440 6326 449492 6332
rect 448244 6248 448296 6254
rect 448244 6190 448296 6196
rect 447140 6112 447192 6118
rect 447140 6054 447192 6060
rect 449900 6112 449952 6118
rect 449900 6054 449952 6060
rect 445852 5840 445904 5846
rect 445852 5782 445904 5788
rect 445944 5840 445996 5846
rect 445944 5782 445996 5788
rect 448612 5840 448664 5846
rect 448612 5782 448664 5788
rect 445392 3460 445444 3466
rect 445392 3402 445444 3408
rect 445484 3460 445536 3466
rect 445484 3402 445536 3408
rect 445404 480 445432 3402
rect 445864 3194 445892 5782
rect 448060 5704 448112 5710
rect 448060 5646 448112 5652
rect 448072 4146 448100 5646
rect 448060 4140 448112 4146
rect 448060 4082 448112 4088
rect 448624 3942 448652 5782
rect 447784 3936 447836 3942
rect 447784 3878 447836 3884
rect 448612 3936 448664 3942
rect 448612 3878 448664 3884
rect 446588 3664 446640 3670
rect 446588 3606 446640 3612
rect 445852 3188 445904 3194
rect 445852 3130 445904 3136
rect 446600 480 446628 3606
rect 447796 480 447824 3878
rect 449912 3738 449940 6054
rect 450822 6012 451386 6032
rect 450822 6010 450836 6012
rect 450892 6010 450916 6012
rect 450972 6010 450996 6012
rect 451052 6010 451076 6012
rect 451132 6010 451156 6012
rect 451212 6010 451236 6012
rect 451292 6010 451316 6012
rect 451372 6010 451386 6012
rect 451066 5958 451076 6010
rect 451132 5958 451142 6010
rect 450822 5956 450836 5958
rect 450892 5956 450916 5958
rect 450972 5956 450996 5958
rect 451052 5956 451076 5958
rect 451132 5956 451156 5958
rect 451212 5956 451236 5958
rect 451292 5956 451316 5958
rect 451372 5956 451386 5958
rect 450822 5936 451386 5956
rect 451752 5642 451780 8092
rect 451740 5636 451792 5642
rect 451740 5578 451792 5584
rect 452856 5574 452884 8092
rect 454052 6118 454080 8092
rect 455156 6186 455184 8092
rect 455144 6180 455196 6186
rect 455144 6122 455196 6128
rect 454040 6112 454092 6118
rect 454040 6054 454092 6060
rect 456352 5846 456380 8092
rect 457260 6248 457312 6254
rect 457260 6190 457312 6196
rect 456340 5840 456392 5846
rect 456340 5782 456392 5788
rect 455328 5636 455380 5642
rect 455328 5578 455380 5584
rect 452844 5568 452896 5574
rect 452844 5510 452896 5516
rect 450822 4924 451386 4944
rect 450822 4922 450836 4924
rect 450892 4922 450916 4924
rect 450972 4922 450996 4924
rect 451052 4922 451076 4924
rect 451132 4922 451156 4924
rect 451212 4922 451236 4924
rect 451292 4922 451316 4924
rect 451372 4922 451386 4924
rect 451066 4870 451076 4922
rect 451132 4870 451142 4922
rect 450822 4868 450836 4870
rect 450892 4868 450916 4870
rect 450972 4868 450996 4870
rect 451052 4868 451076 4870
rect 451132 4868 451156 4870
rect 451212 4868 451236 4870
rect 451292 4868 451316 4870
rect 451372 4868 451386 4870
rect 450822 4848 451386 4868
rect 453672 4140 453724 4146
rect 453672 4082 453724 4088
rect 450822 3836 451386 3856
rect 450822 3834 450836 3836
rect 450892 3834 450916 3836
rect 450972 3834 450996 3836
rect 451052 3834 451076 3836
rect 451132 3834 451156 3836
rect 451212 3834 451236 3836
rect 451292 3834 451316 3836
rect 451372 3834 451386 3836
rect 451066 3782 451076 3834
rect 451132 3782 451142 3834
rect 450822 3780 450836 3782
rect 450892 3780 450916 3782
rect 450972 3780 450996 3782
rect 451052 3780 451076 3782
rect 451132 3780 451156 3782
rect 451212 3780 451236 3782
rect 451292 3780 451316 3782
rect 451372 3780 451386 3782
rect 450822 3760 451386 3780
rect 449900 3732 449952 3738
rect 449900 3674 449952 3680
rect 451464 3460 451516 3466
rect 451464 3402 451516 3408
rect 448980 2984 449032 2990
rect 448980 2926 449032 2932
rect 448992 480 449020 2926
rect 450176 2916 450228 2922
rect 450176 2858 450228 2864
rect 450188 480 450216 2858
rect 450822 2748 451386 2768
rect 450822 2746 450836 2748
rect 450892 2746 450916 2748
rect 450972 2746 450996 2748
rect 451052 2746 451076 2748
rect 451132 2746 451156 2748
rect 451212 2746 451236 2748
rect 451292 2746 451316 2748
rect 451372 2746 451386 2748
rect 451066 2694 451076 2746
rect 451132 2694 451142 2746
rect 450822 2692 450836 2694
rect 450892 2692 450916 2694
rect 450972 2692 450996 2694
rect 451052 2692 451076 2694
rect 451132 2692 451156 2694
rect 451212 2692 451236 2694
rect 451292 2692 451316 2694
rect 451372 2692 451386 2694
rect 450822 2672 451386 2692
rect 451476 2530 451504 3402
rect 452476 3188 452528 3194
rect 452476 3130 452528 3136
rect 451292 2502 451504 2530
rect 451292 480 451320 2502
rect 452488 480 452516 3130
rect 453684 480 453712 4082
rect 454868 3936 454920 3942
rect 454868 3878 454920 3884
rect 454880 480 454908 3878
rect 455340 3058 455368 5578
rect 455420 5568 455472 5574
rect 455420 5510 455472 5516
rect 455432 3126 455460 5510
rect 456064 3732 456116 3738
rect 456064 3674 456116 3680
rect 455420 3120 455472 3126
rect 455420 3062 455472 3068
rect 455328 3052 455380 3058
rect 455328 2994 455380 3000
rect 456076 480 456104 3674
rect 457272 480 457300 6190
rect 457456 5710 457484 8092
rect 458560 6730 458588 8092
rect 459652 6792 459704 6798
rect 459652 6734 459704 6740
rect 458548 6724 458600 6730
rect 458548 6666 458600 6672
rect 458456 6384 458508 6390
rect 458456 6326 458508 6332
rect 457536 6112 457588 6118
rect 457536 6054 457588 6060
rect 457444 5704 457496 5710
rect 457444 5646 457496 5652
rect 457548 4078 457576 6054
rect 457536 4072 457588 4078
rect 457536 4014 457588 4020
rect 458468 480 458496 6326
rect 458640 5840 458692 5846
rect 458640 5782 458692 5788
rect 458652 3466 458680 5782
rect 459560 5704 459612 5710
rect 459560 5646 459612 5652
rect 459572 3534 459600 5646
rect 459560 3528 459612 3534
rect 459560 3470 459612 3476
rect 458640 3460 458692 3466
rect 458640 3402 458692 3408
rect 459664 480 459692 6734
rect 459756 5574 459784 8092
rect 460860 6118 460888 8092
rect 462056 6254 462084 8092
rect 463160 6390 463188 8092
rect 464356 6458 464384 8092
rect 464344 6452 464396 6458
rect 464344 6394 464396 6400
rect 463148 6384 463200 6390
rect 463148 6326 463200 6332
rect 465460 6322 465488 8092
rect 466656 6526 466684 8092
rect 466644 6520 466696 6526
rect 466644 6462 466696 6468
rect 465448 6316 465500 6322
rect 465448 6258 465500 6264
rect 462044 6248 462096 6254
rect 462044 6190 462096 6196
rect 467760 6186 467788 8092
rect 467932 6724 467984 6730
rect 467932 6666 467984 6672
rect 464436 6180 464488 6186
rect 464436 6122 464488 6128
rect 467748 6180 467800 6186
rect 467748 6122 467800 6128
rect 460848 6112 460900 6118
rect 460848 6054 460900 6060
rect 459744 5568 459796 5574
rect 459744 5510 459796 5516
rect 463608 5568 463660 5574
rect 463608 5510 463660 5516
rect 463240 4072 463292 4078
rect 463240 4014 463292 4020
rect 462044 3120 462096 3126
rect 462044 3062 462096 3068
rect 460848 3052 460900 3058
rect 460848 2994 460900 3000
rect 460860 480 460888 2994
rect 462056 480 462084 3062
rect 463252 480 463280 4014
rect 463620 3194 463648 5510
rect 463608 3188 463660 3194
rect 463608 3130 463660 3136
rect 464448 480 464476 6122
rect 466828 3528 466880 3534
rect 466828 3470 466880 3476
rect 465632 3460 465684 3466
rect 465632 3402 465684 3408
rect 465644 480 465672 3402
rect 466840 480 466868 3470
rect 467944 480 467972 6666
rect 468864 6594 468892 8092
rect 470060 6662 470088 8092
rect 470048 6656 470100 6662
rect 470048 6598 470100 6604
rect 468852 6588 468904 6594
rect 468852 6530 468904 6536
rect 470324 6112 470376 6118
rect 470324 6054 470376 6060
rect 468822 5468 469386 5488
rect 468822 5466 468836 5468
rect 468892 5466 468916 5468
rect 468972 5466 468996 5468
rect 469052 5466 469076 5468
rect 469132 5466 469156 5468
rect 469212 5466 469236 5468
rect 469292 5466 469316 5468
rect 469372 5466 469386 5468
rect 469066 5414 469076 5466
rect 469132 5414 469142 5466
rect 468822 5412 468836 5414
rect 468892 5412 468916 5414
rect 468972 5412 468996 5414
rect 469052 5412 469076 5414
rect 469132 5412 469156 5414
rect 469212 5412 469236 5414
rect 469292 5412 469316 5414
rect 469372 5412 469386 5414
rect 468822 5392 469386 5412
rect 468822 4380 469386 4400
rect 468822 4378 468836 4380
rect 468892 4378 468916 4380
rect 468972 4378 468996 4380
rect 469052 4378 469076 4380
rect 469132 4378 469156 4380
rect 469212 4378 469236 4380
rect 469292 4378 469316 4380
rect 469372 4378 469386 4380
rect 469066 4326 469076 4378
rect 469132 4326 469142 4378
rect 468822 4324 468836 4326
rect 468892 4324 468916 4326
rect 468972 4324 468996 4326
rect 469052 4324 469076 4326
rect 469132 4324 469156 4326
rect 469212 4324 469236 4326
rect 469292 4324 469316 4326
rect 469372 4324 469386 4326
rect 468822 4304 469386 4324
rect 468822 3292 469386 3312
rect 468822 3290 468836 3292
rect 468892 3290 468916 3292
rect 468972 3290 468996 3292
rect 469052 3290 469076 3292
rect 469132 3290 469156 3292
rect 469212 3290 469236 3292
rect 469292 3290 469316 3292
rect 469372 3290 469386 3292
rect 469066 3238 469076 3290
rect 469132 3238 469142 3290
rect 468822 3236 468836 3238
rect 468892 3236 468916 3238
rect 468972 3236 468996 3238
rect 469052 3236 469076 3238
rect 469132 3236 469156 3238
rect 469212 3236 469236 3238
rect 469292 3236 469316 3238
rect 469372 3236 469386 3238
rect 468822 3216 469386 3236
rect 468668 3188 468720 3194
rect 468668 3130 468720 3136
rect 468680 1986 468708 3130
rect 468822 2204 469386 2224
rect 468822 2202 468836 2204
rect 468892 2202 468916 2204
rect 468972 2202 468996 2204
rect 469052 2202 469076 2204
rect 469132 2202 469156 2204
rect 469212 2202 469236 2204
rect 469292 2202 469316 2204
rect 469372 2202 469386 2204
rect 469066 2150 469076 2202
rect 469132 2150 469142 2202
rect 468822 2148 468836 2150
rect 468892 2148 468916 2150
rect 468972 2148 468996 2150
rect 469052 2148 469076 2150
rect 469132 2148 469156 2150
rect 469212 2148 469236 2150
rect 469292 2148 469316 2150
rect 469372 2148 469386 2150
rect 468822 2128 469386 2148
rect 468680 1958 469168 1986
rect 469140 480 469168 1958
rect 470336 480 470364 6054
rect 471164 5710 471192 8092
rect 471520 6248 471572 6254
rect 471520 6190 471572 6196
rect 471152 5704 471204 5710
rect 471152 5646 471204 5652
rect 471532 480 471560 6190
rect 472360 5574 472388 8092
rect 472716 6384 472768 6390
rect 472716 6326 472768 6332
rect 472348 5568 472400 5574
rect 472348 5510 472400 5516
rect 472728 480 472756 6326
rect 473464 6254 473492 8092
rect 473912 6452 473964 6458
rect 473912 6394 473964 6400
rect 473452 6248 473504 6254
rect 473452 6190 473504 6196
rect 473360 5704 473412 5710
rect 473360 5646 473412 5652
rect 473372 3466 473400 5646
rect 473360 3460 473412 3466
rect 473360 3402 473412 3408
rect 473924 480 473952 6394
rect 474660 6390 474688 8092
rect 475764 6458 475792 8092
rect 476960 6730 476988 8092
rect 476948 6724 477000 6730
rect 476948 6666 477000 6672
rect 476304 6520 476356 6526
rect 476304 6462 476356 6468
rect 475752 6452 475804 6458
rect 475752 6394 475804 6400
rect 474648 6384 474700 6390
rect 474648 6326 474700 6332
rect 475108 6316 475160 6322
rect 475108 6258 475160 6264
rect 474740 5568 474792 5574
rect 474740 5510 474792 5516
rect 474752 3398 474780 5510
rect 474740 3392 474792 3398
rect 474740 3334 474792 3340
rect 475120 480 475148 6258
rect 476316 480 476344 6462
rect 477500 6180 477552 6186
rect 477500 6122 477552 6128
rect 477512 480 477540 6122
rect 478064 6118 478092 8092
rect 479168 6594 479196 8092
rect 479892 6656 479944 6662
rect 479892 6598 479944 6604
rect 478696 6588 478748 6594
rect 478696 6530 478748 6536
rect 479156 6588 479208 6594
rect 479156 6530 479208 6536
rect 478052 6112 478104 6118
rect 478052 6054 478104 6060
rect 478708 480 478736 6530
rect 479904 480 479932 6598
rect 480364 5914 480392 8092
rect 481468 6322 481496 8092
rect 481456 6316 481508 6322
rect 481456 6258 481508 6264
rect 482664 6186 482692 8092
rect 483768 6526 483796 8092
rect 484964 6866 484992 8092
rect 484952 6860 485004 6866
rect 484952 6802 485004 6808
rect 486068 6662 486096 8092
rect 486700 6724 486752 6730
rect 486700 6666 486752 6672
rect 486056 6656 486108 6662
rect 486056 6598 486108 6604
rect 483756 6520 483808 6526
rect 483756 6462 483808 6468
rect 485688 6452 485740 6458
rect 485688 6394 485740 6400
rect 484584 6384 484636 6390
rect 484584 6326 484636 6332
rect 483480 6248 483532 6254
rect 483480 6190 483532 6196
rect 482652 6180 482704 6186
rect 482652 6122 482704 6128
rect 480352 5908 480404 5914
rect 480352 5850 480404 5856
rect 481088 3460 481140 3466
rect 481088 3402 481140 3408
rect 481100 480 481128 3402
rect 482284 3392 482336 3398
rect 482284 3334 482336 3340
rect 482296 480 482324 3334
rect 483492 480 483520 6190
rect 484596 480 484624 6326
rect 485700 4026 485728 6394
rect 485700 3998 485820 4026
rect 485792 480 485820 3998
rect 486712 2530 486740 6666
rect 487264 6254 487292 8092
rect 487252 6248 487304 6254
rect 487252 6190 487304 6196
rect 488172 6112 488224 6118
rect 488172 6054 488224 6060
rect 486822 6012 487386 6032
rect 486822 6010 486836 6012
rect 486892 6010 486916 6012
rect 486972 6010 486996 6012
rect 487052 6010 487076 6012
rect 487132 6010 487156 6012
rect 487212 6010 487236 6012
rect 487292 6010 487316 6012
rect 487372 6010 487386 6012
rect 487066 5958 487076 6010
rect 487132 5958 487142 6010
rect 486822 5956 486836 5958
rect 486892 5956 486916 5958
rect 486972 5956 486996 5958
rect 487052 5956 487076 5958
rect 487132 5956 487156 5958
rect 487212 5956 487236 5958
rect 487292 5956 487316 5958
rect 487372 5956 487386 5958
rect 486822 5936 487386 5956
rect 486822 4924 487386 4944
rect 486822 4922 486836 4924
rect 486892 4922 486916 4924
rect 486972 4922 486996 4924
rect 487052 4922 487076 4924
rect 487132 4922 487156 4924
rect 487212 4922 487236 4924
rect 487292 4922 487316 4924
rect 487372 4922 487386 4924
rect 487066 4870 487076 4922
rect 487132 4870 487142 4922
rect 486822 4868 486836 4870
rect 486892 4868 486916 4870
rect 486972 4868 486996 4870
rect 487052 4868 487076 4870
rect 487132 4868 487156 4870
rect 487212 4868 487236 4870
rect 487292 4868 487316 4870
rect 487372 4868 487386 4870
rect 486822 4848 487386 4868
rect 486822 3836 487386 3856
rect 486822 3834 486836 3836
rect 486892 3834 486916 3836
rect 486972 3834 486996 3836
rect 487052 3834 487076 3836
rect 487132 3834 487156 3836
rect 487212 3834 487236 3836
rect 487292 3834 487316 3836
rect 487372 3834 487386 3836
rect 487066 3782 487076 3834
rect 487132 3782 487142 3834
rect 486822 3780 486836 3782
rect 486892 3780 486916 3782
rect 486972 3780 486996 3782
rect 487052 3780 487076 3782
rect 487132 3780 487156 3782
rect 487212 3780 487236 3782
rect 487292 3780 487316 3782
rect 487372 3780 487386 3782
rect 486822 3760 487386 3780
rect 486822 2748 487386 2768
rect 486822 2746 486836 2748
rect 486892 2746 486916 2748
rect 486972 2746 486996 2748
rect 487052 2746 487076 2748
rect 487132 2746 487156 2748
rect 487212 2746 487236 2748
rect 487292 2746 487316 2748
rect 487372 2746 487386 2748
rect 487066 2694 487076 2746
rect 487132 2694 487142 2746
rect 486822 2692 486836 2694
rect 486892 2692 486916 2694
rect 486972 2692 486996 2694
rect 487052 2692 487076 2694
rect 487132 2692 487156 2694
rect 487212 2692 487236 2694
rect 487292 2692 487316 2694
rect 487372 2692 487386 2694
rect 486822 2672 487386 2692
rect 486712 2502 487016 2530
rect 486988 480 487016 2502
rect 488184 480 488212 6054
rect 488368 5710 488396 8092
rect 489368 6588 489420 6594
rect 489368 6530 489420 6536
rect 488356 5704 488408 5710
rect 488356 5646 488408 5652
rect 489380 480 489408 6530
rect 489472 6390 489500 8092
rect 490668 6594 490696 8092
rect 491772 6882 491800 8092
rect 491680 6854 491800 6882
rect 490656 6588 490708 6594
rect 490656 6530 490708 6536
rect 489460 6384 489512 6390
rect 489460 6326 489512 6332
rect 490748 6248 490800 6254
rect 490748 6190 490800 6196
rect 490564 5908 490616 5914
rect 490564 5850 490616 5856
rect 490380 5704 490432 5710
rect 490380 5646 490432 5652
rect 490392 3942 490420 5646
rect 490380 3936 490432 3942
rect 490380 3878 490432 3884
rect 490576 480 490604 5850
rect 490760 3126 490788 6190
rect 491680 5914 491708 6854
rect 492968 6730 492996 8092
rect 494072 6798 494100 8092
rect 494060 6792 494112 6798
rect 494060 6734 494112 6740
rect 492956 6724 493008 6730
rect 492956 6666 493008 6672
rect 495268 6526 495296 8092
rect 495348 6860 495400 6866
rect 495348 6802 495400 6808
rect 494152 6520 494204 6526
rect 494152 6462 494204 6468
rect 495256 6520 495308 6526
rect 495256 6462 495308 6468
rect 491760 6316 491812 6322
rect 491760 6258 491812 6264
rect 491668 5908 491720 5914
rect 491668 5850 491720 5856
rect 490748 3120 490800 3126
rect 490748 3062 490800 3068
rect 491772 480 491800 6258
rect 492956 6180 493008 6186
rect 492956 6122 493008 6128
rect 492968 480 492996 6122
rect 494164 480 494192 6462
rect 495360 480 495388 6802
rect 496372 6322 496400 8092
rect 496544 6656 496596 6662
rect 496544 6598 496596 6604
rect 496360 6316 496412 6322
rect 496360 6258 496412 6264
rect 496556 480 496584 6598
rect 497568 6254 497596 8092
rect 497556 6248 497608 6254
rect 497556 6190 497608 6196
rect 498672 6186 498700 8092
rect 499882 8078 500264 8106
rect 500236 6390 500264 8078
rect 500132 6384 500184 6390
rect 500132 6326 500184 6332
rect 500224 6384 500276 6390
rect 500224 6326 500276 6332
rect 498660 6180 498712 6186
rect 498660 6122 498712 6128
rect 498936 3936 498988 3942
rect 498936 3878 498988 3884
rect 497740 3120 497792 3126
rect 497740 3062 497792 3068
rect 497752 480 497780 3062
rect 498948 480 498976 3878
rect 500144 480 500172 6326
rect 500972 6118 501000 8092
rect 501236 6588 501288 6594
rect 501236 6530 501288 6536
rect 500960 6112 501012 6118
rect 500960 6054 501012 6060
rect 501248 480 501276 6530
rect 502076 6458 502104 8092
rect 502064 6452 502116 6458
rect 502064 6394 502116 6400
rect 502248 5908 502300 5914
rect 502248 5850 502300 5856
rect 502260 4026 502288 5850
rect 503272 5574 503300 8092
rect 503628 6724 503680 6730
rect 503628 6666 503680 6672
rect 503260 5568 503312 5574
rect 503260 5510 503312 5516
rect 502260 3998 502472 4026
rect 502444 480 502472 3998
rect 503640 480 503668 6666
rect 504376 6594 504404 8092
rect 504732 6792 504784 6798
rect 504732 6734 504784 6740
rect 504364 6588 504416 6594
rect 504364 6530 504416 6536
rect 504744 1986 504772 6734
rect 505572 6662 505600 8092
rect 506676 6866 506704 8092
rect 506664 6860 506716 6866
rect 506664 6802 506716 6808
rect 507872 6798 507900 8092
rect 507860 6792 507912 6798
rect 507860 6734 507912 6740
rect 505560 6656 505612 6662
rect 505560 6598 505612 6604
rect 506020 6520 506072 6526
rect 506020 6462 506072 6468
rect 504822 5468 505386 5488
rect 504822 5466 504836 5468
rect 504892 5466 504916 5468
rect 504972 5466 504996 5468
rect 505052 5466 505076 5468
rect 505132 5466 505156 5468
rect 505212 5466 505236 5468
rect 505292 5466 505316 5468
rect 505372 5466 505386 5468
rect 505066 5414 505076 5466
rect 505132 5414 505142 5466
rect 504822 5412 504836 5414
rect 504892 5412 504916 5414
rect 504972 5412 504996 5414
rect 505052 5412 505076 5414
rect 505132 5412 505156 5414
rect 505212 5412 505236 5414
rect 505292 5412 505316 5414
rect 505372 5412 505386 5414
rect 504822 5392 505386 5412
rect 504822 4380 505386 4400
rect 504822 4378 504836 4380
rect 504892 4378 504916 4380
rect 504972 4378 504996 4380
rect 505052 4378 505076 4380
rect 505132 4378 505156 4380
rect 505212 4378 505236 4380
rect 505292 4378 505316 4380
rect 505372 4378 505386 4380
rect 505066 4326 505076 4378
rect 505132 4326 505142 4378
rect 504822 4324 504836 4326
rect 504892 4324 504916 4326
rect 504972 4324 504996 4326
rect 505052 4324 505076 4326
rect 505132 4324 505156 4326
rect 505212 4324 505236 4326
rect 505292 4324 505316 4326
rect 505372 4324 505386 4326
rect 504822 4304 505386 4324
rect 504822 3292 505386 3312
rect 504822 3290 504836 3292
rect 504892 3290 504916 3292
rect 504972 3290 504996 3292
rect 505052 3290 505076 3292
rect 505132 3290 505156 3292
rect 505212 3290 505236 3292
rect 505292 3290 505316 3292
rect 505372 3290 505386 3292
rect 505066 3238 505076 3290
rect 505132 3238 505142 3290
rect 504822 3236 504836 3238
rect 504892 3236 504916 3238
rect 504972 3236 504996 3238
rect 505052 3236 505076 3238
rect 505132 3236 505156 3238
rect 505212 3236 505236 3238
rect 505292 3236 505316 3238
rect 505372 3236 505386 3238
rect 504822 3216 505386 3236
rect 504822 2204 505386 2224
rect 504822 2202 504836 2204
rect 504892 2202 504916 2204
rect 504972 2202 504996 2204
rect 505052 2202 505076 2204
rect 505132 2202 505156 2204
rect 505212 2202 505236 2204
rect 505292 2202 505316 2204
rect 505372 2202 505386 2204
rect 505066 2150 505076 2202
rect 505132 2150 505142 2202
rect 504822 2148 504836 2150
rect 504892 2148 504916 2150
rect 504972 2148 504996 2150
rect 505052 2148 505076 2150
rect 505132 2148 505156 2150
rect 505212 2148 505236 2150
rect 505292 2148 505316 2150
rect 505372 2148 505386 2150
rect 504822 2128 505386 2148
rect 504744 1958 504864 1986
rect 504836 480 504864 1958
rect 506032 480 506060 6462
rect 507216 6316 507268 6322
rect 507216 6258 507268 6264
rect 506296 5568 506348 5574
rect 506296 5510 506348 5516
rect 506308 3466 506336 5510
rect 506296 3460 506348 3466
rect 506296 3402 506348 3408
rect 507228 480 507256 6258
rect 508976 6254 509004 8092
rect 510172 6526 510200 8092
rect 511276 6730 511304 8092
rect 511264 6724 511316 6730
rect 511264 6666 511316 6672
rect 510160 6520 510212 6526
rect 510160 6462 510212 6468
rect 512380 6458 512408 8092
rect 510988 6452 511040 6458
rect 510988 6394 511040 6400
rect 512368 6452 512420 6458
rect 512368 6394 512420 6400
rect 510804 6384 510856 6390
rect 510804 6326 510856 6332
rect 508412 6248 508464 6254
rect 508412 6190 508464 6196
rect 508964 6248 509016 6254
rect 508964 6190 509016 6196
rect 508424 480 508452 6190
rect 509608 6180 509660 6186
rect 509608 6122 509660 6128
rect 509620 480 509648 6122
rect 510816 480 510844 6326
rect 511000 3194 511028 6394
rect 513576 6390 513604 8092
rect 513564 6384 513616 6390
rect 513564 6326 513616 6332
rect 514680 6322 514708 8092
rect 515588 6588 515640 6594
rect 515588 6530 515640 6536
rect 514668 6316 514720 6322
rect 514668 6258 514720 6264
rect 511908 6112 511960 6118
rect 511908 6054 511960 6060
rect 511920 4026 511948 6054
rect 511920 3998 512040 4026
rect 510988 3188 511040 3194
rect 510988 3130 511040 3136
rect 512012 480 512040 3998
rect 514392 3460 514444 3466
rect 514392 3402 514444 3408
rect 513196 3188 513248 3194
rect 513196 3130 513248 3136
rect 513208 480 513236 3130
rect 514404 480 514432 3402
rect 515600 480 515628 6530
rect 515876 6186 515904 8092
rect 516140 6860 516192 6866
rect 516140 6802 516192 6808
rect 515864 6180 515916 6186
rect 515864 6122 515916 6128
rect 516152 3602 516180 6802
rect 516784 6656 516836 6662
rect 516784 6598 516836 6604
rect 516140 3596 516192 3602
rect 516140 3538 516192 3544
rect 516796 480 516824 6598
rect 516980 5914 517008 8092
rect 516968 5908 517020 5914
rect 516968 5850 517020 5856
rect 518176 5642 518204 8092
rect 519280 6866 519308 8092
rect 519268 6860 519320 6866
rect 519268 6802 519320 6808
rect 520476 6798 520504 8092
rect 519084 6792 519136 6798
rect 519084 6734 519136 6740
rect 520464 6792 520516 6798
rect 520464 6734 520516 6740
rect 518164 5636 518216 5642
rect 518164 5578 518216 5584
rect 517888 3596 517940 3602
rect 517888 3538 517940 3544
rect 517900 480 517928 3538
rect 519096 480 519124 6734
rect 521580 6594 521608 8092
rect 522592 8078 522698 8106
rect 523894 8078 524184 8106
rect 521568 6588 521620 6594
rect 521568 6530 521620 6536
rect 521476 6520 521528 6526
rect 521476 6462 521528 6468
rect 520188 6248 520240 6254
rect 520188 6190 520240 6196
rect 520200 4026 520228 6190
rect 520200 3998 520320 4026
rect 520292 480 520320 3998
rect 521488 480 521516 6462
rect 522592 6118 522620 8078
rect 522672 6724 522724 6730
rect 522672 6666 522724 6672
rect 522580 6112 522632 6118
rect 522580 6054 522632 6060
rect 521568 5636 521620 5642
rect 521568 5578 521620 5584
rect 521580 3466 521608 5578
rect 521568 3460 521620 3466
rect 521568 3402 521620 3408
rect 522684 480 522712 6666
rect 523868 6452 523920 6458
rect 523868 6394 523920 6400
rect 522822 6012 523386 6032
rect 522822 6010 522836 6012
rect 522892 6010 522916 6012
rect 522972 6010 522996 6012
rect 523052 6010 523076 6012
rect 523132 6010 523156 6012
rect 523212 6010 523236 6012
rect 523292 6010 523316 6012
rect 523372 6010 523386 6012
rect 523066 5958 523076 6010
rect 523132 5958 523142 6010
rect 522822 5956 522836 5958
rect 522892 5956 522916 5958
rect 522972 5956 522996 5958
rect 523052 5956 523076 5958
rect 523132 5956 523156 5958
rect 523212 5956 523236 5958
rect 523292 5956 523316 5958
rect 523372 5956 523386 5958
rect 522822 5936 523386 5956
rect 522822 4924 523386 4944
rect 522822 4922 522836 4924
rect 522892 4922 522916 4924
rect 522972 4922 522996 4924
rect 523052 4922 523076 4924
rect 523132 4922 523156 4924
rect 523212 4922 523236 4924
rect 523292 4922 523316 4924
rect 523372 4922 523386 4924
rect 523066 4870 523076 4922
rect 523132 4870 523142 4922
rect 522822 4868 522836 4870
rect 522892 4868 522916 4870
rect 522972 4868 522996 4870
rect 523052 4868 523076 4870
rect 523132 4868 523156 4870
rect 523212 4868 523236 4870
rect 523292 4868 523316 4870
rect 523372 4868 523386 4870
rect 522822 4848 523386 4868
rect 522822 3836 523386 3856
rect 522822 3834 522836 3836
rect 522892 3834 522916 3836
rect 522972 3834 522996 3836
rect 523052 3834 523076 3836
rect 523132 3834 523156 3836
rect 523212 3834 523236 3836
rect 523292 3834 523316 3836
rect 523372 3834 523386 3836
rect 523066 3782 523076 3834
rect 523132 3782 523142 3834
rect 522822 3780 522836 3782
rect 522892 3780 522916 3782
rect 522972 3780 522996 3782
rect 523052 3780 523076 3782
rect 523132 3780 523156 3782
rect 523212 3780 523236 3782
rect 523292 3780 523316 3782
rect 523372 3780 523386 3782
rect 522822 3760 523386 3780
rect 522822 2748 523386 2768
rect 522822 2746 522836 2748
rect 522892 2746 522916 2748
rect 522972 2746 522996 2748
rect 523052 2746 523076 2748
rect 523132 2746 523156 2748
rect 523212 2746 523236 2748
rect 523292 2746 523316 2748
rect 523372 2746 523386 2748
rect 523066 2694 523076 2746
rect 523132 2694 523142 2746
rect 522822 2692 522836 2694
rect 522892 2692 522916 2694
rect 522972 2692 522996 2694
rect 523052 2692 523076 2694
rect 523132 2692 523156 2694
rect 523212 2692 523236 2694
rect 523292 2692 523316 2694
rect 523372 2692 523386 2694
rect 522822 2672 523386 2692
rect 523880 480 523908 6394
rect 524156 6254 524184 8078
rect 524984 6526 525012 8092
rect 526180 6662 526208 8092
rect 527284 6730 527312 8092
rect 527272 6724 527324 6730
rect 527272 6666 527324 6672
rect 526168 6656 526220 6662
rect 526168 6598 526220 6604
rect 524972 6520 525024 6526
rect 524972 6462 525024 6468
rect 525064 6384 525116 6390
rect 525064 6326 525116 6332
rect 524420 6316 524472 6322
rect 524420 6258 524472 6264
rect 524144 6248 524196 6254
rect 524144 6190 524196 6196
rect 524432 3194 524460 6258
rect 524420 3188 524472 3194
rect 524420 3130 524472 3136
rect 525076 480 525104 6326
rect 528480 6322 528508 8092
rect 529584 6390 529612 8092
rect 530780 6458 530808 8092
rect 531044 6860 531096 6866
rect 531044 6802 531096 6808
rect 530768 6452 530820 6458
rect 530768 6394 530820 6400
rect 529572 6384 529624 6390
rect 529572 6326 529624 6332
rect 528468 6316 528520 6322
rect 528468 6258 528520 6264
rect 527088 6180 527140 6186
rect 527088 6122 527140 6128
rect 525800 5908 525852 5914
rect 525800 5850 525852 5856
rect 525812 3058 525840 5850
rect 527100 3346 527128 6122
rect 529848 3460 529900 3466
rect 529848 3402 529900 3408
rect 527100 3318 527496 3346
rect 526260 3188 526312 3194
rect 526260 3130 526312 3136
rect 525800 3052 525852 3058
rect 525800 2994 525852 3000
rect 526272 480 526300 3130
rect 527468 480 527496 3318
rect 528652 3052 528704 3058
rect 528652 2994 528704 3000
rect 528664 480 528692 2994
rect 529860 480 529888 3402
rect 531056 480 531084 6802
rect 531320 6588 531372 6594
rect 531320 6530 531372 6536
rect 531332 3602 531360 6530
rect 531504 6112 531556 6118
rect 531504 6054 531556 6060
rect 531320 3596 531372 3602
rect 531320 3538 531372 3544
rect 531516 3058 531544 6054
rect 531884 5914 531912 8092
rect 532240 6792 532292 6798
rect 532240 6734 532292 6740
rect 531872 5908 531924 5914
rect 531872 5850 531924 5856
rect 531504 3052 531556 3058
rect 531504 2994 531556 3000
rect 532252 480 532280 6734
rect 532988 5574 533016 8092
rect 534184 6186 534212 8092
rect 535288 6798 535316 8092
rect 535276 6792 535328 6798
rect 535276 6734 535328 6740
rect 536484 6254 536512 8092
rect 537588 6526 537616 8092
rect 538784 6866 538812 8092
rect 538772 6860 538824 6866
rect 538772 6802 538824 6808
rect 539324 6724 539376 6730
rect 539324 6666 539376 6672
rect 538128 6656 538180 6662
rect 538128 6598 538180 6604
rect 536748 6520 536800 6526
rect 536748 6462 536800 6468
rect 537576 6520 537628 6526
rect 537576 6462 537628 6468
rect 535368 6248 535420 6254
rect 535368 6190 535420 6196
rect 536472 6248 536524 6254
rect 536472 6190 536524 6196
rect 534172 6180 534224 6186
rect 534172 6122 534224 6128
rect 532976 5568 533028 5574
rect 532976 5510 533028 5516
rect 533436 3596 533488 3602
rect 533436 3538 533488 3544
rect 533448 480 533476 3538
rect 535380 3210 535408 6190
rect 535460 5568 535512 5574
rect 535460 5510 535512 5516
rect 535472 3466 535500 5510
rect 535460 3460 535512 3466
rect 535460 3402 535512 3408
rect 536760 3346 536788 6462
rect 536760 3318 536972 3346
rect 535380 3182 535776 3210
rect 534540 3052 534592 3058
rect 534540 2994 534592 3000
rect 534552 480 534580 2994
rect 535748 480 535776 3182
rect 536944 480 536972 3318
rect 538140 480 538168 6598
rect 539336 480 539364 6666
rect 539888 6322 539916 8092
rect 541084 6662 541112 8092
rect 541072 6656 541124 6662
rect 541072 6598 541124 6604
rect 541532 6452 541584 6458
rect 541532 6394 541584 6400
rect 539968 6384 540020 6390
rect 539968 6326 540020 6332
rect 539416 6316 539468 6322
rect 539416 6258 539468 6264
rect 539876 6316 539928 6322
rect 539876 6258 539928 6264
rect 539428 4146 539456 6258
rect 539416 4140 539468 4146
rect 539416 4082 539468 4088
rect 539980 3126 540008 6326
rect 541440 5908 541492 5914
rect 541440 5850 541492 5856
rect 540822 5468 541386 5488
rect 540822 5466 540836 5468
rect 540892 5466 540916 5468
rect 540972 5466 540996 5468
rect 541052 5466 541076 5468
rect 541132 5466 541156 5468
rect 541212 5466 541236 5468
rect 541292 5466 541316 5468
rect 541372 5466 541386 5468
rect 541066 5414 541076 5466
rect 541132 5414 541142 5466
rect 540822 5412 540836 5414
rect 540892 5412 540916 5414
rect 540972 5412 540996 5414
rect 541052 5412 541076 5414
rect 541132 5412 541156 5414
rect 541212 5412 541236 5414
rect 541292 5412 541316 5414
rect 541372 5412 541386 5414
rect 540822 5392 541386 5412
rect 540822 4380 541386 4400
rect 540822 4378 540836 4380
rect 540892 4378 540916 4380
rect 540972 4378 540996 4380
rect 541052 4378 541076 4380
rect 541132 4378 541156 4380
rect 541212 4378 541236 4380
rect 541292 4378 541316 4380
rect 541372 4378 541386 4380
rect 541066 4326 541076 4378
rect 541132 4326 541142 4378
rect 540822 4324 540836 4326
rect 540892 4324 540916 4326
rect 540972 4324 540996 4326
rect 541052 4324 541076 4326
rect 541132 4324 541156 4326
rect 541212 4324 541236 4326
rect 541292 4324 541316 4326
rect 541372 4324 541386 4326
rect 540822 4304 541386 4324
rect 540520 4140 540572 4146
rect 540520 4082 540572 4088
rect 539968 3120 540020 3126
rect 539968 3062 540020 3068
rect 540532 480 540560 4082
rect 540822 3292 541386 3312
rect 540822 3290 540836 3292
rect 540892 3290 540916 3292
rect 540972 3290 540996 3292
rect 541052 3290 541076 3292
rect 541132 3290 541156 3292
rect 541212 3290 541236 3292
rect 541292 3290 541316 3292
rect 541372 3290 541386 3292
rect 541066 3238 541076 3290
rect 541132 3238 541142 3290
rect 540822 3236 540836 3238
rect 540892 3236 540916 3238
rect 540972 3236 540996 3238
rect 541052 3236 541076 3238
rect 541132 3236 541156 3238
rect 541212 3236 541236 3238
rect 541292 3236 541316 3238
rect 541372 3236 541386 3238
rect 540822 3216 541386 3236
rect 541452 3194 541480 5850
rect 541544 3398 541572 6394
rect 542188 6390 542216 8092
rect 543384 6594 543412 8092
rect 543372 6588 543424 6594
rect 543372 6530 543424 6536
rect 544488 6458 544516 8092
rect 545120 6792 545172 6798
rect 545120 6734 545172 6740
rect 544476 6452 544528 6458
rect 544476 6394 544528 6400
rect 542176 6384 542228 6390
rect 542176 6326 542228 6332
rect 545132 3602 545160 6734
rect 545592 6730 545620 8092
rect 546788 6798 546816 8092
rect 546776 6792 546828 6798
rect 546776 6734 546828 6740
rect 545580 6724 545632 6730
rect 545580 6666 545632 6672
rect 546592 6520 546644 6526
rect 546592 6462 546644 6468
rect 546500 6248 546552 6254
rect 546500 6190 546552 6196
rect 546408 6180 546460 6186
rect 546408 6122 546460 6128
rect 546420 4026 546448 6122
rect 546512 4146 546540 6190
rect 546500 4140 546552 4146
rect 546500 4082 546552 4088
rect 546420 3998 546540 4026
rect 545120 3596 545172 3602
rect 545120 3538 545172 3544
rect 545304 3460 545356 3466
rect 545304 3402 545356 3408
rect 541532 3392 541584 3398
rect 541532 3334 541584 3340
rect 542912 3392 542964 3398
rect 542912 3334 542964 3340
rect 541440 3188 541492 3194
rect 541440 3130 541492 3136
rect 541716 3120 541768 3126
rect 541716 3062 541768 3068
rect 540822 2204 541386 2224
rect 540822 2202 540836 2204
rect 540892 2202 540916 2204
rect 540972 2202 540996 2204
rect 541052 2202 541076 2204
rect 541132 2202 541156 2204
rect 541212 2202 541236 2204
rect 541292 2202 541316 2204
rect 541372 2202 541386 2204
rect 541066 2150 541076 2202
rect 541132 2150 541142 2202
rect 540822 2148 540836 2150
rect 540892 2148 540916 2150
rect 540972 2148 540996 2150
rect 541052 2148 541076 2150
rect 541132 2148 541156 2150
rect 541212 2148 541236 2150
rect 541292 2148 541316 2150
rect 541372 2148 541386 2150
rect 540822 2128 541386 2148
rect 541728 480 541756 3062
rect 542924 480 542952 3334
rect 544108 3188 544160 3194
rect 544108 3130 544160 3136
rect 544120 480 544148 3130
rect 545316 480 545344 3402
rect 546512 480 546540 3998
rect 546604 3466 546632 6462
rect 547892 5642 547920 8092
rect 547880 5636 547932 5642
rect 547880 5578 547932 5584
rect 549088 5574 549116 8092
rect 549536 6860 549588 6866
rect 549536 6802 549588 6808
rect 549076 5568 549128 5574
rect 549076 5510 549128 5516
rect 548892 4140 548944 4146
rect 548892 4082 548944 4088
rect 547696 3596 547748 3602
rect 547696 3538 547748 3544
rect 546592 3460 546644 3466
rect 546592 3402 546644 3408
rect 547708 480 547736 3538
rect 548904 480 548932 4082
rect 549548 3398 549576 6802
rect 550192 6526 550220 8092
rect 550180 6520 550232 6526
rect 550180 6462 550232 6468
rect 550640 6316 550692 6322
rect 550640 6258 550692 6264
rect 550088 3460 550140 3466
rect 550088 3402 550140 3408
rect 549536 3392 549588 3398
rect 549536 3334 549588 3340
rect 550100 480 550128 3402
rect 550652 3194 550680 6258
rect 551388 6254 551416 8092
rect 552020 6384 552072 6390
rect 552020 6326 552072 6332
rect 551376 6248 551428 6254
rect 551376 6190 551428 6196
rect 551928 5636 551980 5642
rect 551928 5578 551980 5584
rect 550732 5568 550784 5574
rect 550732 5510 550784 5516
rect 550744 3466 550772 5510
rect 551940 3534 551968 5578
rect 551928 3528 551980 3534
rect 551928 3470 551980 3476
rect 550732 3460 550784 3466
rect 550732 3402 550784 3408
rect 551192 3392 551244 3398
rect 551192 3334 551244 3340
rect 550640 3188 550692 3194
rect 550640 3130 550692 3136
rect 551204 480 551232 3334
rect 552032 3126 552060 6326
rect 552492 6118 552520 8092
rect 553308 6656 553360 6662
rect 553308 6598 553360 6604
rect 552480 6112 552532 6118
rect 552480 6054 552532 6060
rect 553320 3584 553348 6598
rect 553400 6588 553452 6594
rect 553400 6530 553452 6536
rect 553412 3738 553440 6530
rect 553688 6186 553716 8092
rect 554792 6322 554820 8092
rect 554872 6452 554924 6458
rect 554872 6394 554924 6400
rect 554780 6316 554832 6322
rect 554780 6258 554832 6264
rect 553676 6180 553728 6186
rect 553676 6122 553728 6128
rect 553400 3732 553452 3738
rect 553400 3674 553452 3680
rect 553320 3556 553624 3584
rect 552388 3188 552440 3194
rect 552388 3130 552440 3136
rect 552020 3120 552072 3126
rect 552020 3062 552072 3068
rect 552400 480 552428 3130
rect 553596 480 553624 3556
rect 554884 3194 554912 6394
rect 555896 5914 555924 8092
rect 556160 6792 556212 6798
rect 556160 6734 556212 6740
rect 555884 5908 555936 5914
rect 555884 5850 555936 5856
rect 555976 3732 556028 3738
rect 555976 3674 556028 3680
rect 554872 3188 554924 3194
rect 554872 3130 554924 3136
rect 554780 3120 554832 3126
rect 554780 3062 554832 3068
rect 554792 480 554820 3062
rect 555988 480 556016 3674
rect 556172 3602 556200 6734
rect 556252 6724 556304 6730
rect 556252 6666 556304 6672
rect 556160 3596 556212 3602
rect 556160 3538 556212 3544
rect 556264 3398 556292 6666
rect 557092 6662 557120 8092
rect 558196 6730 558224 8092
rect 558184 6724 558236 6730
rect 558184 6666 558236 6672
rect 557080 6656 557132 6662
rect 557080 6598 557132 6604
rect 559392 6594 559420 8092
rect 560496 6866 560524 8092
rect 560484 6860 560536 6866
rect 560484 6802 560536 6808
rect 561692 6798 561720 8092
rect 561680 6792 561732 6798
rect 561680 6734 561732 6740
rect 559380 6588 559432 6594
rect 559380 6530 559432 6536
rect 560392 6520 560444 6526
rect 560392 6462 560444 6468
rect 558822 6012 559386 6032
rect 558822 6010 558836 6012
rect 558892 6010 558916 6012
rect 558972 6010 558996 6012
rect 559052 6010 559076 6012
rect 559132 6010 559156 6012
rect 559212 6010 559236 6012
rect 559292 6010 559316 6012
rect 559372 6010 559386 6012
rect 559066 5958 559076 6010
rect 559132 5958 559142 6010
rect 558822 5956 558836 5958
rect 558892 5956 558916 5958
rect 558972 5956 558996 5958
rect 559052 5956 559076 5958
rect 559132 5956 559156 5958
rect 559212 5956 559236 5958
rect 559292 5956 559316 5958
rect 559372 5956 559386 5958
rect 558822 5936 559386 5956
rect 558822 4924 559386 4944
rect 558822 4922 558836 4924
rect 558892 4922 558916 4924
rect 558972 4922 558996 4924
rect 559052 4922 559076 4924
rect 559132 4922 559156 4924
rect 559212 4922 559236 4924
rect 559292 4922 559316 4924
rect 559372 4922 559386 4924
rect 559066 4870 559076 4922
rect 559132 4870 559142 4922
rect 558822 4868 558836 4870
rect 558892 4868 558916 4870
rect 558972 4868 558996 4870
rect 559052 4868 559076 4870
rect 559132 4868 559156 4870
rect 559212 4868 559236 4870
rect 559292 4868 559316 4870
rect 559372 4868 559386 4870
rect 558822 4848 559386 4868
rect 558822 3836 559386 3856
rect 558822 3834 558836 3836
rect 558892 3834 558916 3836
rect 558972 3834 558996 3836
rect 559052 3834 559076 3836
rect 559132 3834 559156 3836
rect 559212 3834 559236 3836
rect 559292 3834 559316 3836
rect 559372 3834 559386 3836
rect 559066 3782 559076 3834
rect 559132 3782 559142 3834
rect 558822 3780 558836 3782
rect 558892 3780 558916 3782
rect 558972 3780 558996 3782
rect 559052 3780 559076 3782
rect 559132 3780 559156 3782
rect 559212 3780 559236 3782
rect 559292 3780 559316 3782
rect 559372 3780 559386 3782
rect 558822 3760 559386 3780
rect 559564 3596 559616 3602
rect 559564 3538 559616 3544
rect 556252 3392 556304 3398
rect 556252 3334 556304 3340
rect 558368 3392 558420 3398
rect 558368 3334 558420 3340
rect 557172 3188 557224 3194
rect 557172 3130 557224 3136
rect 557184 480 557212 3130
rect 558380 480 558408 3334
rect 558822 2748 559386 2768
rect 558822 2746 558836 2748
rect 558892 2746 558916 2748
rect 558972 2746 558996 2748
rect 559052 2746 559076 2748
rect 559132 2746 559156 2748
rect 559212 2746 559236 2748
rect 559292 2746 559316 2748
rect 559372 2746 559386 2748
rect 559066 2694 559076 2746
rect 559132 2694 559142 2746
rect 558822 2692 558836 2694
rect 558892 2692 558916 2694
rect 558972 2692 558996 2694
rect 559052 2692 559076 2694
rect 559132 2692 559156 2694
rect 559212 2692 559236 2694
rect 559292 2692 559316 2694
rect 559372 2692 559386 2694
rect 558822 2672 559386 2692
rect 559576 480 559604 3538
rect 560404 3398 560432 6462
rect 562796 6390 562824 8092
rect 563992 6526 564020 8092
rect 563980 6520 564032 6526
rect 563980 6462 564032 6468
rect 565096 6458 565124 8092
rect 565084 6452 565136 6458
rect 565084 6394 565136 6400
rect 562784 6384 562836 6390
rect 562784 6326 562836 6332
rect 566200 6322 566228 8092
rect 564440 6316 564492 6322
rect 564440 6258 564492 6264
rect 566188 6316 566240 6322
rect 566188 6258 566240 6264
rect 561772 6248 561824 6254
rect 561772 6190 561824 6196
rect 561680 6112 561732 6118
rect 561680 6054 561732 6060
rect 560760 3528 560812 3534
rect 560760 3470 560812 3476
rect 560392 3392 560444 3398
rect 560392 3334 560444 3340
rect 560772 480 560800 3470
rect 561692 3194 561720 6054
rect 561680 3188 561732 3194
rect 561680 3130 561732 3136
rect 561784 3126 561812 6190
rect 564452 4078 564480 6258
rect 567396 6254 567424 8092
rect 568212 6724 568264 6730
rect 568212 6666 568264 6672
rect 567384 6248 567436 6254
rect 567384 6190 567436 6196
rect 564624 6180 564676 6186
rect 564624 6122 564676 6128
rect 564532 5908 564584 5914
rect 564532 5850 564584 5856
rect 564440 4072 564492 4078
rect 564440 4014 564492 4020
rect 561956 3460 562008 3466
rect 561956 3402 562008 3408
rect 561772 3120 561824 3126
rect 561772 3062 561824 3068
rect 561968 480 561996 3402
rect 563152 3392 563204 3398
rect 563152 3334 563204 3340
rect 563164 480 563192 3334
rect 564348 3120 564400 3126
rect 564348 3062 564400 3068
rect 564360 480 564388 3062
rect 564544 3058 564572 5850
rect 564636 3126 564664 6122
rect 568224 4146 568252 6666
rect 568396 6656 568448 6662
rect 568396 6598 568448 6604
rect 568212 4140 568264 4146
rect 568212 4082 568264 4088
rect 567844 4072 567896 4078
rect 567844 4014 567896 4020
rect 565544 3188 565596 3194
rect 565544 3130 565596 3136
rect 564624 3120 564676 3126
rect 564624 3062 564676 3068
rect 564532 3052 564584 3058
rect 564532 2994 564584 3000
rect 565556 480 565584 3130
rect 566740 3120 566792 3126
rect 566740 3062 566792 3068
rect 566752 480 566780 3062
rect 567856 480 567884 4014
rect 568408 3466 568436 6598
rect 568500 6186 568528 8092
rect 570144 6860 570196 6866
rect 570144 6802 570196 6808
rect 568488 6180 568540 6186
rect 568488 6122 568540 6128
rect 570156 4078 570184 6802
rect 571340 6792 571392 6798
rect 571340 6734 571392 6740
rect 570144 4072 570196 4078
rect 570144 4014 570196 4020
rect 571352 4010 571380 6734
rect 572628 6588 572680 6594
rect 572628 6530 572680 6536
rect 571432 4140 571484 4146
rect 571432 4082 571484 4088
rect 571340 4004 571392 4010
rect 571340 3946 571392 3952
rect 568396 3460 568448 3466
rect 568396 3402 568448 3408
rect 570236 3460 570288 3466
rect 570236 3402 570288 3408
rect 569040 3052 569092 3058
rect 569040 2994 569092 3000
rect 569052 480 569080 2994
rect 570248 480 570276 3402
rect 571444 480 571472 4082
rect 572640 480 572668 6530
rect 575480 6520 575532 6526
rect 575480 6462 575532 6468
rect 573824 4072 573876 4078
rect 573824 4014 573876 4020
rect 573836 480 573864 4014
rect 575020 4004 575072 4010
rect 575020 3946 575072 3952
rect 575032 480 575060 3946
rect 575492 3194 575520 6462
rect 577688 6452 577740 6458
rect 577688 6394 577740 6400
rect 576216 6384 576268 6390
rect 576216 6326 576268 6332
rect 575480 3188 575532 3194
rect 575480 3130 575532 3136
rect 576228 480 576256 6326
rect 576822 5468 577386 5488
rect 576822 5466 576836 5468
rect 576892 5466 576916 5468
rect 576972 5466 576996 5468
rect 577052 5466 577076 5468
rect 577132 5466 577156 5468
rect 577212 5466 577236 5468
rect 577292 5466 577316 5468
rect 577372 5466 577386 5468
rect 577066 5414 577076 5466
rect 577132 5414 577142 5466
rect 576822 5412 576836 5414
rect 576892 5412 576916 5414
rect 576972 5412 576996 5414
rect 577052 5412 577076 5414
rect 577132 5412 577156 5414
rect 577212 5412 577236 5414
rect 577292 5412 577316 5414
rect 577372 5412 577386 5414
rect 576822 5392 577386 5412
rect 576822 4380 577386 4400
rect 576822 4378 576836 4380
rect 576892 4378 576916 4380
rect 576972 4378 576996 4380
rect 577052 4378 577076 4380
rect 577132 4378 577156 4380
rect 577212 4378 577236 4380
rect 577292 4378 577316 4380
rect 577372 4378 577386 4380
rect 577066 4326 577076 4378
rect 577132 4326 577142 4378
rect 576822 4324 576836 4326
rect 576892 4324 576916 4326
rect 576972 4324 576996 4326
rect 577052 4324 577076 4326
rect 577132 4324 577156 4326
rect 577212 4324 577236 4326
rect 577292 4324 577316 4326
rect 577372 4324 577386 4326
rect 576822 4304 577386 4324
rect 576822 3292 577386 3312
rect 576822 3290 576836 3292
rect 576892 3290 576916 3292
rect 576972 3290 576996 3292
rect 577052 3290 577076 3292
rect 577132 3290 577156 3292
rect 577212 3290 577236 3292
rect 577292 3290 577316 3292
rect 577372 3290 577386 3292
rect 577066 3238 577076 3290
rect 577132 3238 577142 3290
rect 576822 3236 576836 3238
rect 576892 3236 576916 3238
rect 576972 3236 576996 3238
rect 577052 3236 577076 3238
rect 577132 3236 577156 3238
rect 577212 3236 577236 3238
rect 577292 3236 577316 3238
rect 577372 3236 577386 3238
rect 576822 3216 577386 3236
rect 577700 3194 577728 6394
rect 579804 6316 579856 6322
rect 579804 6258 579856 6264
rect 577412 3188 577464 3194
rect 577412 3130 577464 3136
rect 577688 3188 577740 3194
rect 577688 3130 577740 3136
rect 578608 3188 578660 3194
rect 578608 3130 578660 3136
rect 576822 2204 577386 2224
rect 576822 2202 576836 2204
rect 576892 2202 576916 2204
rect 576972 2202 576996 2204
rect 577052 2202 577076 2204
rect 577132 2202 577156 2204
rect 577212 2202 577236 2204
rect 577292 2202 577316 2204
rect 577372 2202 577386 2204
rect 577066 2150 577076 2202
rect 577132 2150 577142 2202
rect 576822 2148 576836 2150
rect 576892 2148 576916 2150
rect 576972 2148 576996 2150
rect 577052 2148 577076 2150
rect 577132 2148 577156 2150
rect 577212 2148 577236 2150
rect 577292 2148 577316 2150
rect 577372 2148 577386 2150
rect 576822 2128 577386 2148
rect 577424 480 577452 3130
rect 578620 480 578648 3130
rect 579816 480 579844 6258
rect 581000 6248 581052 6254
rect 581000 6190 581052 6196
rect 581012 480 581040 6190
rect 582196 6180 582248 6186
rect 582196 6122 582248 6128
rect 582208 480 582236 6122
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 18836 701242 18892 701244
rect 18916 701242 18972 701244
rect 18996 701242 19052 701244
rect 19076 701242 19132 701244
rect 19156 701242 19212 701244
rect 19236 701242 19292 701244
rect 19316 701242 19372 701244
rect 18836 701190 18874 701242
rect 18874 701190 18886 701242
rect 18886 701190 18892 701242
rect 18916 701190 18938 701242
rect 18938 701190 18950 701242
rect 18950 701190 18972 701242
rect 18996 701190 19002 701242
rect 19002 701190 19014 701242
rect 19014 701190 19052 701242
rect 19076 701190 19078 701242
rect 19078 701190 19130 701242
rect 19130 701190 19132 701242
rect 19156 701190 19194 701242
rect 19194 701190 19206 701242
rect 19206 701190 19212 701242
rect 19236 701190 19258 701242
rect 19258 701190 19270 701242
rect 19270 701190 19292 701242
rect 19316 701190 19322 701242
rect 19322 701190 19334 701242
rect 19334 701190 19372 701242
rect 18836 701188 18892 701190
rect 18916 701188 18972 701190
rect 18996 701188 19052 701190
rect 19076 701188 19132 701190
rect 19156 701188 19212 701190
rect 19236 701188 19292 701190
rect 19316 701188 19372 701190
rect 36836 701786 36892 701788
rect 36916 701786 36972 701788
rect 36996 701786 37052 701788
rect 37076 701786 37132 701788
rect 37156 701786 37212 701788
rect 37236 701786 37292 701788
rect 37316 701786 37372 701788
rect 36836 701734 36874 701786
rect 36874 701734 36886 701786
rect 36886 701734 36892 701786
rect 36916 701734 36938 701786
rect 36938 701734 36950 701786
rect 36950 701734 36972 701786
rect 36996 701734 37002 701786
rect 37002 701734 37014 701786
rect 37014 701734 37052 701786
rect 37076 701734 37078 701786
rect 37078 701734 37130 701786
rect 37130 701734 37132 701786
rect 37156 701734 37194 701786
rect 37194 701734 37206 701786
rect 37206 701734 37212 701786
rect 37236 701734 37258 701786
rect 37258 701734 37270 701786
rect 37270 701734 37292 701786
rect 37316 701734 37322 701786
rect 37322 701734 37334 701786
rect 37334 701734 37372 701786
rect 36836 701732 36892 701734
rect 36916 701732 36972 701734
rect 36996 701732 37052 701734
rect 37076 701732 37132 701734
rect 37156 701732 37212 701734
rect 37236 701732 37292 701734
rect 37316 701732 37372 701734
rect 54836 701242 54892 701244
rect 54916 701242 54972 701244
rect 54996 701242 55052 701244
rect 55076 701242 55132 701244
rect 55156 701242 55212 701244
rect 55236 701242 55292 701244
rect 55316 701242 55372 701244
rect 54836 701190 54874 701242
rect 54874 701190 54886 701242
rect 54886 701190 54892 701242
rect 54916 701190 54938 701242
rect 54938 701190 54950 701242
rect 54950 701190 54972 701242
rect 54996 701190 55002 701242
rect 55002 701190 55014 701242
rect 55014 701190 55052 701242
rect 55076 701190 55078 701242
rect 55078 701190 55130 701242
rect 55130 701190 55132 701242
rect 55156 701190 55194 701242
rect 55194 701190 55206 701242
rect 55206 701190 55212 701242
rect 55236 701190 55258 701242
rect 55258 701190 55270 701242
rect 55270 701190 55292 701242
rect 55316 701190 55322 701242
rect 55322 701190 55334 701242
rect 55334 701190 55372 701242
rect 54836 701188 54892 701190
rect 54916 701188 54972 701190
rect 54996 701188 55052 701190
rect 55076 701188 55132 701190
rect 55156 701188 55212 701190
rect 55236 701188 55292 701190
rect 55316 701188 55372 701190
rect 40498 700984 40554 701040
rect 36836 700698 36892 700700
rect 36916 700698 36972 700700
rect 36996 700698 37052 700700
rect 37076 700698 37132 700700
rect 37156 700698 37212 700700
rect 37236 700698 37292 700700
rect 37316 700698 37372 700700
rect 36836 700646 36874 700698
rect 36874 700646 36886 700698
rect 36886 700646 36892 700698
rect 36916 700646 36938 700698
rect 36938 700646 36950 700698
rect 36950 700646 36972 700698
rect 36996 700646 37002 700698
rect 37002 700646 37014 700698
rect 37014 700646 37052 700698
rect 37076 700646 37078 700698
rect 37078 700646 37130 700698
rect 37130 700646 37132 700698
rect 37156 700646 37194 700698
rect 37194 700646 37206 700698
rect 37206 700646 37212 700698
rect 37236 700646 37258 700698
rect 37258 700646 37270 700698
rect 37270 700646 37292 700698
rect 37316 700646 37322 700698
rect 37322 700646 37334 700698
rect 37334 700646 37372 700698
rect 36836 700644 36892 700646
rect 36916 700644 36972 700646
rect 36996 700644 37052 700646
rect 37076 700644 37132 700646
rect 37156 700644 37212 700646
rect 37236 700644 37292 700646
rect 37316 700644 37372 700646
rect 24306 700440 24362 700496
rect 8114 700304 8170 700360
rect 72836 701786 72892 701788
rect 72916 701786 72972 701788
rect 72996 701786 73052 701788
rect 73076 701786 73132 701788
rect 73156 701786 73212 701788
rect 73236 701786 73292 701788
rect 73316 701786 73372 701788
rect 72836 701734 72874 701786
rect 72874 701734 72886 701786
rect 72886 701734 72892 701786
rect 72916 701734 72938 701786
rect 72938 701734 72950 701786
rect 72950 701734 72972 701786
rect 72996 701734 73002 701786
rect 73002 701734 73014 701786
rect 73014 701734 73052 701786
rect 73076 701734 73078 701786
rect 73078 701734 73130 701786
rect 73130 701734 73132 701786
rect 73156 701734 73194 701786
rect 73194 701734 73206 701786
rect 73206 701734 73212 701786
rect 73236 701734 73258 701786
rect 73258 701734 73270 701786
rect 73270 701734 73292 701786
rect 73316 701734 73322 701786
rect 73322 701734 73334 701786
rect 73334 701734 73372 701786
rect 72836 701732 72892 701734
rect 72916 701732 72972 701734
rect 72996 701732 73052 701734
rect 73076 701732 73132 701734
rect 73156 701732 73212 701734
rect 73236 701732 73292 701734
rect 73316 701732 73372 701734
rect 72836 700698 72892 700700
rect 72916 700698 72972 700700
rect 72996 700698 73052 700700
rect 73076 700698 73132 700700
rect 73156 700698 73212 700700
rect 73236 700698 73292 700700
rect 73316 700698 73372 700700
rect 72836 700646 72874 700698
rect 72874 700646 72886 700698
rect 72886 700646 72892 700698
rect 72916 700646 72938 700698
rect 72938 700646 72950 700698
rect 72950 700646 72972 700698
rect 72996 700646 73002 700698
rect 73002 700646 73014 700698
rect 73014 700646 73052 700698
rect 73076 700646 73078 700698
rect 73078 700646 73130 700698
rect 73130 700646 73132 700698
rect 73156 700646 73194 700698
rect 73194 700646 73206 700698
rect 73206 700646 73212 700698
rect 73236 700646 73258 700698
rect 73258 700646 73270 700698
rect 73270 700646 73292 700698
rect 73316 700646 73322 700698
rect 73322 700646 73334 700698
rect 73334 700646 73372 700698
rect 72836 700644 72892 700646
rect 72916 700644 72972 700646
rect 72996 700644 73052 700646
rect 73076 700644 73132 700646
rect 73156 700644 73212 700646
rect 73236 700644 73292 700646
rect 73316 700644 73372 700646
rect 90836 701242 90892 701244
rect 90916 701242 90972 701244
rect 90996 701242 91052 701244
rect 91076 701242 91132 701244
rect 91156 701242 91212 701244
rect 91236 701242 91292 701244
rect 91316 701242 91372 701244
rect 90836 701190 90874 701242
rect 90874 701190 90886 701242
rect 90886 701190 90892 701242
rect 90916 701190 90938 701242
rect 90938 701190 90950 701242
rect 90950 701190 90972 701242
rect 90996 701190 91002 701242
rect 91002 701190 91014 701242
rect 91014 701190 91052 701242
rect 91076 701190 91078 701242
rect 91078 701190 91130 701242
rect 91130 701190 91132 701242
rect 91156 701190 91194 701242
rect 91194 701190 91206 701242
rect 91206 701190 91212 701242
rect 91236 701190 91258 701242
rect 91258 701190 91270 701242
rect 91270 701190 91292 701242
rect 91316 701190 91322 701242
rect 91322 701190 91334 701242
rect 91334 701190 91372 701242
rect 90836 701188 90892 701190
rect 90916 701188 90972 701190
rect 90996 701188 91052 701190
rect 91076 701188 91132 701190
rect 91156 701188 91212 701190
rect 91236 701188 91292 701190
rect 91316 701188 91372 701190
rect 108836 701786 108892 701788
rect 108916 701786 108972 701788
rect 108996 701786 109052 701788
rect 109076 701786 109132 701788
rect 109156 701786 109212 701788
rect 109236 701786 109292 701788
rect 109316 701786 109372 701788
rect 108836 701734 108874 701786
rect 108874 701734 108886 701786
rect 108886 701734 108892 701786
rect 108916 701734 108938 701786
rect 108938 701734 108950 701786
rect 108950 701734 108972 701786
rect 108996 701734 109002 701786
rect 109002 701734 109014 701786
rect 109014 701734 109052 701786
rect 109076 701734 109078 701786
rect 109078 701734 109130 701786
rect 109130 701734 109132 701786
rect 109156 701734 109194 701786
rect 109194 701734 109206 701786
rect 109206 701734 109212 701786
rect 109236 701734 109258 701786
rect 109258 701734 109270 701786
rect 109270 701734 109292 701786
rect 109316 701734 109322 701786
rect 109322 701734 109334 701786
rect 109334 701734 109372 701786
rect 108836 701732 108892 701734
rect 108916 701732 108972 701734
rect 108996 701732 109052 701734
rect 109076 701732 109132 701734
rect 109156 701732 109212 701734
rect 109236 701732 109292 701734
rect 109316 701732 109372 701734
rect 126836 701242 126892 701244
rect 126916 701242 126972 701244
rect 126996 701242 127052 701244
rect 127076 701242 127132 701244
rect 127156 701242 127212 701244
rect 127236 701242 127292 701244
rect 127316 701242 127372 701244
rect 126836 701190 126874 701242
rect 126874 701190 126886 701242
rect 126886 701190 126892 701242
rect 126916 701190 126938 701242
rect 126938 701190 126950 701242
rect 126950 701190 126972 701242
rect 126996 701190 127002 701242
rect 127002 701190 127014 701242
rect 127014 701190 127052 701242
rect 127076 701190 127078 701242
rect 127078 701190 127130 701242
rect 127130 701190 127132 701242
rect 127156 701190 127194 701242
rect 127194 701190 127206 701242
rect 127206 701190 127212 701242
rect 127236 701190 127258 701242
rect 127258 701190 127270 701242
rect 127270 701190 127292 701242
rect 127316 701190 127322 701242
rect 127322 701190 127334 701242
rect 127334 701190 127372 701242
rect 126836 701188 126892 701190
rect 126916 701188 126972 701190
rect 126996 701188 127052 701190
rect 127076 701188 127132 701190
rect 127156 701188 127212 701190
rect 127236 701188 127292 701190
rect 127316 701188 127372 701190
rect 144836 701786 144892 701788
rect 144916 701786 144972 701788
rect 144996 701786 145052 701788
rect 145076 701786 145132 701788
rect 145156 701786 145212 701788
rect 145236 701786 145292 701788
rect 145316 701786 145372 701788
rect 144836 701734 144874 701786
rect 144874 701734 144886 701786
rect 144886 701734 144892 701786
rect 144916 701734 144938 701786
rect 144938 701734 144950 701786
rect 144950 701734 144972 701786
rect 144996 701734 145002 701786
rect 145002 701734 145014 701786
rect 145014 701734 145052 701786
rect 145076 701734 145078 701786
rect 145078 701734 145130 701786
rect 145130 701734 145132 701786
rect 145156 701734 145194 701786
rect 145194 701734 145206 701786
rect 145206 701734 145212 701786
rect 145236 701734 145258 701786
rect 145258 701734 145270 701786
rect 145270 701734 145292 701786
rect 145316 701734 145322 701786
rect 145322 701734 145334 701786
rect 145334 701734 145372 701786
rect 144836 701732 144892 701734
rect 144916 701732 144972 701734
rect 144996 701732 145052 701734
rect 145076 701732 145132 701734
rect 145156 701732 145212 701734
rect 145236 701732 145292 701734
rect 145316 701732 145372 701734
rect 162836 701242 162892 701244
rect 162916 701242 162972 701244
rect 162996 701242 163052 701244
rect 163076 701242 163132 701244
rect 163156 701242 163212 701244
rect 163236 701242 163292 701244
rect 163316 701242 163372 701244
rect 162836 701190 162874 701242
rect 162874 701190 162886 701242
rect 162886 701190 162892 701242
rect 162916 701190 162938 701242
rect 162938 701190 162950 701242
rect 162950 701190 162972 701242
rect 162996 701190 163002 701242
rect 163002 701190 163014 701242
rect 163014 701190 163052 701242
rect 163076 701190 163078 701242
rect 163078 701190 163130 701242
rect 163130 701190 163132 701242
rect 163156 701190 163194 701242
rect 163194 701190 163206 701242
rect 163206 701190 163212 701242
rect 163236 701190 163258 701242
rect 163258 701190 163270 701242
rect 163270 701190 163292 701242
rect 163316 701190 163322 701242
rect 163322 701190 163334 701242
rect 163334 701190 163372 701242
rect 162836 701188 162892 701190
rect 162916 701188 162972 701190
rect 162996 701188 163052 701190
rect 163076 701188 163132 701190
rect 163156 701188 163212 701190
rect 163236 701188 163292 701190
rect 163316 701188 163372 701190
rect 108836 700698 108892 700700
rect 108916 700698 108972 700700
rect 108996 700698 109052 700700
rect 109076 700698 109132 700700
rect 109156 700698 109212 700700
rect 109236 700698 109292 700700
rect 109316 700698 109372 700700
rect 108836 700646 108874 700698
rect 108874 700646 108886 700698
rect 108886 700646 108892 700698
rect 108916 700646 108938 700698
rect 108938 700646 108950 700698
rect 108950 700646 108972 700698
rect 108996 700646 109002 700698
rect 109002 700646 109014 700698
rect 109014 700646 109052 700698
rect 109076 700646 109078 700698
rect 109078 700646 109130 700698
rect 109130 700646 109132 700698
rect 109156 700646 109194 700698
rect 109194 700646 109206 700698
rect 109206 700646 109212 700698
rect 109236 700646 109258 700698
rect 109258 700646 109270 700698
rect 109270 700646 109292 700698
rect 109316 700646 109322 700698
rect 109322 700646 109334 700698
rect 109334 700646 109372 700698
rect 108836 700644 108892 700646
rect 108916 700644 108972 700646
rect 108996 700644 109052 700646
rect 109076 700644 109132 700646
rect 109156 700644 109212 700646
rect 109236 700644 109292 700646
rect 109316 700644 109372 700646
rect 144836 700698 144892 700700
rect 144916 700698 144972 700700
rect 144996 700698 145052 700700
rect 145076 700698 145132 700700
rect 145156 700698 145212 700700
rect 145236 700698 145292 700700
rect 145316 700698 145372 700700
rect 144836 700646 144874 700698
rect 144874 700646 144886 700698
rect 144886 700646 144892 700698
rect 144916 700646 144938 700698
rect 144938 700646 144950 700698
rect 144950 700646 144972 700698
rect 144996 700646 145002 700698
rect 145002 700646 145014 700698
rect 145014 700646 145052 700698
rect 145076 700646 145078 700698
rect 145078 700646 145130 700698
rect 145130 700646 145132 700698
rect 145156 700646 145194 700698
rect 145194 700646 145206 700698
rect 145206 700646 145212 700698
rect 145236 700646 145258 700698
rect 145258 700646 145270 700698
rect 145270 700646 145292 700698
rect 145316 700646 145322 700698
rect 145322 700646 145334 700698
rect 145334 700646 145372 700698
rect 144836 700644 144892 700646
rect 144916 700644 144972 700646
rect 144996 700644 145052 700646
rect 145076 700644 145132 700646
rect 145156 700644 145212 700646
rect 145236 700644 145292 700646
rect 145316 700644 145372 700646
rect 180836 701786 180892 701788
rect 180916 701786 180972 701788
rect 180996 701786 181052 701788
rect 181076 701786 181132 701788
rect 181156 701786 181212 701788
rect 181236 701786 181292 701788
rect 181316 701786 181372 701788
rect 180836 701734 180874 701786
rect 180874 701734 180886 701786
rect 180886 701734 180892 701786
rect 180916 701734 180938 701786
rect 180938 701734 180950 701786
rect 180950 701734 180972 701786
rect 180996 701734 181002 701786
rect 181002 701734 181014 701786
rect 181014 701734 181052 701786
rect 181076 701734 181078 701786
rect 181078 701734 181130 701786
rect 181130 701734 181132 701786
rect 181156 701734 181194 701786
rect 181194 701734 181206 701786
rect 181206 701734 181212 701786
rect 181236 701734 181258 701786
rect 181258 701734 181270 701786
rect 181270 701734 181292 701786
rect 181316 701734 181322 701786
rect 181322 701734 181334 701786
rect 181334 701734 181372 701786
rect 180836 701732 180892 701734
rect 180916 701732 180972 701734
rect 180996 701732 181052 701734
rect 181076 701732 181132 701734
rect 181156 701732 181212 701734
rect 181236 701732 181292 701734
rect 181316 701732 181372 701734
rect 198836 701242 198892 701244
rect 198916 701242 198972 701244
rect 198996 701242 199052 701244
rect 199076 701242 199132 701244
rect 199156 701242 199212 701244
rect 199236 701242 199292 701244
rect 199316 701242 199372 701244
rect 198836 701190 198874 701242
rect 198874 701190 198886 701242
rect 198886 701190 198892 701242
rect 198916 701190 198938 701242
rect 198938 701190 198950 701242
rect 198950 701190 198972 701242
rect 198996 701190 199002 701242
rect 199002 701190 199014 701242
rect 199014 701190 199052 701242
rect 199076 701190 199078 701242
rect 199078 701190 199130 701242
rect 199130 701190 199132 701242
rect 199156 701190 199194 701242
rect 199194 701190 199206 701242
rect 199206 701190 199212 701242
rect 199236 701190 199258 701242
rect 199258 701190 199270 701242
rect 199270 701190 199292 701242
rect 199316 701190 199322 701242
rect 199322 701190 199334 701242
rect 199334 701190 199372 701242
rect 198836 701188 198892 701190
rect 198916 701188 198972 701190
rect 198996 701188 199052 701190
rect 199076 701188 199132 701190
rect 199156 701188 199212 701190
rect 199236 701188 199292 701190
rect 199316 701188 199372 701190
rect 180836 700698 180892 700700
rect 180916 700698 180972 700700
rect 180996 700698 181052 700700
rect 181076 700698 181132 700700
rect 181156 700698 181212 700700
rect 181236 700698 181292 700700
rect 181316 700698 181372 700700
rect 180836 700646 180874 700698
rect 180874 700646 180886 700698
rect 180886 700646 180892 700698
rect 180916 700646 180938 700698
rect 180938 700646 180950 700698
rect 180950 700646 180972 700698
rect 180996 700646 181002 700698
rect 181002 700646 181014 700698
rect 181014 700646 181052 700698
rect 181076 700646 181078 700698
rect 181078 700646 181130 700698
rect 181130 700646 181132 700698
rect 181156 700646 181194 700698
rect 181194 700646 181206 700698
rect 181206 700646 181212 700698
rect 181236 700646 181258 700698
rect 181258 700646 181270 700698
rect 181270 700646 181292 700698
rect 181316 700646 181322 700698
rect 181322 700646 181334 700698
rect 181334 700646 181372 700698
rect 180836 700644 180892 700646
rect 180916 700644 180972 700646
rect 180996 700644 181052 700646
rect 181076 700644 181132 700646
rect 181156 700644 181212 700646
rect 181236 700644 181292 700646
rect 181316 700644 181372 700646
rect 216836 701786 216892 701788
rect 216916 701786 216972 701788
rect 216996 701786 217052 701788
rect 217076 701786 217132 701788
rect 217156 701786 217212 701788
rect 217236 701786 217292 701788
rect 217316 701786 217372 701788
rect 216836 701734 216874 701786
rect 216874 701734 216886 701786
rect 216886 701734 216892 701786
rect 216916 701734 216938 701786
rect 216938 701734 216950 701786
rect 216950 701734 216972 701786
rect 216996 701734 217002 701786
rect 217002 701734 217014 701786
rect 217014 701734 217052 701786
rect 217076 701734 217078 701786
rect 217078 701734 217130 701786
rect 217130 701734 217132 701786
rect 217156 701734 217194 701786
rect 217194 701734 217206 701786
rect 217206 701734 217212 701786
rect 217236 701734 217258 701786
rect 217258 701734 217270 701786
rect 217270 701734 217292 701786
rect 217316 701734 217322 701786
rect 217322 701734 217334 701786
rect 217334 701734 217372 701786
rect 216836 701732 216892 701734
rect 216916 701732 216972 701734
rect 216996 701732 217052 701734
rect 217076 701732 217132 701734
rect 217156 701732 217212 701734
rect 217236 701732 217292 701734
rect 217316 701732 217372 701734
rect 216836 700698 216892 700700
rect 216916 700698 216972 700700
rect 216996 700698 217052 700700
rect 217076 700698 217132 700700
rect 217156 700698 217212 700700
rect 217236 700698 217292 700700
rect 217316 700698 217372 700700
rect 216836 700646 216874 700698
rect 216874 700646 216886 700698
rect 216886 700646 216892 700698
rect 216916 700646 216938 700698
rect 216938 700646 216950 700698
rect 216950 700646 216972 700698
rect 216996 700646 217002 700698
rect 217002 700646 217014 700698
rect 217014 700646 217052 700698
rect 217076 700646 217078 700698
rect 217078 700646 217130 700698
rect 217130 700646 217132 700698
rect 217156 700646 217194 700698
rect 217194 700646 217206 700698
rect 217206 700646 217212 700698
rect 217236 700646 217258 700698
rect 217258 700646 217270 700698
rect 217270 700646 217292 700698
rect 217316 700646 217322 700698
rect 217322 700646 217334 700698
rect 217334 700646 217372 700698
rect 216836 700644 216892 700646
rect 216916 700644 216972 700646
rect 216996 700644 217052 700646
rect 217076 700644 217132 700646
rect 217156 700644 217212 700646
rect 217236 700644 217292 700646
rect 217316 700644 217372 700646
rect 18836 700154 18892 700156
rect 18916 700154 18972 700156
rect 18996 700154 19052 700156
rect 19076 700154 19132 700156
rect 19156 700154 19212 700156
rect 19236 700154 19292 700156
rect 19316 700154 19372 700156
rect 18836 700102 18874 700154
rect 18874 700102 18886 700154
rect 18886 700102 18892 700154
rect 18916 700102 18938 700154
rect 18938 700102 18950 700154
rect 18950 700102 18972 700154
rect 18996 700102 19002 700154
rect 19002 700102 19014 700154
rect 19014 700102 19052 700154
rect 19076 700102 19078 700154
rect 19078 700102 19130 700154
rect 19130 700102 19132 700154
rect 19156 700102 19194 700154
rect 19194 700102 19206 700154
rect 19206 700102 19212 700154
rect 19236 700102 19258 700154
rect 19258 700102 19270 700154
rect 19270 700102 19292 700154
rect 19316 700102 19322 700154
rect 19322 700102 19334 700154
rect 19334 700102 19372 700154
rect 18836 700100 18892 700102
rect 18916 700100 18972 700102
rect 18996 700100 19052 700102
rect 19076 700100 19132 700102
rect 19156 700100 19212 700102
rect 19236 700100 19292 700102
rect 19316 700100 19372 700102
rect 54836 700154 54892 700156
rect 54916 700154 54972 700156
rect 54996 700154 55052 700156
rect 55076 700154 55132 700156
rect 55156 700154 55212 700156
rect 55236 700154 55292 700156
rect 55316 700154 55372 700156
rect 54836 700102 54874 700154
rect 54874 700102 54886 700154
rect 54886 700102 54892 700154
rect 54916 700102 54938 700154
rect 54938 700102 54950 700154
rect 54950 700102 54972 700154
rect 54996 700102 55002 700154
rect 55002 700102 55014 700154
rect 55014 700102 55052 700154
rect 55076 700102 55078 700154
rect 55078 700102 55130 700154
rect 55130 700102 55132 700154
rect 55156 700102 55194 700154
rect 55194 700102 55206 700154
rect 55206 700102 55212 700154
rect 55236 700102 55258 700154
rect 55258 700102 55270 700154
rect 55270 700102 55292 700154
rect 55316 700102 55322 700154
rect 55322 700102 55334 700154
rect 55334 700102 55372 700154
rect 54836 700100 54892 700102
rect 54916 700100 54972 700102
rect 54996 700100 55052 700102
rect 55076 700100 55132 700102
rect 55156 700100 55212 700102
rect 55236 700100 55292 700102
rect 55316 700100 55372 700102
rect 90836 700154 90892 700156
rect 90916 700154 90972 700156
rect 90996 700154 91052 700156
rect 91076 700154 91132 700156
rect 91156 700154 91212 700156
rect 91236 700154 91292 700156
rect 91316 700154 91372 700156
rect 90836 700102 90874 700154
rect 90874 700102 90886 700154
rect 90886 700102 90892 700154
rect 90916 700102 90938 700154
rect 90938 700102 90950 700154
rect 90950 700102 90972 700154
rect 90996 700102 91002 700154
rect 91002 700102 91014 700154
rect 91014 700102 91052 700154
rect 91076 700102 91078 700154
rect 91078 700102 91130 700154
rect 91130 700102 91132 700154
rect 91156 700102 91194 700154
rect 91194 700102 91206 700154
rect 91206 700102 91212 700154
rect 91236 700102 91258 700154
rect 91258 700102 91270 700154
rect 91270 700102 91292 700154
rect 91316 700102 91322 700154
rect 91322 700102 91334 700154
rect 91334 700102 91372 700154
rect 90836 700100 90892 700102
rect 90916 700100 90972 700102
rect 90996 700100 91052 700102
rect 91076 700100 91132 700102
rect 91156 700100 91212 700102
rect 91236 700100 91292 700102
rect 91316 700100 91372 700102
rect 126836 700154 126892 700156
rect 126916 700154 126972 700156
rect 126996 700154 127052 700156
rect 127076 700154 127132 700156
rect 127156 700154 127212 700156
rect 127236 700154 127292 700156
rect 127316 700154 127372 700156
rect 126836 700102 126874 700154
rect 126874 700102 126886 700154
rect 126886 700102 126892 700154
rect 126916 700102 126938 700154
rect 126938 700102 126950 700154
rect 126950 700102 126972 700154
rect 126996 700102 127002 700154
rect 127002 700102 127014 700154
rect 127014 700102 127052 700154
rect 127076 700102 127078 700154
rect 127078 700102 127130 700154
rect 127130 700102 127132 700154
rect 127156 700102 127194 700154
rect 127194 700102 127206 700154
rect 127206 700102 127212 700154
rect 127236 700102 127258 700154
rect 127258 700102 127270 700154
rect 127270 700102 127292 700154
rect 127316 700102 127322 700154
rect 127322 700102 127334 700154
rect 127334 700102 127372 700154
rect 126836 700100 126892 700102
rect 126916 700100 126972 700102
rect 126996 700100 127052 700102
rect 127076 700100 127132 700102
rect 127156 700100 127212 700102
rect 127236 700100 127292 700102
rect 127316 700100 127372 700102
rect 162836 700154 162892 700156
rect 162916 700154 162972 700156
rect 162996 700154 163052 700156
rect 163076 700154 163132 700156
rect 163156 700154 163212 700156
rect 163236 700154 163292 700156
rect 163316 700154 163372 700156
rect 162836 700102 162874 700154
rect 162874 700102 162886 700154
rect 162886 700102 162892 700154
rect 162916 700102 162938 700154
rect 162938 700102 162950 700154
rect 162950 700102 162972 700154
rect 162996 700102 163002 700154
rect 163002 700102 163014 700154
rect 163014 700102 163052 700154
rect 163076 700102 163078 700154
rect 163078 700102 163130 700154
rect 163130 700102 163132 700154
rect 163156 700102 163194 700154
rect 163194 700102 163206 700154
rect 163206 700102 163212 700154
rect 163236 700102 163258 700154
rect 163258 700102 163270 700154
rect 163270 700102 163292 700154
rect 163316 700102 163322 700154
rect 163322 700102 163334 700154
rect 163334 700102 163372 700154
rect 162836 700100 162892 700102
rect 162916 700100 162972 700102
rect 162996 700100 163052 700102
rect 163076 700100 163132 700102
rect 163156 700100 163212 700102
rect 163236 700100 163292 700102
rect 163316 700100 163372 700102
rect 198836 700154 198892 700156
rect 198916 700154 198972 700156
rect 198996 700154 199052 700156
rect 199076 700154 199132 700156
rect 199156 700154 199212 700156
rect 199236 700154 199292 700156
rect 199316 700154 199372 700156
rect 198836 700102 198874 700154
rect 198874 700102 198886 700154
rect 198886 700102 198892 700154
rect 198916 700102 198938 700154
rect 198938 700102 198950 700154
rect 198950 700102 198972 700154
rect 198996 700102 199002 700154
rect 199002 700102 199014 700154
rect 199014 700102 199052 700154
rect 199076 700102 199078 700154
rect 199078 700102 199130 700154
rect 199130 700102 199132 700154
rect 199156 700102 199194 700154
rect 199194 700102 199206 700154
rect 199206 700102 199212 700154
rect 199236 700102 199258 700154
rect 199258 700102 199270 700154
rect 199270 700102 199292 700154
rect 199316 700102 199322 700154
rect 199322 700102 199334 700154
rect 199334 700102 199372 700154
rect 198836 700100 198892 700102
rect 198916 700100 198972 700102
rect 198996 700100 199052 700102
rect 199076 700100 199132 700102
rect 199156 700100 199212 700102
rect 199236 700100 199292 700102
rect 199316 700100 199372 700102
rect 36836 699610 36892 699612
rect 36916 699610 36972 699612
rect 36996 699610 37052 699612
rect 37076 699610 37132 699612
rect 37156 699610 37212 699612
rect 37236 699610 37292 699612
rect 37316 699610 37372 699612
rect 36836 699558 36874 699610
rect 36874 699558 36886 699610
rect 36886 699558 36892 699610
rect 36916 699558 36938 699610
rect 36938 699558 36950 699610
rect 36950 699558 36972 699610
rect 36996 699558 37002 699610
rect 37002 699558 37014 699610
rect 37014 699558 37052 699610
rect 37076 699558 37078 699610
rect 37078 699558 37130 699610
rect 37130 699558 37132 699610
rect 37156 699558 37194 699610
rect 37194 699558 37206 699610
rect 37206 699558 37212 699610
rect 37236 699558 37258 699610
rect 37258 699558 37270 699610
rect 37270 699558 37292 699610
rect 37316 699558 37322 699610
rect 37322 699558 37334 699610
rect 37334 699558 37372 699610
rect 36836 699556 36892 699558
rect 36916 699556 36972 699558
rect 36996 699556 37052 699558
rect 37076 699556 37132 699558
rect 37156 699556 37212 699558
rect 37236 699556 37292 699558
rect 37316 699556 37372 699558
rect 72836 699610 72892 699612
rect 72916 699610 72972 699612
rect 72996 699610 73052 699612
rect 73076 699610 73132 699612
rect 73156 699610 73212 699612
rect 73236 699610 73292 699612
rect 73316 699610 73372 699612
rect 72836 699558 72874 699610
rect 72874 699558 72886 699610
rect 72886 699558 72892 699610
rect 72916 699558 72938 699610
rect 72938 699558 72950 699610
rect 72950 699558 72972 699610
rect 72996 699558 73002 699610
rect 73002 699558 73014 699610
rect 73014 699558 73052 699610
rect 73076 699558 73078 699610
rect 73078 699558 73130 699610
rect 73130 699558 73132 699610
rect 73156 699558 73194 699610
rect 73194 699558 73206 699610
rect 73206 699558 73212 699610
rect 73236 699558 73258 699610
rect 73258 699558 73270 699610
rect 73270 699558 73292 699610
rect 73316 699558 73322 699610
rect 73322 699558 73334 699610
rect 73334 699558 73372 699610
rect 72836 699556 72892 699558
rect 72916 699556 72972 699558
rect 72996 699556 73052 699558
rect 73076 699556 73132 699558
rect 73156 699556 73212 699558
rect 73236 699556 73292 699558
rect 73316 699556 73372 699558
rect 108836 699610 108892 699612
rect 108916 699610 108972 699612
rect 108996 699610 109052 699612
rect 109076 699610 109132 699612
rect 109156 699610 109212 699612
rect 109236 699610 109292 699612
rect 109316 699610 109372 699612
rect 108836 699558 108874 699610
rect 108874 699558 108886 699610
rect 108886 699558 108892 699610
rect 108916 699558 108938 699610
rect 108938 699558 108950 699610
rect 108950 699558 108972 699610
rect 108996 699558 109002 699610
rect 109002 699558 109014 699610
rect 109014 699558 109052 699610
rect 109076 699558 109078 699610
rect 109078 699558 109130 699610
rect 109130 699558 109132 699610
rect 109156 699558 109194 699610
rect 109194 699558 109206 699610
rect 109206 699558 109212 699610
rect 109236 699558 109258 699610
rect 109258 699558 109270 699610
rect 109270 699558 109292 699610
rect 109316 699558 109322 699610
rect 109322 699558 109334 699610
rect 109334 699558 109372 699610
rect 108836 699556 108892 699558
rect 108916 699556 108972 699558
rect 108996 699556 109052 699558
rect 109076 699556 109132 699558
rect 109156 699556 109212 699558
rect 109236 699556 109292 699558
rect 109316 699556 109372 699558
rect 144836 699610 144892 699612
rect 144916 699610 144972 699612
rect 144996 699610 145052 699612
rect 145076 699610 145132 699612
rect 145156 699610 145212 699612
rect 145236 699610 145292 699612
rect 145316 699610 145372 699612
rect 144836 699558 144874 699610
rect 144874 699558 144886 699610
rect 144886 699558 144892 699610
rect 144916 699558 144938 699610
rect 144938 699558 144950 699610
rect 144950 699558 144972 699610
rect 144996 699558 145002 699610
rect 145002 699558 145014 699610
rect 145014 699558 145052 699610
rect 145076 699558 145078 699610
rect 145078 699558 145130 699610
rect 145130 699558 145132 699610
rect 145156 699558 145194 699610
rect 145194 699558 145206 699610
rect 145206 699558 145212 699610
rect 145236 699558 145258 699610
rect 145258 699558 145270 699610
rect 145270 699558 145292 699610
rect 145316 699558 145322 699610
rect 145322 699558 145334 699610
rect 145334 699558 145372 699610
rect 144836 699556 144892 699558
rect 144916 699556 144972 699558
rect 144996 699556 145052 699558
rect 145076 699556 145132 699558
rect 145156 699556 145212 699558
rect 145236 699556 145292 699558
rect 145316 699556 145372 699558
rect 4802 699216 4858 699272
rect 2870 682216 2926 682272
rect 2778 667936 2834 667992
rect 3054 653556 3056 653576
rect 3056 653556 3108 653576
rect 3108 653556 3110 653576
rect 3054 653520 3110 653556
rect 2962 624860 2964 624880
rect 2964 624860 3016 624880
rect 3016 624860 3018 624880
rect 2962 624824 3018 624860
rect 2778 610408 2834 610464
rect 3054 596028 3056 596048
rect 3056 596028 3108 596048
rect 3108 596028 3110 596048
rect 3054 595992 3110 596028
rect 2962 567296 3018 567352
rect 3146 553016 3202 553072
rect 3238 538600 3294 538656
rect 3054 509904 3110 509960
rect 3238 481108 3240 481128
rect 3240 481108 3292 481128
rect 3292 481108 3294 481128
rect 3238 481072 3294 481108
rect 3054 452412 3056 452432
rect 3056 452412 3108 452432
rect 3108 452412 3110 452432
rect 3054 452376 3110 452412
rect 3422 695680 3478 695736
rect 3330 437960 3386 438016
rect 3330 423680 3386 423736
rect 3330 394984 3386 395040
rect 3330 366188 3332 366208
rect 3332 366188 3384 366208
rect 3384 366188 3386 366208
rect 3330 366152 3386 366188
rect 3330 337456 3386 337512
rect 2778 323040 2834 323096
rect 3330 294344 3386 294400
rect 2778 280084 2834 280120
rect 2778 280064 2780 280084
rect 2780 280064 2832 280084
rect 2832 280064 2834 280084
rect 3146 265648 3202 265704
rect 3238 251232 3294 251288
rect 3146 208156 3148 208176
rect 3148 208156 3200 208176
rect 3200 208156 3202 208176
rect 3146 208120 3202 208156
rect 2778 193840 2834 193896
rect 1122 165008 1178 165064
rect 2778 150728 2834 150784
rect 3330 136348 3332 136368
rect 3332 136348 3384 136368
rect 3384 136348 3386 136368
rect 3330 136312 3386 136348
rect 3330 122068 3332 122088
rect 3332 122068 3384 122088
rect 3384 122068 3386 122088
rect 3330 122032 3386 122068
rect 3054 78920 3110 78976
rect 2778 64540 2780 64560
rect 2780 64540 2832 64560
rect 2832 64540 2834 64560
rect 2778 64504 2834 64540
rect 3514 693912 3570 693968
rect 3974 495488 4030 495544
rect 3882 308760 3938 308816
rect 3790 222536 3846 222592
rect 3698 179424 3754 179480
rect 4066 380568 4122 380624
rect 4066 236952 4122 237008
rect 3974 107616 4030 107672
rect 3606 93200 3662 93256
rect 18836 699066 18892 699068
rect 18916 699066 18972 699068
rect 18996 699066 19052 699068
rect 19076 699066 19132 699068
rect 19156 699066 19212 699068
rect 19236 699066 19292 699068
rect 19316 699066 19372 699068
rect 18836 699014 18874 699066
rect 18874 699014 18886 699066
rect 18886 699014 18892 699066
rect 18916 699014 18938 699066
rect 18938 699014 18950 699066
rect 18950 699014 18972 699066
rect 18996 699014 19002 699066
rect 19002 699014 19014 699066
rect 19014 699014 19052 699066
rect 19076 699014 19078 699066
rect 19078 699014 19130 699066
rect 19130 699014 19132 699066
rect 19156 699014 19194 699066
rect 19194 699014 19206 699066
rect 19206 699014 19212 699066
rect 19236 699014 19258 699066
rect 19258 699014 19270 699066
rect 19270 699014 19292 699066
rect 19316 699014 19322 699066
rect 19322 699014 19334 699066
rect 19334 699014 19372 699066
rect 18836 699012 18892 699014
rect 18916 699012 18972 699014
rect 18996 699012 19052 699014
rect 19076 699012 19132 699014
rect 19156 699012 19212 699014
rect 19236 699012 19292 699014
rect 19316 699012 19372 699014
rect 54836 699066 54892 699068
rect 54916 699066 54972 699068
rect 54996 699066 55052 699068
rect 55076 699066 55132 699068
rect 55156 699066 55212 699068
rect 55236 699066 55292 699068
rect 55316 699066 55372 699068
rect 54836 699014 54874 699066
rect 54874 699014 54886 699066
rect 54886 699014 54892 699066
rect 54916 699014 54938 699066
rect 54938 699014 54950 699066
rect 54950 699014 54972 699066
rect 54996 699014 55002 699066
rect 55002 699014 55014 699066
rect 55014 699014 55052 699066
rect 55076 699014 55078 699066
rect 55078 699014 55130 699066
rect 55130 699014 55132 699066
rect 55156 699014 55194 699066
rect 55194 699014 55206 699066
rect 55206 699014 55212 699066
rect 55236 699014 55258 699066
rect 55258 699014 55270 699066
rect 55270 699014 55292 699066
rect 55316 699014 55322 699066
rect 55322 699014 55334 699066
rect 55334 699014 55372 699066
rect 54836 699012 54892 699014
rect 54916 699012 54972 699014
rect 54996 699012 55052 699014
rect 55076 699012 55132 699014
rect 55156 699012 55212 699014
rect 55236 699012 55292 699014
rect 55316 699012 55372 699014
rect 43442 698808 43498 698864
rect 5354 698672 5410 698728
rect 29182 698264 29238 698320
rect 6182 697040 6238 697096
rect 3514 50088 3570 50144
rect 3514 35828 3570 35864
rect 3514 35808 3516 35828
rect 3516 35808 3568 35828
rect 3568 35808 3570 35828
rect 3422 21392 3478 21448
rect 7654 693640 7710 693696
rect 10322 696904 10378 696960
rect 36836 698522 36892 698524
rect 36916 698522 36972 698524
rect 36996 698522 37052 698524
rect 37076 698522 37132 698524
rect 37156 698522 37212 698524
rect 37236 698522 37292 698524
rect 37316 698522 37372 698524
rect 36836 698470 36874 698522
rect 36874 698470 36886 698522
rect 36886 698470 36892 698522
rect 36916 698470 36938 698522
rect 36938 698470 36950 698522
rect 36950 698470 36972 698522
rect 36996 698470 37002 698522
rect 37002 698470 37014 698522
rect 37014 698470 37052 698522
rect 37076 698470 37078 698522
rect 37078 698470 37130 698522
rect 37130 698470 37132 698522
rect 37156 698470 37194 698522
rect 37194 698470 37206 698522
rect 37206 698470 37212 698522
rect 37236 698470 37258 698522
rect 37258 698470 37270 698522
rect 37270 698470 37292 698522
rect 37316 698470 37322 698522
rect 37322 698470 37334 698522
rect 37334 698470 37372 698522
rect 36836 698468 36892 698470
rect 36916 698468 36972 698470
rect 36996 698468 37052 698470
rect 37076 698468 37132 698470
rect 37156 698468 37212 698470
rect 37236 698468 37292 698470
rect 37316 698468 37372 698470
rect 72836 698522 72892 698524
rect 72916 698522 72972 698524
rect 72996 698522 73052 698524
rect 73076 698522 73132 698524
rect 73156 698522 73212 698524
rect 73236 698522 73292 698524
rect 73316 698522 73372 698524
rect 72836 698470 72874 698522
rect 72874 698470 72886 698522
rect 72886 698470 72892 698522
rect 72916 698470 72938 698522
rect 72938 698470 72950 698522
rect 72950 698470 72972 698522
rect 72996 698470 73002 698522
rect 73002 698470 73014 698522
rect 73014 698470 73052 698522
rect 73076 698470 73078 698522
rect 73078 698470 73130 698522
rect 73130 698470 73132 698522
rect 73156 698470 73194 698522
rect 73194 698470 73206 698522
rect 73206 698470 73212 698522
rect 73236 698470 73258 698522
rect 73258 698470 73270 698522
rect 73270 698470 73292 698522
rect 73316 698470 73322 698522
rect 73322 698470 73334 698522
rect 73334 698470 73372 698522
rect 72836 698468 72892 698470
rect 72916 698468 72972 698470
rect 72996 698468 73052 698470
rect 73076 698468 73132 698470
rect 73156 698468 73212 698470
rect 73236 698468 73292 698470
rect 73316 698468 73372 698470
rect 90836 699066 90892 699068
rect 90916 699066 90972 699068
rect 90996 699066 91052 699068
rect 91076 699066 91132 699068
rect 91156 699066 91212 699068
rect 91236 699066 91292 699068
rect 91316 699066 91372 699068
rect 90836 699014 90874 699066
rect 90874 699014 90886 699066
rect 90886 699014 90892 699066
rect 90916 699014 90938 699066
rect 90938 699014 90950 699066
rect 90950 699014 90972 699066
rect 90996 699014 91002 699066
rect 91002 699014 91014 699066
rect 91014 699014 91052 699066
rect 91076 699014 91078 699066
rect 91078 699014 91130 699066
rect 91130 699014 91132 699066
rect 91156 699014 91194 699066
rect 91194 699014 91206 699066
rect 91206 699014 91212 699066
rect 91236 699014 91258 699066
rect 91258 699014 91270 699066
rect 91270 699014 91292 699066
rect 91316 699014 91322 699066
rect 91322 699014 91334 699066
rect 91334 699014 91372 699066
rect 90836 699012 90892 699014
rect 90916 699012 90972 699014
rect 90996 699012 91052 699014
rect 91076 699012 91132 699014
rect 91156 699012 91212 699014
rect 91236 699012 91292 699014
rect 91316 699012 91372 699014
rect 108836 698522 108892 698524
rect 108916 698522 108972 698524
rect 108996 698522 109052 698524
rect 109076 698522 109132 698524
rect 109156 698522 109212 698524
rect 109236 698522 109292 698524
rect 109316 698522 109372 698524
rect 108836 698470 108874 698522
rect 108874 698470 108886 698522
rect 108886 698470 108892 698522
rect 108916 698470 108938 698522
rect 108938 698470 108950 698522
rect 108950 698470 108972 698522
rect 108996 698470 109002 698522
rect 109002 698470 109014 698522
rect 109014 698470 109052 698522
rect 109076 698470 109078 698522
rect 109078 698470 109130 698522
rect 109130 698470 109132 698522
rect 109156 698470 109194 698522
rect 109194 698470 109206 698522
rect 109206 698470 109212 698522
rect 109236 698470 109258 698522
rect 109258 698470 109270 698522
rect 109270 698470 109292 698522
rect 109316 698470 109322 698522
rect 109322 698470 109334 698522
rect 109334 698470 109372 698522
rect 108836 698468 108892 698470
rect 108916 698468 108972 698470
rect 108996 698468 109052 698470
rect 109076 698468 109132 698470
rect 109156 698468 109212 698470
rect 109236 698468 109292 698470
rect 109316 698468 109372 698470
rect 126836 699066 126892 699068
rect 126916 699066 126972 699068
rect 126996 699066 127052 699068
rect 127076 699066 127132 699068
rect 127156 699066 127212 699068
rect 127236 699066 127292 699068
rect 127316 699066 127372 699068
rect 126836 699014 126874 699066
rect 126874 699014 126886 699066
rect 126886 699014 126892 699066
rect 126916 699014 126938 699066
rect 126938 699014 126950 699066
rect 126950 699014 126972 699066
rect 126996 699014 127002 699066
rect 127002 699014 127014 699066
rect 127014 699014 127052 699066
rect 127076 699014 127078 699066
rect 127078 699014 127130 699066
rect 127130 699014 127132 699066
rect 127156 699014 127194 699066
rect 127194 699014 127206 699066
rect 127206 699014 127212 699066
rect 127236 699014 127258 699066
rect 127258 699014 127270 699066
rect 127270 699014 127292 699066
rect 127316 699014 127322 699066
rect 127322 699014 127334 699066
rect 127334 699014 127372 699066
rect 126836 699012 126892 699014
rect 126916 699012 126972 699014
rect 126996 699012 127052 699014
rect 127076 699012 127132 699014
rect 127156 699012 127212 699014
rect 127236 699012 127292 699014
rect 127316 699012 127372 699014
rect 144836 698522 144892 698524
rect 144916 698522 144972 698524
rect 144996 698522 145052 698524
rect 145076 698522 145132 698524
rect 145156 698522 145212 698524
rect 145236 698522 145292 698524
rect 145316 698522 145372 698524
rect 144836 698470 144874 698522
rect 144874 698470 144886 698522
rect 144886 698470 144892 698522
rect 144916 698470 144938 698522
rect 144938 698470 144950 698522
rect 144950 698470 144972 698522
rect 144996 698470 145002 698522
rect 145002 698470 145014 698522
rect 145014 698470 145052 698522
rect 145076 698470 145078 698522
rect 145078 698470 145130 698522
rect 145130 698470 145132 698522
rect 145156 698470 145194 698522
rect 145194 698470 145206 698522
rect 145206 698470 145212 698522
rect 145236 698470 145258 698522
rect 145258 698470 145270 698522
rect 145270 698470 145292 698522
rect 145316 698470 145322 698522
rect 145322 698470 145334 698522
rect 145334 698470 145372 698522
rect 144836 698468 144892 698470
rect 144916 698468 144972 698470
rect 144996 698468 145052 698470
rect 145076 698468 145132 698470
rect 145156 698468 145212 698470
rect 145236 698468 145292 698470
rect 145316 698468 145372 698470
rect 162836 699066 162892 699068
rect 162916 699066 162972 699068
rect 162996 699066 163052 699068
rect 163076 699066 163132 699068
rect 163156 699066 163212 699068
rect 163236 699066 163292 699068
rect 163316 699066 163372 699068
rect 162836 699014 162874 699066
rect 162874 699014 162886 699066
rect 162886 699014 162892 699066
rect 162916 699014 162938 699066
rect 162938 699014 162950 699066
rect 162950 699014 162972 699066
rect 162996 699014 163002 699066
rect 163002 699014 163014 699066
rect 163014 699014 163052 699066
rect 163076 699014 163078 699066
rect 163078 699014 163130 699066
rect 163130 699014 163132 699066
rect 163156 699014 163194 699066
rect 163194 699014 163206 699066
rect 163206 699014 163212 699066
rect 163236 699014 163258 699066
rect 163258 699014 163270 699066
rect 163270 699014 163292 699066
rect 163316 699014 163322 699066
rect 163322 699014 163334 699066
rect 163334 699014 163372 699066
rect 162836 699012 162892 699014
rect 162916 699012 162972 699014
rect 162996 699012 163052 699014
rect 163076 699012 163132 699014
rect 163156 699012 163212 699014
rect 163236 699012 163292 699014
rect 163316 699012 163372 699014
rect 173898 695988 173900 696008
rect 173900 695988 173952 696008
rect 173952 695988 173954 696008
rect 173898 695952 173954 695988
rect 174266 695988 174268 696008
rect 174268 695988 174320 696008
rect 174320 695988 174322 696008
rect 174266 695952 174322 695988
rect 19982 695544 20038 695600
rect 15290 695272 15346 695328
rect 176198 695272 176254 695328
rect 180836 699610 180892 699612
rect 180916 699610 180972 699612
rect 180996 699610 181052 699612
rect 181076 699610 181132 699612
rect 181156 699610 181212 699612
rect 181236 699610 181292 699612
rect 181316 699610 181372 699612
rect 180836 699558 180874 699610
rect 180874 699558 180886 699610
rect 180886 699558 180892 699610
rect 180916 699558 180938 699610
rect 180938 699558 180950 699610
rect 180950 699558 180972 699610
rect 180996 699558 181002 699610
rect 181002 699558 181014 699610
rect 181014 699558 181052 699610
rect 181076 699558 181078 699610
rect 181078 699558 181130 699610
rect 181130 699558 181132 699610
rect 181156 699558 181194 699610
rect 181194 699558 181206 699610
rect 181206 699558 181212 699610
rect 181236 699558 181258 699610
rect 181258 699558 181270 699610
rect 181270 699558 181292 699610
rect 181316 699558 181322 699610
rect 181322 699558 181334 699610
rect 181334 699558 181372 699610
rect 180836 699556 180892 699558
rect 180916 699556 180972 699558
rect 180996 699556 181052 699558
rect 181076 699556 181132 699558
rect 181156 699556 181212 699558
rect 181236 699556 181292 699558
rect 181316 699556 181372 699558
rect 216836 699610 216892 699612
rect 216916 699610 216972 699612
rect 216996 699610 217052 699612
rect 217076 699610 217132 699612
rect 217156 699610 217212 699612
rect 217236 699610 217292 699612
rect 217316 699610 217372 699612
rect 216836 699558 216874 699610
rect 216874 699558 216886 699610
rect 216886 699558 216892 699610
rect 216916 699558 216938 699610
rect 216938 699558 216950 699610
rect 216950 699558 216972 699610
rect 216996 699558 217002 699610
rect 217002 699558 217014 699610
rect 217014 699558 217052 699610
rect 217076 699558 217078 699610
rect 217078 699558 217130 699610
rect 217130 699558 217132 699610
rect 217156 699558 217194 699610
rect 217194 699558 217206 699610
rect 217206 699558 217212 699610
rect 217236 699558 217258 699610
rect 217258 699558 217270 699610
rect 217270 699558 217292 699610
rect 217316 699558 217322 699610
rect 217322 699558 217334 699610
rect 217334 699558 217372 699610
rect 216836 699556 216892 699558
rect 216916 699556 216972 699558
rect 216996 699556 217052 699558
rect 217076 699556 217132 699558
rect 217156 699556 217212 699558
rect 217236 699556 217292 699558
rect 217316 699556 217372 699558
rect 190458 699352 190514 699408
rect 200026 699352 200082 699408
rect 180798 699116 180800 699136
rect 180800 699116 180852 699136
rect 180852 699116 180854 699136
rect 180798 699080 180854 699116
rect 190366 699116 190368 699136
rect 190368 699116 190420 699136
rect 190420 699116 190422 699136
rect 190366 699080 190422 699116
rect 209778 699116 209780 699136
rect 209780 699116 209832 699136
rect 209832 699116 209834 699136
rect 209778 699080 209834 699116
rect 219346 699116 219348 699136
rect 219348 699116 219400 699136
rect 219400 699116 219402 699136
rect 219346 699080 219402 699116
rect 198836 699066 198892 699068
rect 198916 699066 198972 699068
rect 198996 699066 199052 699068
rect 199076 699066 199132 699068
rect 199156 699066 199212 699068
rect 199236 699066 199292 699068
rect 199316 699066 199372 699068
rect 198836 699014 198874 699066
rect 198874 699014 198886 699066
rect 198886 699014 198892 699066
rect 198916 699014 198938 699066
rect 198938 699014 198950 699066
rect 198950 699014 198972 699066
rect 198996 699014 199002 699066
rect 199002 699014 199014 699066
rect 199014 699014 199052 699066
rect 199076 699014 199078 699066
rect 199078 699014 199130 699066
rect 199130 699014 199132 699066
rect 199156 699014 199194 699066
rect 199194 699014 199206 699066
rect 199206 699014 199212 699066
rect 199236 699014 199258 699066
rect 199258 699014 199270 699066
rect 199270 699014 199292 699066
rect 199316 699014 199322 699066
rect 199322 699014 199334 699066
rect 199334 699014 199372 699066
rect 198836 699012 198892 699014
rect 198916 699012 198972 699014
rect 198996 699012 199052 699014
rect 199076 699012 199132 699014
rect 199156 699012 199212 699014
rect 199236 699012 199292 699014
rect 199316 699012 199372 699014
rect 180836 698522 180892 698524
rect 180916 698522 180972 698524
rect 180996 698522 181052 698524
rect 181076 698522 181132 698524
rect 181156 698522 181212 698524
rect 181236 698522 181292 698524
rect 181316 698522 181372 698524
rect 180836 698470 180874 698522
rect 180874 698470 180886 698522
rect 180886 698470 180892 698522
rect 180916 698470 180938 698522
rect 180938 698470 180950 698522
rect 180950 698470 180972 698522
rect 180996 698470 181002 698522
rect 181002 698470 181014 698522
rect 181014 698470 181052 698522
rect 181076 698470 181078 698522
rect 181078 698470 181130 698522
rect 181130 698470 181132 698522
rect 181156 698470 181194 698522
rect 181194 698470 181206 698522
rect 181206 698470 181212 698522
rect 181236 698470 181258 698522
rect 181258 698470 181270 698522
rect 181270 698470 181292 698522
rect 181316 698470 181322 698522
rect 181322 698470 181334 698522
rect 181334 698470 181372 698522
rect 180836 698468 180892 698470
rect 180916 698468 180972 698470
rect 180996 698468 181052 698470
rect 181076 698468 181132 698470
rect 181156 698468 181212 698470
rect 181236 698468 181292 698470
rect 181316 698468 181372 698470
rect 216836 698522 216892 698524
rect 216916 698522 216972 698524
rect 216996 698522 217052 698524
rect 217076 698522 217132 698524
rect 217156 698522 217212 698524
rect 217236 698522 217292 698524
rect 217316 698522 217372 698524
rect 216836 698470 216874 698522
rect 216874 698470 216886 698522
rect 216886 698470 216892 698522
rect 216916 698470 216938 698522
rect 216938 698470 216950 698522
rect 216950 698470 216972 698522
rect 216996 698470 217002 698522
rect 217002 698470 217014 698522
rect 217014 698470 217052 698522
rect 217076 698470 217078 698522
rect 217078 698470 217130 698522
rect 217130 698470 217132 698522
rect 217156 698470 217194 698522
rect 217194 698470 217206 698522
rect 217206 698470 217212 698522
rect 217236 698470 217258 698522
rect 217258 698470 217270 698522
rect 217270 698470 217292 698522
rect 217316 698470 217322 698522
rect 217322 698470 217334 698522
rect 217334 698470 217372 698522
rect 216836 698468 216892 698470
rect 216916 698468 216972 698470
rect 216996 698468 217052 698470
rect 217076 698468 217132 698470
rect 217156 698468 217212 698470
rect 217236 698468 217292 698470
rect 217316 698468 217372 698470
rect 234836 701242 234892 701244
rect 234916 701242 234972 701244
rect 234996 701242 235052 701244
rect 235076 701242 235132 701244
rect 235156 701242 235212 701244
rect 235236 701242 235292 701244
rect 235316 701242 235372 701244
rect 234836 701190 234874 701242
rect 234874 701190 234886 701242
rect 234886 701190 234892 701242
rect 234916 701190 234938 701242
rect 234938 701190 234950 701242
rect 234950 701190 234972 701242
rect 234996 701190 235002 701242
rect 235002 701190 235014 701242
rect 235014 701190 235052 701242
rect 235076 701190 235078 701242
rect 235078 701190 235130 701242
rect 235130 701190 235132 701242
rect 235156 701190 235194 701242
rect 235194 701190 235206 701242
rect 235206 701190 235212 701242
rect 235236 701190 235258 701242
rect 235258 701190 235270 701242
rect 235270 701190 235292 701242
rect 235316 701190 235322 701242
rect 235322 701190 235334 701242
rect 235334 701190 235372 701242
rect 234836 701188 234892 701190
rect 234916 701188 234972 701190
rect 234996 701188 235052 701190
rect 235076 701188 235132 701190
rect 235156 701188 235212 701190
rect 235236 701188 235292 701190
rect 235316 701188 235372 701190
rect 227994 700848 228050 700904
rect 234836 700154 234892 700156
rect 234916 700154 234972 700156
rect 234996 700154 235052 700156
rect 235076 700154 235132 700156
rect 235156 700154 235212 700156
rect 235236 700154 235292 700156
rect 235316 700154 235372 700156
rect 234836 700102 234874 700154
rect 234874 700102 234886 700154
rect 234886 700102 234892 700154
rect 234916 700102 234938 700154
rect 234938 700102 234950 700154
rect 234950 700102 234972 700154
rect 234996 700102 235002 700154
rect 235002 700102 235014 700154
rect 235014 700102 235052 700154
rect 235076 700102 235078 700154
rect 235078 700102 235130 700154
rect 235130 700102 235132 700154
rect 235156 700102 235194 700154
rect 235194 700102 235206 700154
rect 235206 700102 235212 700154
rect 235236 700102 235258 700154
rect 235258 700102 235270 700154
rect 235270 700102 235292 700154
rect 235316 700102 235322 700154
rect 235322 700102 235334 700154
rect 235334 700102 235372 700154
rect 234836 700100 234892 700102
rect 234916 700100 234972 700102
rect 234996 700100 235052 700102
rect 235076 700100 235132 700102
rect 235156 700100 235212 700102
rect 235236 700100 235292 700102
rect 235316 700100 235372 700102
rect 229098 699352 229154 699408
rect 234836 699066 234892 699068
rect 234916 699066 234972 699068
rect 234996 699066 235052 699068
rect 235076 699066 235132 699068
rect 235156 699066 235212 699068
rect 235236 699066 235292 699068
rect 235316 699066 235372 699068
rect 234836 699014 234874 699066
rect 234874 699014 234886 699066
rect 234886 699014 234892 699066
rect 234916 699014 234938 699066
rect 234938 699014 234950 699066
rect 234950 699014 234972 699066
rect 234996 699014 235002 699066
rect 235002 699014 235014 699066
rect 235014 699014 235052 699066
rect 235076 699014 235078 699066
rect 235078 699014 235130 699066
rect 235130 699014 235132 699066
rect 235156 699014 235194 699066
rect 235194 699014 235206 699066
rect 235206 699014 235212 699066
rect 235236 699014 235258 699066
rect 235258 699014 235270 699066
rect 235270 699014 235292 699066
rect 235316 699014 235322 699066
rect 235322 699014 235334 699066
rect 235334 699014 235372 699066
rect 234836 699012 234892 699014
rect 234916 699012 234972 699014
rect 234996 699012 235052 699014
rect 235076 699012 235132 699014
rect 235156 699012 235212 699014
rect 235236 699012 235292 699014
rect 235316 699012 235372 699014
rect 233054 698808 233110 698864
rect 234710 698808 234766 698864
rect 241518 699624 241574 699680
rect 244186 700032 244242 700088
rect 244186 699352 244242 699408
rect 244094 698944 244150 699000
rect 251086 700032 251142 700088
rect 251086 699624 251142 699680
rect 252836 701786 252892 701788
rect 252916 701786 252972 701788
rect 252996 701786 253052 701788
rect 253076 701786 253132 701788
rect 253156 701786 253212 701788
rect 253236 701786 253292 701788
rect 253316 701786 253372 701788
rect 252836 701734 252874 701786
rect 252874 701734 252886 701786
rect 252886 701734 252892 701786
rect 252916 701734 252938 701786
rect 252938 701734 252950 701786
rect 252950 701734 252972 701786
rect 252996 701734 253002 701786
rect 253002 701734 253014 701786
rect 253014 701734 253052 701786
rect 253076 701734 253078 701786
rect 253078 701734 253130 701786
rect 253130 701734 253132 701786
rect 253156 701734 253194 701786
rect 253194 701734 253206 701786
rect 253206 701734 253212 701786
rect 253236 701734 253258 701786
rect 253258 701734 253270 701786
rect 253270 701734 253292 701786
rect 253316 701734 253322 701786
rect 253322 701734 253334 701786
rect 253334 701734 253372 701786
rect 252836 701732 252892 701734
rect 252916 701732 252972 701734
rect 252996 701732 253052 701734
rect 253076 701732 253132 701734
rect 253156 701732 253212 701734
rect 253236 701732 253292 701734
rect 253316 701732 253372 701734
rect 252836 700698 252892 700700
rect 252916 700698 252972 700700
rect 252996 700698 253052 700700
rect 253076 700698 253132 700700
rect 253156 700698 253212 700700
rect 253236 700698 253292 700700
rect 253316 700698 253372 700700
rect 252836 700646 252874 700698
rect 252874 700646 252886 700698
rect 252886 700646 252892 700698
rect 252916 700646 252938 700698
rect 252938 700646 252950 700698
rect 252950 700646 252972 700698
rect 252996 700646 253002 700698
rect 253002 700646 253014 700698
rect 253014 700646 253052 700698
rect 253076 700646 253078 700698
rect 253078 700646 253130 700698
rect 253130 700646 253132 700698
rect 253156 700646 253194 700698
rect 253194 700646 253206 700698
rect 253206 700646 253212 700698
rect 253236 700646 253258 700698
rect 253258 700646 253270 700698
rect 253270 700646 253292 700698
rect 253316 700646 253322 700698
rect 253322 700646 253334 700698
rect 253334 700646 253372 700698
rect 252836 700644 252892 700646
rect 252916 700644 252972 700646
rect 252996 700644 253052 700646
rect 253076 700644 253132 700646
rect 253156 700644 253212 700646
rect 253236 700644 253292 700646
rect 253316 700644 253372 700646
rect 252836 699610 252892 699612
rect 252916 699610 252972 699612
rect 252996 699610 253052 699612
rect 253076 699610 253132 699612
rect 253156 699610 253212 699612
rect 253236 699610 253292 699612
rect 253316 699610 253372 699612
rect 252836 699558 252874 699610
rect 252874 699558 252886 699610
rect 252886 699558 252892 699610
rect 252916 699558 252938 699610
rect 252938 699558 252950 699610
rect 252950 699558 252972 699610
rect 252996 699558 253002 699610
rect 253002 699558 253014 699610
rect 253014 699558 253052 699610
rect 253076 699558 253078 699610
rect 253078 699558 253130 699610
rect 253130 699558 253132 699610
rect 253156 699558 253194 699610
rect 253194 699558 253206 699610
rect 253206 699558 253212 699610
rect 253236 699558 253258 699610
rect 253258 699558 253270 699610
rect 253270 699558 253292 699610
rect 253316 699558 253322 699610
rect 253322 699558 253334 699610
rect 253334 699558 253372 699610
rect 252836 699556 252892 699558
rect 252916 699556 252972 699558
rect 252996 699556 253052 699558
rect 253076 699556 253132 699558
rect 253156 699556 253212 699558
rect 253236 699556 253292 699558
rect 253316 699556 253372 699558
rect 253662 699116 253664 699136
rect 253664 699116 253716 699136
rect 253716 699116 253718 699136
rect 253662 699080 253718 699116
rect 253846 698944 253902 699000
rect 253754 698844 253756 698864
rect 253756 698844 253808 698864
rect 253808 698844 253810 698864
rect 253754 698808 253810 698844
rect 252836 698522 252892 698524
rect 252916 698522 252972 698524
rect 252996 698522 253052 698524
rect 253076 698522 253132 698524
rect 253156 698522 253212 698524
rect 253236 698522 253292 698524
rect 253316 698522 253372 698524
rect 252836 698470 252874 698522
rect 252874 698470 252886 698522
rect 252886 698470 252892 698522
rect 252916 698470 252938 698522
rect 252938 698470 252950 698522
rect 252950 698470 252972 698522
rect 252996 698470 253002 698522
rect 253002 698470 253014 698522
rect 253014 698470 253052 698522
rect 253076 698470 253078 698522
rect 253078 698470 253130 698522
rect 253130 698470 253132 698522
rect 253156 698470 253194 698522
rect 253194 698470 253206 698522
rect 253206 698470 253212 698522
rect 253236 698470 253258 698522
rect 253258 698470 253270 698522
rect 253270 698470 253292 698522
rect 253316 698470 253322 698522
rect 253322 698470 253334 698522
rect 253334 698470 253372 698522
rect 252836 698468 252892 698470
rect 252916 698468 252972 698470
rect 252996 698468 253052 698470
rect 253076 698468 253132 698470
rect 253156 698468 253212 698470
rect 253236 698468 253292 698470
rect 253316 698468 253372 698470
rect 270836 701242 270892 701244
rect 270916 701242 270972 701244
rect 270996 701242 271052 701244
rect 271076 701242 271132 701244
rect 271156 701242 271212 701244
rect 271236 701242 271292 701244
rect 271316 701242 271372 701244
rect 270836 701190 270874 701242
rect 270874 701190 270886 701242
rect 270886 701190 270892 701242
rect 270916 701190 270938 701242
rect 270938 701190 270950 701242
rect 270950 701190 270972 701242
rect 270996 701190 271002 701242
rect 271002 701190 271014 701242
rect 271014 701190 271052 701242
rect 271076 701190 271078 701242
rect 271078 701190 271130 701242
rect 271130 701190 271132 701242
rect 271156 701190 271194 701242
rect 271194 701190 271206 701242
rect 271206 701190 271212 701242
rect 271236 701190 271258 701242
rect 271258 701190 271270 701242
rect 271270 701190 271292 701242
rect 271316 701190 271322 701242
rect 271322 701190 271334 701242
rect 271334 701190 271372 701242
rect 270836 701188 270892 701190
rect 270916 701188 270972 701190
rect 270996 701188 271052 701190
rect 271076 701188 271132 701190
rect 271156 701188 271212 701190
rect 271236 701188 271292 701190
rect 271316 701188 271372 701190
rect 270836 700154 270892 700156
rect 270916 700154 270972 700156
rect 270996 700154 271052 700156
rect 271076 700154 271132 700156
rect 271156 700154 271212 700156
rect 271236 700154 271292 700156
rect 271316 700154 271372 700156
rect 270836 700102 270874 700154
rect 270874 700102 270886 700154
rect 270886 700102 270892 700154
rect 270916 700102 270938 700154
rect 270938 700102 270950 700154
rect 270950 700102 270972 700154
rect 270996 700102 271002 700154
rect 271002 700102 271014 700154
rect 271014 700102 271052 700154
rect 271076 700102 271078 700154
rect 271078 700102 271130 700154
rect 271130 700102 271132 700154
rect 271156 700102 271194 700154
rect 271194 700102 271206 700154
rect 271206 700102 271212 700154
rect 271236 700102 271258 700154
rect 271258 700102 271270 700154
rect 271270 700102 271292 700154
rect 271316 700102 271322 700154
rect 271322 700102 271334 700154
rect 271334 700102 271372 700154
rect 270836 700100 270892 700102
rect 270916 700100 270972 700102
rect 270996 700100 271052 700102
rect 271076 700100 271132 700102
rect 271156 700100 271212 700102
rect 271236 700100 271292 700102
rect 271316 700100 271372 700102
rect 280066 700032 280122 700088
rect 288836 701786 288892 701788
rect 288916 701786 288972 701788
rect 288996 701786 289052 701788
rect 289076 701786 289132 701788
rect 289156 701786 289212 701788
rect 289236 701786 289292 701788
rect 289316 701786 289372 701788
rect 288836 701734 288874 701786
rect 288874 701734 288886 701786
rect 288886 701734 288892 701786
rect 288916 701734 288938 701786
rect 288938 701734 288950 701786
rect 288950 701734 288972 701786
rect 288996 701734 289002 701786
rect 289002 701734 289014 701786
rect 289014 701734 289052 701786
rect 289076 701734 289078 701786
rect 289078 701734 289130 701786
rect 289130 701734 289132 701786
rect 289156 701734 289194 701786
rect 289194 701734 289206 701786
rect 289206 701734 289212 701786
rect 289236 701734 289258 701786
rect 289258 701734 289270 701786
rect 289270 701734 289292 701786
rect 289316 701734 289322 701786
rect 289322 701734 289334 701786
rect 289334 701734 289372 701786
rect 288836 701732 288892 701734
rect 288916 701732 288972 701734
rect 288996 701732 289052 701734
rect 289076 701732 289132 701734
rect 289156 701732 289212 701734
rect 289236 701732 289292 701734
rect 289316 701732 289372 701734
rect 288836 700698 288892 700700
rect 288916 700698 288972 700700
rect 288996 700698 289052 700700
rect 289076 700698 289132 700700
rect 289156 700698 289212 700700
rect 289236 700698 289292 700700
rect 289316 700698 289372 700700
rect 288836 700646 288874 700698
rect 288874 700646 288886 700698
rect 288886 700646 288892 700698
rect 288916 700646 288938 700698
rect 288938 700646 288950 700698
rect 288950 700646 288972 700698
rect 288996 700646 289002 700698
rect 289002 700646 289014 700698
rect 289014 700646 289052 700698
rect 289076 700646 289078 700698
rect 289078 700646 289130 700698
rect 289130 700646 289132 700698
rect 289156 700646 289194 700698
rect 289194 700646 289206 700698
rect 289206 700646 289212 700698
rect 289236 700646 289258 700698
rect 289258 700646 289270 700698
rect 289270 700646 289292 700698
rect 289316 700646 289322 700698
rect 289322 700646 289334 700698
rect 289334 700646 289372 700698
rect 288836 700644 288892 700646
rect 288916 700644 288972 700646
rect 288996 700644 289052 700646
rect 289076 700644 289132 700646
rect 289156 700644 289212 700646
rect 289236 700644 289292 700646
rect 289316 700644 289372 700646
rect 324836 701786 324892 701788
rect 324916 701786 324972 701788
rect 324996 701786 325052 701788
rect 325076 701786 325132 701788
rect 325156 701786 325212 701788
rect 325236 701786 325292 701788
rect 325316 701786 325372 701788
rect 324836 701734 324874 701786
rect 324874 701734 324886 701786
rect 324886 701734 324892 701786
rect 324916 701734 324938 701786
rect 324938 701734 324950 701786
rect 324950 701734 324972 701786
rect 324996 701734 325002 701786
rect 325002 701734 325014 701786
rect 325014 701734 325052 701786
rect 325076 701734 325078 701786
rect 325078 701734 325130 701786
rect 325130 701734 325132 701786
rect 325156 701734 325194 701786
rect 325194 701734 325206 701786
rect 325206 701734 325212 701786
rect 325236 701734 325258 701786
rect 325258 701734 325270 701786
rect 325270 701734 325292 701786
rect 325316 701734 325322 701786
rect 325322 701734 325334 701786
rect 325334 701734 325372 701786
rect 324836 701732 324892 701734
rect 324916 701732 324972 701734
rect 324996 701732 325052 701734
rect 325076 701732 325132 701734
rect 325156 701732 325212 701734
rect 325236 701732 325292 701734
rect 325316 701732 325372 701734
rect 306836 701242 306892 701244
rect 306916 701242 306972 701244
rect 306996 701242 307052 701244
rect 307076 701242 307132 701244
rect 307156 701242 307212 701244
rect 307236 701242 307292 701244
rect 307316 701242 307372 701244
rect 306836 701190 306874 701242
rect 306874 701190 306886 701242
rect 306886 701190 306892 701242
rect 306916 701190 306938 701242
rect 306938 701190 306950 701242
rect 306950 701190 306972 701242
rect 306996 701190 307002 701242
rect 307002 701190 307014 701242
rect 307014 701190 307052 701242
rect 307076 701190 307078 701242
rect 307078 701190 307130 701242
rect 307130 701190 307132 701242
rect 307156 701190 307194 701242
rect 307194 701190 307206 701242
rect 307206 701190 307212 701242
rect 307236 701190 307258 701242
rect 307258 701190 307270 701242
rect 307270 701190 307292 701242
rect 307316 701190 307322 701242
rect 307322 701190 307334 701242
rect 307334 701190 307372 701242
rect 306836 701188 306892 701190
rect 306916 701188 306972 701190
rect 306996 701188 307052 701190
rect 307076 701188 307132 701190
rect 307156 701188 307212 701190
rect 307236 701188 307292 701190
rect 307316 701188 307372 701190
rect 292578 700168 292634 700224
rect 263598 699488 263654 699544
rect 261390 698944 261446 699000
rect 263690 699352 263746 699408
rect 263690 699080 263746 699136
rect 263874 698944 263930 699000
rect 263690 698844 263692 698864
rect 263692 698844 263744 698864
rect 263744 698844 263746 698864
rect 263690 698808 263746 698844
rect 270498 699796 270500 699816
rect 270500 699796 270552 699816
rect 270552 699796 270554 699816
rect 270498 699760 270554 699796
rect 273166 699760 273222 699816
rect 273350 699388 273352 699408
rect 273352 699388 273404 699408
rect 273404 699388 273406 699408
rect 273350 699352 273406 699388
rect 273258 699080 273314 699136
rect 270836 699066 270892 699068
rect 270916 699066 270972 699068
rect 270996 699066 271052 699068
rect 271076 699066 271132 699068
rect 271156 699066 271212 699068
rect 271236 699066 271292 699068
rect 271316 699066 271372 699068
rect 270836 699014 270874 699066
rect 270874 699014 270886 699066
rect 270886 699014 270892 699066
rect 270916 699014 270938 699066
rect 270938 699014 270950 699066
rect 270950 699014 270972 699066
rect 270996 699014 271002 699066
rect 271002 699014 271014 699066
rect 271014 699014 271052 699066
rect 271076 699014 271078 699066
rect 271078 699014 271130 699066
rect 271130 699014 271132 699066
rect 271156 699014 271194 699066
rect 271194 699014 271206 699066
rect 271206 699014 271212 699066
rect 271236 699014 271258 699066
rect 271258 699014 271270 699066
rect 271270 699014 271292 699066
rect 271316 699014 271322 699066
rect 271322 699014 271334 699066
rect 271334 699014 271372 699066
rect 270836 699012 270892 699014
rect 270916 699012 270972 699014
rect 270996 699012 271052 699014
rect 271076 699012 271132 699014
rect 271156 699012 271212 699014
rect 271236 699012 271292 699014
rect 271316 699012 271372 699014
rect 273534 698944 273590 699000
rect 289542 700052 289598 700088
rect 298650 700168 298706 700224
rect 289542 700032 289544 700052
rect 289544 700032 289596 700052
rect 289596 700032 289598 700052
rect 282734 699488 282790 699544
rect 282734 699352 282790 699408
rect 282918 699488 282974 699544
rect 283010 699388 283012 699408
rect 283012 699388 283064 699408
rect 283064 699388 283066 699408
rect 283010 699352 283066 699388
rect 282918 698808 282974 698864
rect 283286 698944 283342 699000
rect 283010 698536 283066 698592
rect 288836 699610 288892 699612
rect 288916 699610 288972 699612
rect 288996 699610 289052 699612
rect 289076 699610 289132 699612
rect 289156 699610 289212 699612
rect 289236 699610 289292 699612
rect 289316 699610 289372 699612
rect 288836 699558 288874 699610
rect 288874 699558 288886 699610
rect 288886 699558 288892 699610
rect 288916 699558 288938 699610
rect 288938 699558 288950 699610
rect 288950 699558 288972 699610
rect 288996 699558 289002 699610
rect 289002 699558 289014 699610
rect 289014 699558 289052 699610
rect 289076 699558 289078 699610
rect 289078 699558 289130 699610
rect 289130 699558 289132 699610
rect 289156 699558 289194 699610
rect 289194 699558 289206 699610
rect 289206 699558 289212 699610
rect 289236 699558 289258 699610
rect 289258 699558 289270 699610
rect 289270 699558 289292 699610
rect 289316 699558 289322 699610
rect 289322 699558 289334 699610
rect 289334 699558 289372 699610
rect 288836 699556 288892 699558
rect 288916 699556 288972 699558
rect 288996 699556 289052 699558
rect 289076 699556 289132 699558
rect 289156 699556 289212 699558
rect 289236 699556 289292 699558
rect 289316 699556 289372 699558
rect 288438 699080 288494 699136
rect 288836 698522 288892 698524
rect 288916 698522 288972 698524
rect 288996 698522 289052 698524
rect 289076 698522 289132 698524
rect 289156 698522 289212 698524
rect 289236 698522 289292 698524
rect 289316 698522 289372 698524
rect 288836 698470 288874 698522
rect 288874 698470 288886 698522
rect 288886 698470 288892 698522
rect 288916 698470 288938 698522
rect 288938 698470 288950 698522
rect 288950 698470 288972 698522
rect 288996 698470 289002 698522
rect 289002 698470 289014 698522
rect 289014 698470 289052 698522
rect 289076 698470 289078 698522
rect 289078 698470 289130 698522
rect 289130 698470 289132 698522
rect 289156 698470 289194 698522
rect 289194 698470 289206 698522
rect 289206 698470 289212 698522
rect 289236 698470 289258 698522
rect 289258 698470 289270 698522
rect 289270 698470 289292 698522
rect 289316 698470 289322 698522
rect 289322 698470 289334 698522
rect 289334 698470 289372 698522
rect 288836 698468 288892 698470
rect 288916 698468 288972 698470
rect 288996 698468 289052 698470
rect 289076 698468 289132 698470
rect 289156 698468 289212 698470
rect 289236 698468 289292 698470
rect 289316 698468 289372 698470
rect 292302 699896 292358 699952
rect 292486 699796 292488 699816
rect 292488 699796 292540 699816
rect 292540 699796 292542 699816
rect 292486 699760 292542 699796
rect 292670 699896 292726 699952
rect 289726 699488 289782 699544
rect 292670 699488 292726 699544
rect 294050 699352 294106 699408
rect 292394 699116 292396 699136
rect 292396 699116 292448 699136
rect 292448 699116 292450 699136
rect 292394 699080 292450 699116
rect 292486 698944 292542 699000
rect 306836 700154 306892 700156
rect 306916 700154 306972 700156
rect 306996 700154 307052 700156
rect 307076 700154 307132 700156
rect 307156 700154 307212 700156
rect 307236 700154 307292 700156
rect 307316 700154 307372 700156
rect 306836 700102 306874 700154
rect 306874 700102 306886 700154
rect 306886 700102 306892 700154
rect 306916 700102 306938 700154
rect 306938 700102 306950 700154
rect 306950 700102 306972 700154
rect 306996 700102 307002 700154
rect 307002 700102 307014 700154
rect 307014 700102 307052 700154
rect 307076 700102 307078 700154
rect 307078 700102 307130 700154
rect 307130 700102 307132 700154
rect 307156 700102 307194 700154
rect 307194 700102 307206 700154
rect 307206 700102 307212 700154
rect 307236 700102 307258 700154
rect 307258 700102 307270 700154
rect 307270 700102 307292 700154
rect 307316 700102 307322 700154
rect 307322 700102 307334 700154
rect 307334 700102 307372 700154
rect 306836 700100 306892 700102
rect 306916 700100 306972 700102
rect 306996 700100 307052 700102
rect 307076 700100 307132 700102
rect 307156 700100 307212 700102
rect 307236 700100 307292 700102
rect 307316 700100 307372 700102
rect 302054 699916 302110 699952
rect 302054 699896 302056 699916
rect 302056 699896 302108 699916
rect 302108 699896 302110 699916
rect 303618 699896 303674 699952
rect 301962 699796 301964 699816
rect 301964 699796 302016 699816
rect 302016 699796 302018 699816
rect 301962 699760 302018 699796
rect 302146 699080 302202 699136
rect 300214 698808 300270 698864
rect 306836 699066 306892 699068
rect 306916 699066 306972 699068
rect 306996 699066 307052 699068
rect 307076 699066 307132 699068
rect 307156 699066 307212 699068
rect 307236 699066 307292 699068
rect 307316 699066 307372 699068
rect 306836 699014 306874 699066
rect 306874 699014 306886 699066
rect 306886 699014 306892 699066
rect 306916 699014 306938 699066
rect 306938 699014 306950 699066
rect 306950 699014 306972 699066
rect 306996 699014 307002 699066
rect 307002 699014 307014 699066
rect 307014 699014 307052 699066
rect 307076 699014 307078 699066
rect 307078 699014 307130 699066
rect 307130 699014 307132 699066
rect 307156 699014 307194 699066
rect 307194 699014 307206 699066
rect 307206 699014 307212 699066
rect 307236 699014 307258 699066
rect 307258 699014 307270 699066
rect 307270 699014 307292 699066
rect 307316 699014 307322 699066
rect 307322 699014 307334 699066
rect 307334 699014 307372 699066
rect 306836 699012 306892 699014
rect 306916 699012 306972 699014
rect 306996 699012 307052 699014
rect 307076 699012 307132 699014
rect 307156 699012 307212 699014
rect 307236 699012 307292 699014
rect 307316 699012 307372 699014
rect 306378 698844 306380 698864
rect 306380 698844 306432 698864
rect 306432 698844 306434 698864
rect 306378 698808 306434 698844
rect 311898 699080 311954 699136
rect 324836 700698 324892 700700
rect 324916 700698 324972 700700
rect 324996 700698 325052 700700
rect 325076 700698 325132 700700
rect 325156 700698 325212 700700
rect 325236 700698 325292 700700
rect 325316 700698 325372 700700
rect 324836 700646 324874 700698
rect 324874 700646 324886 700698
rect 324886 700646 324892 700698
rect 324916 700646 324938 700698
rect 324938 700646 324950 700698
rect 324950 700646 324972 700698
rect 324996 700646 325002 700698
rect 325002 700646 325014 700698
rect 325014 700646 325052 700698
rect 325076 700646 325078 700698
rect 325078 700646 325130 700698
rect 325130 700646 325132 700698
rect 325156 700646 325194 700698
rect 325194 700646 325206 700698
rect 325206 700646 325212 700698
rect 325236 700646 325258 700698
rect 325258 700646 325270 700698
rect 325270 700646 325292 700698
rect 325316 700646 325322 700698
rect 325322 700646 325334 700698
rect 325334 700646 325372 700698
rect 324836 700644 324892 700646
rect 324916 700644 324972 700646
rect 324996 700644 325052 700646
rect 325076 700644 325132 700646
rect 325156 700644 325212 700646
rect 325236 700644 325292 700646
rect 325316 700644 325372 700646
rect 324836 699610 324892 699612
rect 324916 699610 324972 699612
rect 324996 699610 325052 699612
rect 325076 699610 325132 699612
rect 325156 699610 325212 699612
rect 325236 699610 325292 699612
rect 325316 699610 325372 699612
rect 324836 699558 324874 699610
rect 324874 699558 324886 699610
rect 324886 699558 324892 699610
rect 324916 699558 324938 699610
rect 324938 699558 324950 699610
rect 324950 699558 324972 699610
rect 324996 699558 325002 699610
rect 325002 699558 325014 699610
rect 325014 699558 325052 699610
rect 325076 699558 325078 699610
rect 325078 699558 325130 699610
rect 325130 699558 325132 699610
rect 325156 699558 325194 699610
rect 325194 699558 325206 699610
rect 325206 699558 325212 699610
rect 325236 699558 325258 699610
rect 325258 699558 325270 699610
rect 325270 699558 325292 699610
rect 325316 699558 325322 699610
rect 325322 699558 325334 699610
rect 325334 699558 325372 699610
rect 324836 699556 324892 699558
rect 324916 699556 324972 699558
rect 324996 699556 325052 699558
rect 325076 699556 325132 699558
rect 325156 699556 325212 699558
rect 325236 699556 325292 699558
rect 325316 699556 325372 699558
rect 325514 699116 325516 699136
rect 325516 699116 325568 699136
rect 325568 699116 325570 699136
rect 325514 699080 325570 699116
rect 325698 699116 325700 699136
rect 325700 699116 325752 699136
rect 325752 699116 325754 699136
rect 325698 699080 325754 699116
rect 325606 698844 325608 698864
rect 325608 698844 325660 698864
rect 325660 698844 325662 698864
rect 325606 698808 325662 698844
rect 324836 698522 324892 698524
rect 324916 698522 324972 698524
rect 324996 698522 325052 698524
rect 325076 698522 325132 698524
rect 325156 698522 325212 698524
rect 325236 698522 325292 698524
rect 325316 698522 325372 698524
rect 324836 698470 324874 698522
rect 324874 698470 324886 698522
rect 324886 698470 324892 698522
rect 324916 698470 324938 698522
rect 324938 698470 324950 698522
rect 324950 698470 324972 698522
rect 324996 698470 325002 698522
rect 325002 698470 325014 698522
rect 325014 698470 325052 698522
rect 325076 698470 325078 698522
rect 325078 698470 325130 698522
rect 325130 698470 325132 698522
rect 325156 698470 325194 698522
rect 325194 698470 325206 698522
rect 325206 698470 325212 698522
rect 325236 698470 325258 698522
rect 325258 698470 325270 698522
rect 325270 698470 325292 698522
rect 325316 698470 325322 698522
rect 325322 698470 325334 698522
rect 325334 698470 325372 698522
rect 324836 698468 324892 698470
rect 324916 698468 324972 698470
rect 324996 698468 325052 698470
rect 325076 698468 325132 698470
rect 325156 698468 325212 698470
rect 325236 698468 325292 698470
rect 325316 698468 325372 698470
rect 331218 699080 331274 699136
rect 342836 701242 342892 701244
rect 342916 701242 342972 701244
rect 342996 701242 343052 701244
rect 343076 701242 343132 701244
rect 343156 701242 343212 701244
rect 343236 701242 343292 701244
rect 343316 701242 343372 701244
rect 342836 701190 342874 701242
rect 342874 701190 342886 701242
rect 342886 701190 342892 701242
rect 342916 701190 342938 701242
rect 342938 701190 342950 701242
rect 342950 701190 342972 701242
rect 342996 701190 343002 701242
rect 343002 701190 343014 701242
rect 343014 701190 343052 701242
rect 343076 701190 343078 701242
rect 343078 701190 343130 701242
rect 343130 701190 343132 701242
rect 343156 701190 343194 701242
rect 343194 701190 343206 701242
rect 343206 701190 343212 701242
rect 343236 701190 343258 701242
rect 343258 701190 343270 701242
rect 343270 701190 343292 701242
rect 343316 701190 343322 701242
rect 343322 701190 343334 701242
rect 343334 701190 343372 701242
rect 342836 701188 342892 701190
rect 342916 701188 342972 701190
rect 342996 701188 343052 701190
rect 343076 701188 343132 701190
rect 343156 701188 343212 701190
rect 343236 701188 343292 701190
rect 343316 701188 343372 701190
rect 336922 700984 336978 701040
rect 346306 700440 346362 700496
rect 341614 700304 341670 700360
rect 340694 698844 340696 698864
rect 340696 698844 340748 698864
rect 340748 698844 340750 698864
rect 340694 698808 340750 698844
rect 342836 700154 342892 700156
rect 342916 700154 342972 700156
rect 342996 700154 343052 700156
rect 343076 700154 343132 700156
rect 343156 700154 343212 700156
rect 343236 700154 343292 700156
rect 343316 700154 343372 700156
rect 342836 700102 342874 700154
rect 342874 700102 342886 700154
rect 342886 700102 342892 700154
rect 342916 700102 342938 700154
rect 342938 700102 342950 700154
rect 342950 700102 342972 700154
rect 342996 700102 343002 700154
rect 343002 700102 343014 700154
rect 343014 700102 343052 700154
rect 343076 700102 343078 700154
rect 343078 700102 343130 700154
rect 343130 700102 343132 700154
rect 343156 700102 343194 700154
rect 343194 700102 343206 700154
rect 343206 700102 343212 700154
rect 343236 700102 343258 700154
rect 343258 700102 343270 700154
rect 343270 700102 343292 700154
rect 343316 700102 343322 700154
rect 343322 700102 343334 700154
rect 343334 700102 343372 700154
rect 342836 700100 342892 700102
rect 342916 700100 342972 700102
rect 342996 700100 343052 700102
rect 343076 700100 343132 700102
rect 343156 700100 343212 700102
rect 343236 700100 343292 700102
rect 343316 700100 343372 700102
rect 343546 699080 343602 699136
rect 342836 699066 342892 699068
rect 342916 699066 342972 699068
rect 342996 699066 343052 699068
rect 343076 699066 343132 699068
rect 343156 699066 343212 699068
rect 343236 699066 343292 699068
rect 343316 699066 343372 699068
rect 342836 699014 342874 699066
rect 342874 699014 342886 699066
rect 342886 699014 342892 699066
rect 342916 699014 342938 699066
rect 342938 699014 342950 699066
rect 342950 699014 342972 699066
rect 342996 699014 343002 699066
rect 343002 699014 343014 699066
rect 343014 699014 343052 699066
rect 343076 699014 343078 699066
rect 343078 699014 343130 699066
rect 343130 699014 343132 699066
rect 343156 699014 343194 699066
rect 343194 699014 343206 699066
rect 343206 699014 343212 699066
rect 343236 699014 343258 699066
rect 343258 699014 343270 699066
rect 343270 699014 343292 699066
rect 343316 699014 343322 699066
rect 343322 699014 343334 699066
rect 343334 699014 343372 699066
rect 342836 699012 342892 699014
rect 342916 699012 342972 699014
rect 342996 699012 343052 699014
rect 343076 699012 343132 699014
rect 343156 699012 343212 699014
rect 343236 699012 343292 699014
rect 343316 699012 343372 699014
rect 360836 701786 360892 701788
rect 360916 701786 360972 701788
rect 360996 701786 361052 701788
rect 361076 701786 361132 701788
rect 361156 701786 361212 701788
rect 361236 701786 361292 701788
rect 361316 701786 361372 701788
rect 360836 701734 360874 701786
rect 360874 701734 360886 701786
rect 360886 701734 360892 701786
rect 360916 701734 360938 701786
rect 360938 701734 360950 701786
rect 360950 701734 360972 701786
rect 360996 701734 361002 701786
rect 361002 701734 361014 701786
rect 361014 701734 361052 701786
rect 361076 701734 361078 701786
rect 361078 701734 361130 701786
rect 361130 701734 361132 701786
rect 361156 701734 361194 701786
rect 361194 701734 361206 701786
rect 361206 701734 361212 701786
rect 361236 701734 361258 701786
rect 361258 701734 361270 701786
rect 361270 701734 361292 701786
rect 361316 701734 361322 701786
rect 361322 701734 361334 701786
rect 361334 701734 361372 701786
rect 360836 701732 360892 701734
rect 360916 701732 360972 701734
rect 360996 701732 361052 701734
rect 361076 701732 361132 701734
rect 361156 701732 361212 701734
rect 361236 701732 361292 701734
rect 361316 701732 361372 701734
rect 360836 700698 360892 700700
rect 360916 700698 360972 700700
rect 360996 700698 361052 700700
rect 361076 700698 361132 700700
rect 361156 700698 361212 700700
rect 361236 700698 361292 700700
rect 361316 700698 361372 700700
rect 360836 700646 360874 700698
rect 360874 700646 360886 700698
rect 360886 700646 360892 700698
rect 360916 700646 360938 700698
rect 360938 700646 360950 700698
rect 360950 700646 360972 700698
rect 360996 700646 361002 700698
rect 361002 700646 361014 700698
rect 361014 700646 361052 700698
rect 361076 700646 361078 700698
rect 361078 700646 361130 700698
rect 361130 700646 361132 700698
rect 361156 700646 361194 700698
rect 361194 700646 361206 700698
rect 361206 700646 361212 700698
rect 361236 700646 361258 700698
rect 361258 700646 361270 700698
rect 361270 700646 361292 700698
rect 361316 700646 361322 700698
rect 361322 700646 361334 700698
rect 361334 700646 361372 700698
rect 360836 700644 360892 700646
rect 360916 700644 360972 700646
rect 360996 700644 361052 700646
rect 361076 700644 361132 700646
rect 361156 700644 361212 700646
rect 361236 700644 361292 700646
rect 361316 700644 361372 700646
rect 396836 701786 396892 701788
rect 396916 701786 396972 701788
rect 396996 701786 397052 701788
rect 397076 701786 397132 701788
rect 397156 701786 397212 701788
rect 397236 701786 397292 701788
rect 397316 701786 397372 701788
rect 396836 701734 396874 701786
rect 396874 701734 396886 701786
rect 396886 701734 396892 701786
rect 396916 701734 396938 701786
rect 396938 701734 396950 701786
rect 396950 701734 396972 701786
rect 396996 701734 397002 701786
rect 397002 701734 397014 701786
rect 397014 701734 397052 701786
rect 397076 701734 397078 701786
rect 397078 701734 397130 701786
rect 397130 701734 397132 701786
rect 397156 701734 397194 701786
rect 397194 701734 397206 701786
rect 397206 701734 397212 701786
rect 397236 701734 397258 701786
rect 397258 701734 397270 701786
rect 397270 701734 397292 701786
rect 397316 701734 397322 701786
rect 397322 701734 397334 701786
rect 397334 701734 397372 701786
rect 396836 701732 396892 701734
rect 396916 701732 396972 701734
rect 396996 701732 397052 701734
rect 397076 701732 397132 701734
rect 397156 701732 397212 701734
rect 397236 701732 397292 701734
rect 397316 701732 397372 701734
rect 378836 701242 378892 701244
rect 378916 701242 378972 701244
rect 378996 701242 379052 701244
rect 379076 701242 379132 701244
rect 379156 701242 379212 701244
rect 379236 701242 379292 701244
rect 379316 701242 379372 701244
rect 378836 701190 378874 701242
rect 378874 701190 378886 701242
rect 378886 701190 378892 701242
rect 378916 701190 378938 701242
rect 378938 701190 378950 701242
rect 378950 701190 378972 701242
rect 378996 701190 379002 701242
rect 379002 701190 379014 701242
rect 379014 701190 379052 701242
rect 379076 701190 379078 701242
rect 379078 701190 379130 701242
rect 379130 701190 379132 701242
rect 379156 701190 379194 701242
rect 379194 701190 379206 701242
rect 379206 701190 379212 701242
rect 379236 701190 379258 701242
rect 379258 701190 379270 701242
rect 379270 701190 379292 701242
rect 379316 701190 379322 701242
rect 379322 701190 379334 701242
rect 379334 701190 379372 701242
rect 378836 701188 378892 701190
rect 378916 701188 378972 701190
rect 378996 701188 379052 701190
rect 379076 701188 379132 701190
rect 379156 701188 379212 701190
rect 379236 701188 379292 701190
rect 379316 701188 379372 701190
rect 396836 700698 396892 700700
rect 396916 700698 396972 700700
rect 396996 700698 397052 700700
rect 397076 700698 397132 700700
rect 397156 700698 397212 700700
rect 397236 700698 397292 700700
rect 397316 700698 397372 700700
rect 396836 700646 396874 700698
rect 396874 700646 396886 700698
rect 396886 700646 396892 700698
rect 396916 700646 396938 700698
rect 396938 700646 396950 700698
rect 396950 700646 396972 700698
rect 396996 700646 397002 700698
rect 397002 700646 397014 700698
rect 397014 700646 397052 700698
rect 397076 700646 397078 700698
rect 397078 700646 397130 700698
rect 397130 700646 397132 700698
rect 397156 700646 397194 700698
rect 397194 700646 397206 700698
rect 397206 700646 397212 700698
rect 397236 700646 397258 700698
rect 397258 700646 397270 700698
rect 397270 700646 397292 700698
rect 397316 700646 397322 700698
rect 397322 700646 397334 700698
rect 397334 700646 397372 700698
rect 396836 700644 396892 700646
rect 396916 700644 396972 700646
rect 396996 700644 397052 700646
rect 397076 700644 397132 700646
rect 397156 700644 397212 700646
rect 397236 700644 397292 700646
rect 397316 700644 397372 700646
rect 378836 700154 378892 700156
rect 378916 700154 378972 700156
rect 378996 700154 379052 700156
rect 379076 700154 379132 700156
rect 379156 700154 379212 700156
rect 379236 700154 379292 700156
rect 379316 700154 379372 700156
rect 378836 700102 378874 700154
rect 378874 700102 378886 700154
rect 378886 700102 378892 700154
rect 378916 700102 378938 700154
rect 378938 700102 378950 700154
rect 378950 700102 378972 700154
rect 378996 700102 379002 700154
rect 379002 700102 379014 700154
rect 379014 700102 379052 700154
rect 379076 700102 379078 700154
rect 379078 700102 379130 700154
rect 379130 700102 379132 700154
rect 379156 700102 379194 700154
rect 379194 700102 379206 700154
rect 379206 700102 379212 700154
rect 379236 700102 379258 700154
rect 379258 700102 379270 700154
rect 379270 700102 379292 700154
rect 379316 700102 379322 700154
rect 379322 700102 379334 700154
rect 379334 700102 379372 700154
rect 378836 700100 378892 700102
rect 378916 700100 378972 700102
rect 378996 700100 379052 700102
rect 379076 700100 379132 700102
rect 379156 700100 379212 700102
rect 379236 700100 379292 700102
rect 379316 700100 379372 700102
rect 432836 701786 432892 701788
rect 432916 701786 432972 701788
rect 432996 701786 433052 701788
rect 433076 701786 433132 701788
rect 433156 701786 433212 701788
rect 433236 701786 433292 701788
rect 433316 701786 433372 701788
rect 432836 701734 432874 701786
rect 432874 701734 432886 701786
rect 432886 701734 432892 701786
rect 432916 701734 432938 701786
rect 432938 701734 432950 701786
rect 432950 701734 432972 701786
rect 432996 701734 433002 701786
rect 433002 701734 433014 701786
rect 433014 701734 433052 701786
rect 433076 701734 433078 701786
rect 433078 701734 433130 701786
rect 433130 701734 433132 701786
rect 433156 701734 433194 701786
rect 433194 701734 433206 701786
rect 433206 701734 433212 701786
rect 433236 701734 433258 701786
rect 433258 701734 433270 701786
rect 433270 701734 433292 701786
rect 433316 701734 433322 701786
rect 433322 701734 433334 701786
rect 433334 701734 433372 701786
rect 432836 701732 432892 701734
rect 432916 701732 432972 701734
rect 432996 701732 433052 701734
rect 433076 701732 433132 701734
rect 433156 701732 433212 701734
rect 433236 701732 433292 701734
rect 433316 701732 433372 701734
rect 414836 701242 414892 701244
rect 414916 701242 414972 701244
rect 414996 701242 415052 701244
rect 415076 701242 415132 701244
rect 415156 701242 415212 701244
rect 415236 701242 415292 701244
rect 415316 701242 415372 701244
rect 414836 701190 414874 701242
rect 414874 701190 414886 701242
rect 414886 701190 414892 701242
rect 414916 701190 414938 701242
rect 414938 701190 414950 701242
rect 414950 701190 414972 701242
rect 414996 701190 415002 701242
rect 415002 701190 415014 701242
rect 415014 701190 415052 701242
rect 415076 701190 415078 701242
rect 415078 701190 415130 701242
rect 415130 701190 415132 701242
rect 415156 701190 415194 701242
rect 415194 701190 415206 701242
rect 415206 701190 415212 701242
rect 415236 701190 415258 701242
rect 415258 701190 415270 701242
rect 415270 701190 415292 701242
rect 415316 701190 415322 701242
rect 415322 701190 415334 701242
rect 415334 701190 415372 701242
rect 414836 701188 414892 701190
rect 414916 701188 414972 701190
rect 414996 701188 415052 701190
rect 415076 701188 415132 701190
rect 415156 701188 415212 701190
rect 415236 701188 415292 701190
rect 415316 701188 415372 701190
rect 450836 701242 450892 701244
rect 450916 701242 450972 701244
rect 450996 701242 451052 701244
rect 451076 701242 451132 701244
rect 451156 701242 451212 701244
rect 451236 701242 451292 701244
rect 451316 701242 451372 701244
rect 450836 701190 450874 701242
rect 450874 701190 450886 701242
rect 450886 701190 450892 701242
rect 450916 701190 450938 701242
rect 450938 701190 450950 701242
rect 450950 701190 450972 701242
rect 450996 701190 451002 701242
rect 451002 701190 451014 701242
rect 451014 701190 451052 701242
rect 451076 701190 451078 701242
rect 451078 701190 451130 701242
rect 451130 701190 451132 701242
rect 451156 701190 451194 701242
rect 451194 701190 451206 701242
rect 451206 701190 451212 701242
rect 451236 701190 451258 701242
rect 451258 701190 451270 701242
rect 451270 701190 451292 701242
rect 451316 701190 451322 701242
rect 451322 701190 451334 701242
rect 451334 701190 451372 701242
rect 450836 701188 450892 701190
rect 450916 701188 450972 701190
rect 450996 701188 451052 701190
rect 451076 701188 451132 701190
rect 451156 701188 451212 701190
rect 451236 701188 451292 701190
rect 451316 701188 451372 701190
rect 432836 700698 432892 700700
rect 432916 700698 432972 700700
rect 432996 700698 433052 700700
rect 433076 700698 433132 700700
rect 433156 700698 433212 700700
rect 433236 700698 433292 700700
rect 433316 700698 433372 700700
rect 432836 700646 432874 700698
rect 432874 700646 432886 700698
rect 432886 700646 432892 700698
rect 432916 700646 432938 700698
rect 432938 700646 432950 700698
rect 432950 700646 432972 700698
rect 432996 700646 433002 700698
rect 433002 700646 433014 700698
rect 433014 700646 433052 700698
rect 433076 700646 433078 700698
rect 433078 700646 433130 700698
rect 433130 700646 433132 700698
rect 433156 700646 433194 700698
rect 433194 700646 433206 700698
rect 433206 700646 433212 700698
rect 433236 700646 433258 700698
rect 433258 700646 433270 700698
rect 433270 700646 433292 700698
rect 433316 700646 433322 700698
rect 433322 700646 433334 700698
rect 433334 700646 433372 700698
rect 432836 700644 432892 700646
rect 432916 700644 432972 700646
rect 432996 700644 433052 700646
rect 433076 700644 433132 700646
rect 433156 700644 433212 700646
rect 433236 700644 433292 700646
rect 433316 700644 433372 700646
rect 468836 701786 468892 701788
rect 468916 701786 468972 701788
rect 468996 701786 469052 701788
rect 469076 701786 469132 701788
rect 469156 701786 469212 701788
rect 469236 701786 469292 701788
rect 469316 701786 469372 701788
rect 468836 701734 468874 701786
rect 468874 701734 468886 701786
rect 468886 701734 468892 701786
rect 468916 701734 468938 701786
rect 468938 701734 468950 701786
rect 468950 701734 468972 701786
rect 468996 701734 469002 701786
rect 469002 701734 469014 701786
rect 469014 701734 469052 701786
rect 469076 701734 469078 701786
rect 469078 701734 469130 701786
rect 469130 701734 469132 701786
rect 469156 701734 469194 701786
rect 469194 701734 469206 701786
rect 469206 701734 469212 701786
rect 469236 701734 469258 701786
rect 469258 701734 469270 701786
rect 469270 701734 469292 701786
rect 469316 701734 469322 701786
rect 469322 701734 469334 701786
rect 469334 701734 469372 701786
rect 468836 701732 468892 701734
rect 468916 701732 468972 701734
rect 468996 701732 469052 701734
rect 469076 701732 469132 701734
rect 469156 701732 469212 701734
rect 469236 701732 469292 701734
rect 469316 701732 469372 701734
rect 468836 700698 468892 700700
rect 468916 700698 468972 700700
rect 468996 700698 469052 700700
rect 469076 700698 469132 700700
rect 469156 700698 469212 700700
rect 469236 700698 469292 700700
rect 469316 700698 469372 700700
rect 468836 700646 468874 700698
rect 468874 700646 468886 700698
rect 468886 700646 468892 700698
rect 468916 700646 468938 700698
rect 468938 700646 468950 700698
rect 468950 700646 468972 700698
rect 468996 700646 469002 700698
rect 469002 700646 469014 700698
rect 469014 700646 469052 700698
rect 469076 700646 469078 700698
rect 469078 700646 469130 700698
rect 469130 700646 469132 700698
rect 469156 700646 469194 700698
rect 469194 700646 469206 700698
rect 469206 700646 469212 700698
rect 469236 700646 469258 700698
rect 469258 700646 469270 700698
rect 469270 700646 469292 700698
rect 469316 700646 469322 700698
rect 469322 700646 469334 700698
rect 469334 700646 469372 700698
rect 468836 700644 468892 700646
rect 468916 700644 468972 700646
rect 468996 700644 469052 700646
rect 469076 700644 469132 700646
rect 469156 700644 469212 700646
rect 469236 700644 469292 700646
rect 469316 700644 469372 700646
rect 504836 701786 504892 701788
rect 504916 701786 504972 701788
rect 504996 701786 505052 701788
rect 505076 701786 505132 701788
rect 505156 701786 505212 701788
rect 505236 701786 505292 701788
rect 505316 701786 505372 701788
rect 504836 701734 504874 701786
rect 504874 701734 504886 701786
rect 504886 701734 504892 701786
rect 504916 701734 504938 701786
rect 504938 701734 504950 701786
rect 504950 701734 504972 701786
rect 504996 701734 505002 701786
rect 505002 701734 505014 701786
rect 505014 701734 505052 701786
rect 505076 701734 505078 701786
rect 505078 701734 505130 701786
rect 505130 701734 505132 701786
rect 505156 701734 505194 701786
rect 505194 701734 505206 701786
rect 505206 701734 505212 701786
rect 505236 701734 505258 701786
rect 505258 701734 505270 701786
rect 505270 701734 505292 701786
rect 505316 701734 505322 701786
rect 505322 701734 505334 701786
rect 505334 701734 505372 701786
rect 504836 701732 504892 701734
rect 504916 701732 504972 701734
rect 504996 701732 505052 701734
rect 505076 701732 505132 701734
rect 505156 701732 505212 701734
rect 505236 701732 505292 701734
rect 505316 701732 505372 701734
rect 486836 701242 486892 701244
rect 486916 701242 486972 701244
rect 486996 701242 487052 701244
rect 487076 701242 487132 701244
rect 487156 701242 487212 701244
rect 487236 701242 487292 701244
rect 487316 701242 487372 701244
rect 486836 701190 486874 701242
rect 486874 701190 486886 701242
rect 486886 701190 486892 701242
rect 486916 701190 486938 701242
rect 486938 701190 486950 701242
rect 486950 701190 486972 701242
rect 486996 701190 487002 701242
rect 487002 701190 487014 701242
rect 487014 701190 487052 701242
rect 487076 701190 487078 701242
rect 487078 701190 487130 701242
rect 487130 701190 487132 701242
rect 487156 701190 487194 701242
rect 487194 701190 487206 701242
rect 487206 701190 487212 701242
rect 487236 701190 487258 701242
rect 487258 701190 487270 701242
rect 487270 701190 487292 701242
rect 487316 701190 487322 701242
rect 487322 701190 487334 701242
rect 487334 701190 487372 701242
rect 486836 701188 486892 701190
rect 486916 701188 486972 701190
rect 486996 701188 487052 701190
rect 487076 701188 487132 701190
rect 487156 701188 487212 701190
rect 487236 701188 487292 701190
rect 487316 701188 487372 701190
rect 522836 701242 522892 701244
rect 522916 701242 522972 701244
rect 522996 701242 523052 701244
rect 523076 701242 523132 701244
rect 523156 701242 523212 701244
rect 523236 701242 523292 701244
rect 523316 701242 523372 701244
rect 522836 701190 522874 701242
rect 522874 701190 522886 701242
rect 522886 701190 522892 701242
rect 522916 701190 522938 701242
rect 522938 701190 522950 701242
rect 522950 701190 522972 701242
rect 522996 701190 523002 701242
rect 523002 701190 523014 701242
rect 523014 701190 523052 701242
rect 523076 701190 523078 701242
rect 523078 701190 523130 701242
rect 523130 701190 523132 701242
rect 523156 701190 523194 701242
rect 523194 701190 523206 701242
rect 523206 701190 523212 701242
rect 523236 701190 523258 701242
rect 523258 701190 523270 701242
rect 523270 701190 523292 701242
rect 523316 701190 523322 701242
rect 523322 701190 523334 701242
rect 523334 701190 523372 701242
rect 522836 701188 522892 701190
rect 522916 701188 522972 701190
rect 522996 701188 523052 701190
rect 523076 701188 523132 701190
rect 523156 701188 523212 701190
rect 523236 701188 523292 701190
rect 523316 701188 523372 701190
rect 540836 701786 540892 701788
rect 540916 701786 540972 701788
rect 540996 701786 541052 701788
rect 541076 701786 541132 701788
rect 541156 701786 541212 701788
rect 541236 701786 541292 701788
rect 541316 701786 541372 701788
rect 540836 701734 540874 701786
rect 540874 701734 540886 701786
rect 540886 701734 540892 701786
rect 540916 701734 540938 701786
rect 540938 701734 540950 701786
rect 540950 701734 540972 701786
rect 540996 701734 541002 701786
rect 541002 701734 541014 701786
rect 541014 701734 541052 701786
rect 541076 701734 541078 701786
rect 541078 701734 541130 701786
rect 541130 701734 541132 701786
rect 541156 701734 541194 701786
rect 541194 701734 541206 701786
rect 541206 701734 541212 701786
rect 541236 701734 541258 701786
rect 541258 701734 541270 701786
rect 541270 701734 541292 701786
rect 541316 701734 541322 701786
rect 541322 701734 541334 701786
rect 541334 701734 541372 701786
rect 540836 701732 540892 701734
rect 540916 701732 540972 701734
rect 540996 701732 541052 701734
rect 541076 701732 541132 701734
rect 541156 701732 541212 701734
rect 541236 701732 541292 701734
rect 541316 701732 541372 701734
rect 527178 700848 527234 700904
rect 504836 700698 504892 700700
rect 504916 700698 504972 700700
rect 504996 700698 505052 700700
rect 505076 700698 505132 700700
rect 505156 700698 505212 700700
rect 505236 700698 505292 700700
rect 505316 700698 505372 700700
rect 504836 700646 504874 700698
rect 504874 700646 504886 700698
rect 504886 700646 504892 700698
rect 504916 700646 504938 700698
rect 504938 700646 504950 700698
rect 504950 700646 504972 700698
rect 504996 700646 505002 700698
rect 505002 700646 505014 700698
rect 505014 700646 505052 700698
rect 505076 700646 505078 700698
rect 505078 700646 505130 700698
rect 505130 700646 505132 700698
rect 505156 700646 505194 700698
rect 505194 700646 505206 700698
rect 505206 700646 505212 700698
rect 505236 700646 505258 700698
rect 505258 700646 505270 700698
rect 505270 700646 505292 700698
rect 505316 700646 505322 700698
rect 505322 700646 505334 700698
rect 505334 700646 505372 700698
rect 504836 700644 504892 700646
rect 504916 700644 504972 700646
rect 504996 700644 505052 700646
rect 505076 700644 505132 700646
rect 505156 700644 505212 700646
rect 505236 700644 505292 700646
rect 505316 700644 505372 700646
rect 540836 700698 540892 700700
rect 540916 700698 540972 700700
rect 540996 700698 541052 700700
rect 541076 700698 541132 700700
rect 541156 700698 541212 700700
rect 541236 700698 541292 700700
rect 541316 700698 541372 700700
rect 540836 700646 540874 700698
rect 540874 700646 540886 700698
rect 540886 700646 540892 700698
rect 540916 700646 540938 700698
rect 540938 700646 540950 700698
rect 540950 700646 540972 700698
rect 540996 700646 541002 700698
rect 541002 700646 541014 700698
rect 541014 700646 541052 700698
rect 541076 700646 541078 700698
rect 541078 700646 541130 700698
rect 541130 700646 541132 700698
rect 541156 700646 541194 700698
rect 541194 700646 541206 700698
rect 541206 700646 541212 700698
rect 541236 700646 541258 700698
rect 541258 700646 541270 700698
rect 541270 700646 541292 700698
rect 541316 700646 541322 700698
rect 541322 700646 541334 700698
rect 541334 700646 541372 700698
rect 540836 700644 540892 700646
rect 540916 700644 540972 700646
rect 540996 700644 541052 700646
rect 541076 700644 541132 700646
rect 541156 700644 541212 700646
rect 541236 700644 541292 700646
rect 541316 700644 541372 700646
rect 576836 701786 576892 701788
rect 576916 701786 576972 701788
rect 576996 701786 577052 701788
rect 577076 701786 577132 701788
rect 577156 701786 577212 701788
rect 577236 701786 577292 701788
rect 577316 701786 577372 701788
rect 576836 701734 576874 701786
rect 576874 701734 576886 701786
rect 576886 701734 576892 701786
rect 576916 701734 576938 701786
rect 576938 701734 576950 701786
rect 576950 701734 576972 701786
rect 576996 701734 577002 701786
rect 577002 701734 577014 701786
rect 577014 701734 577052 701786
rect 577076 701734 577078 701786
rect 577078 701734 577130 701786
rect 577130 701734 577132 701786
rect 577156 701734 577194 701786
rect 577194 701734 577206 701786
rect 577206 701734 577212 701786
rect 577236 701734 577258 701786
rect 577258 701734 577270 701786
rect 577270 701734 577292 701786
rect 577316 701734 577322 701786
rect 577322 701734 577334 701786
rect 577334 701734 577372 701786
rect 576836 701732 576892 701734
rect 576916 701732 576972 701734
rect 576996 701732 577052 701734
rect 577076 701732 577132 701734
rect 577156 701732 577212 701734
rect 577236 701732 577292 701734
rect 577316 701732 577372 701734
rect 558836 701242 558892 701244
rect 558916 701242 558972 701244
rect 558996 701242 559052 701244
rect 559076 701242 559132 701244
rect 559156 701242 559212 701244
rect 559236 701242 559292 701244
rect 559316 701242 559372 701244
rect 558836 701190 558874 701242
rect 558874 701190 558886 701242
rect 558886 701190 558892 701242
rect 558916 701190 558938 701242
rect 558938 701190 558950 701242
rect 558950 701190 558972 701242
rect 558996 701190 559002 701242
rect 559002 701190 559014 701242
rect 559014 701190 559052 701242
rect 559076 701190 559078 701242
rect 559078 701190 559130 701242
rect 559130 701190 559132 701242
rect 559156 701190 559194 701242
rect 559194 701190 559206 701242
rect 559206 701190 559212 701242
rect 559236 701190 559258 701242
rect 559258 701190 559270 701242
rect 559270 701190 559292 701242
rect 559316 701190 559322 701242
rect 559322 701190 559334 701242
rect 559334 701190 559372 701242
rect 558836 701188 558892 701190
rect 558916 701188 558972 701190
rect 558996 701188 559052 701190
rect 559076 701188 559132 701190
rect 559156 701188 559212 701190
rect 559236 701188 559292 701190
rect 559316 701188 559372 701190
rect 576836 700698 576892 700700
rect 576916 700698 576972 700700
rect 576996 700698 577052 700700
rect 577076 700698 577132 700700
rect 577156 700698 577212 700700
rect 577236 700698 577292 700700
rect 577316 700698 577372 700700
rect 576836 700646 576874 700698
rect 576874 700646 576886 700698
rect 576886 700646 576892 700698
rect 576916 700646 576938 700698
rect 576938 700646 576950 700698
rect 576950 700646 576972 700698
rect 576996 700646 577002 700698
rect 577002 700646 577014 700698
rect 577014 700646 577052 700698
rect 577076 700646 577078 700698
rect 577078 700646 577130 700698
rect 577130 700646 577132 700698
rect 577156 700646 577194 700698
rect 577194 700646 577206 700698
rect 577206 700646 577212 700698
rect 577236 700646 577258 700698
rect 577258 700646 577270 700698
rect 577270 700646 577292 700698
rect 577316 700646 577322 700698
rect 577322 700646 577334 700698
rect 577334 700646 577372 700698
rect 576836 700644 576892 700646
rect 576916 700644 576972 700646
rect 576996 700644 577052 700646
rect 577076 700644 577132 700646
rect 577156 700644 577212 700646
rect 577236 700644 577292 700646
rect 577316 700644 577372 700646
rect 414836 700154 414892 700156
rect 414916 700154 414972 700156
rect 414996 700154 415052 700156
rect 415076 700154 415132 700156
rect 415156 700154 415212 700156
rect 415236 700154 415292 700156
rect 415316 700154 415372 700156
rect 414836 700102 414874 700154
rect 414874 700102 414886 700154
rect 414886 700102 414892 700154
rect 414916 700102 414938 700154
rect 414938 700102 414950 700154
rect 414950 700102 414972 700154
rect 414996 700102 415002 700154
rect 415002 700102 415014 700154
rect 415014 700102 415052 700154
rect 415076 700102 415078 700154
rect 415078 700102 415130 700154
rect 415130 700102 415132 700154
rect 415156 700102 415194 700154
rect 415194 700102 415206 700154
rect 415206 700102 415212 700154
rect 415236 700102 415258 700154
rect 415258 700102 415270 700154
rect 415270 700102 415292 700154
rect 415316 700102 415322 700154
rect 415322 700102 415334 700154
rect 415334 700102 415372 700154
rect 414836 700100 414892 700102
rect 414916 700100 414972 700102
rect 414996 700100 415052 700102
rect 415076 700100 415132 700102
rect 415156 700100 415212 700102
rect 415236 700100 415292 700102
rect 415316 700100 415372 700102
rect 450836 700154 450892 700156
rect 450916 700154 450972 700156
rect 450996 700154 451052 700156
rect 451076 700154 451132 700156
rect 451156 700154 451212 700156
rect 451236 700154 451292 700156
rect 451316 700154 451372 700156
rect 450836 700102 450874 700154
rect 450874 700102 450886 700154
rect 450886 700102 450892 700154
rect 450916 700102 450938 700154
rect 450938 700102 450950 700154
rect 450950 700102 450972 700154
rect 450996 700102 451002 700154
rect 451002 700102 451014 700154
rect 451014 700102 451052 700154
rect 451076 700102 451078 700154
rect 451078 700102 451130 700154
rect 451130 700102 451132 700154
rect 451156 700102 451194 700154
rect 451194 700102 451206 700154
rect 451206 700102 451212 700154
rect 451236 700102 451258 700154
rect 451258 700102 451270 700154
rect 451270 700102 451292 700154
rect 451316 700102 451322 700154
rect 451322 700102 451334 700154
rect 451334 700102 451372 700154
rect 450836 700100 450892 700102
rect 450916 700100 450972 700102
rect 450996 700100 451052 700102
rect 451076 700100 451132 700102
rect 451156 700100 451212 700102
rect 451236 700100 451292 700102
rect 451316 700100 451372 700102
rect 486836 700154 486892 700156
rect 486916 700154 486972 700156
rect 486996 700154 487052 700156
rect 487076 700154 487132 700156
rect 487156 700154 487212 700156
rect 487236 700154 487292 700156
rect 487316 700154 487372 700156
rect 486836 700102 486874 700154
rect 486874 700102 486886 700154
rect 486886 700102 486892 700154
rect 486916 700102 486938 700154
rect 486938 700102 486950 700154
rect 486950 700102 486972 700154
rect 486996 700102 487002 700154
rect 487002 700102 487014 700154
rect 487014 700102 487052 700154
rect 487076 700102 487078 700154
rect 487078 700102 487130 700154
rect 487130 700102 487132 700154
rect 487156 700102 487194 700154
rect 487194 700102 487206 700154
rect 487206 700102 487212 700154
rect 487236 700102 487258 700154
rect 487258 700102 487270 700154
rect 487270 700102 487292 700154
rect 487316 700102 487322 700154
rect 487322 700102 487334 700154
rect 487334 700102 487372 700154
rect 486836 700100 486892 700102
rect 486916 700100 486972 700102
rect 486996 700100 487052 700102
rect 487076 700100 487132 700102
rect 487156 700100 487212 700102
rect 487236 700100 487292 700102
rect 487316 700100 487372 700102
rect 522836 700154 522892 700156
rect 522916 700154 522972 700156
rect 522996 700154 523052 700156
rect 523076 700154 523132 700156
rect 523156 700154 523212 700156
rect 523236 700154 523292 700156
rect 523316 700154 523372 700156
rect 522836 700102 522874 700154
rect 522874 700102 522886 700154
rect 522886 700102 522892 700154
rect 522916 700102 522938 700154
rect 522938 700102 522950 700154
rect 522950 700102 522972 700154
rect 522996 700102 523002 700154
rect 523002 700102 523014 700154
rect 523014 700102 523052 700154
rect 523076 700102 523078 700154
rect 523078 700102 523130 700154
rect 523130 700102 523132 700154
rect 523156 700102 523194 700154
rect 523194 700102 523206 700154
rect 523206 700102 523212 700154
rect 523236 700102 523258 700154
rect 523258 700102 523270 700154
rect 523270 700102 523292 700154
rect 523316 700102 523322 700154
rect 523322 700102 523334 700154
rect 523334 700102 523372 700154
rect 522836 700100 522892 700102
rect 522916 700100 522972 700102
rect 522996 700100 523052 700102
rect 523076 700100 523132 700102
rect 523156 700100 523212 700102
rect 523236 700100 523292 700102
rect 523316 700100 523372 700102
rect 558836 700154 558892 700156
rect 558916 700154 558972 700156
rect 558996 700154 559052 700156
rect 559076 700154 559132 700156
rect 559156 700154 559212 700156
rect 559236 700154 559292 700156
rect 559316 700154 559372 700156
rect 558836 700102 558874 700154
rect 558874 700102 558886 700154
rect 558886 700102 558892 700154
rect 558916 700102 558938 700154
rect 558938 700102 558950 700154
rect 558950 700102 558972 700154
rect 558996 700102 559002 700154
rect 559002 700102 559014 700154
rect 559014 700102 559052 700154
rect 559076 700102 559078 700154
rect 559078 700102 559130 700154
rect 559130 700102 559132 700154
rect 559156 700102 559194 700154
rect 559194 700102 559206 700154
rect 559206 700102 559212 700154
rect 559236 700102 559258 700154
rect 559258 700102 559270 700154
rect 559270 700102 559292 700154
rect 559316 700102 559322 700154
rect 559322 700102 559334 700154
rect 559334 700102 559372 700154
rect 558836 700100 558892 700102
rect 558916 700100 558972 700102
rect 558996 700100 559052 700102
rect 559076 700100 559132 700102
rect 559156 700100 559212 700102
rect 559236 700100 559292 700102
rect 559316 700100 559372 700102
rect 360836 699610 360892 699612
rect 360916 699610 360972 699612
rect 360996 699610 361052 699612
rect 361076 699610 361132 699612
rect 361156 699610 361212 699612
rect 361236 699610 361292 699612
rect 361316 699610 361372 699612
rect 360836 699558 360874 699610
rect 360874 699558 360886 699610
rect 360886 699558 360892 699610
rect 360916 699558 360938 699610
rect 360938 699558 360950 699610
rect 360950 699558 360972 699610
rect 360996 699558 361002 699610
rect 361002 699558 361014 699610
rect 361014 699558 361052 699610
rect 361076 699558 361078 699610
rect 361078 699558 361130 699610
rect 361130 699558 361132 699610
rect 361156 699558 361194 699610
rect 361194 699558 361206 699610
rect 361206 699558 361212 699610
rect 361236 699558 361258 699610
rect 361258 699558 361270 699610
rect 361270 699558 361292 699610
rect 361316 699558 361322 699610
rect 361322 699558 361334 699610
rect 361334 699558 361372 699610
rect 360836 699556 360892 699558
rect 360916 699556 360972 699558
rect 360996 699556 361052 699558
rect 361076 699556 361132 699558
rect 361156 699556 361212 699558
rect 361236 699556 361292 699558
rect 361316 699556 361372 699558
rect 354494 699116 354496 699136
rect 354496 699116 354548 699136
rect 354548 699116 354550 699136
rect 354494 699080 354550 699116
rect 354586 698844 354588 698864
rect 354588 698844 354640 698864
rect 354640 698844 354642 698864
rect 354586 698808 354642 698844
rect 360836 698522 360892 698524
rect 360916 698522 360972 698524
rect 360996 698522 361052 698524
rect 361076 698522 361132 698524
rect 361156 698522 361212 698524
rect 361236 698522 361292 698524
rect 361316 698522 361372 698524
rect 360836 698470 360874 698522
rect 360874 698470 360886 698522
rect 360886 698470 360892 698522
rect 360916 698470 360938 698522
rect 360938 698470 360950 698522
rect 360950 698470 360972 698522
rect 360996 698470 361002 698522
rect 361002 698470 361014 698522
rect 361014 698470 361052 698522
rect 361076 698470 361078 698522
rect 361078 698470 361130 698522
rect 361130 698470 361132 698522
rect 361156 698470 361194 698522
rect 361194 698470 361206 698522
rect 361206 698470 361212 698522
rect 361236 698470 361258 698522
rect 361258 698470 361270 698522
rect 361270 698470 361292 698522
rect 361316 698470 361322 698522
rect 361322 698470 361334 698522
rect 361334 698470 361372 698522
rect 360836 698468 360892 698470
rect 360916 698468 360972 698470
rect 360996 698468 361052 698470
rect 361076 698468 361132 698470
rect 361156 698468 361212 698470
rect 361236 698468 361292 698470
rect 361316 698468 361372 698470
rect 396836 699610 396892 699612
rect 396916 699610 396972 699612
rect 396996 699610 397052 699612
rect 397076 699610 397132 699612
rect 397156 699610 397212 699612
rect 397236 699610 397292 699612
rect 397316 699610 397372 699612
rect 396836 699558 396874 699610
rect 396874 699558 396886 699610
rect 396886 699558 396892 699610
rect 396916 699558 396938 699610
rect 396938 699558 396950 699610
rect 396950 699558 396972 699610
rect 396996 699558 397002 699610
rect 397002 699558 397014 699610
rect 397014 699558 397052 699610
rect 397076 699558 397078 699610
rect 397078 699558 397130 699610
rect 397130 699558 397132 699610
rect 397156 699558 397194 699610
rect 397194 699558 397206 699610
rect 397206 699558 397212 699610
rect 397236 699558 397258 699610
rect 397258 699558 397270 699610
rect 397270 699558 397292 699610
rect 397316 699558 397322 699610
rect 397322 699558 397334 699610
rect 397334 699558 397372 699610
rect 396836 699556 396892 699558
rect 396916 699556 396972 699558
rect 396996 699556 397052 699558
rect 397076 699556 397132 699558
rect 397156 699556 397212 699558
rect 397236 699556 397292 699558
rect 397316 699556 397372 699558
rect 432836 699610 432892 699612
rect 432916 699610 432972 699612
rect 432996 699610 433052 699612
rect 433076 699610 433132 699612
rect 433156 699610 433212 699612
rect 433236 699610 433292 699612
rect 433316 699610 433372 699612
rect 432836 699558 432874 699610
rect 432874 699558 432886 699610
rect 432886 699558 432892 699610
rect 432916 699558 432938 699610
rect 432938 699558 432950 699610
rect 432950 699558 432972 699610
rect 432996 699558 433002 699610
rect 433002 699558 433014 699610
rect 433014 699558 433052 699610
rect 433076 699558 433078 699610
rect 433078 699558 433130 699610
rect 433130 699558 433132 699610
rect 433156 699558 433194 699610
rect 433194 699558 433206 699610
rect 433206 699558 433212 699610
rect 433236 699558 433258 699610
rect 433258 699558 433270 699610
rect 433270 699558 433292 699610
rect 433316 699558 433322 699610
rect 433322 699558 433334 699610
rect 433334 699558 433372 699610
rect 432836 699556 432892 699558
rect 432916 699556 432972 699558
rect 432996 699556 433052 699558
rect 433076 699556 433132 699558
rect 433156 699556 433212 699558
rect 433236 699556 433292 699558
rect 433316 699556 433372 699558
rect 468836 699610 468892 699612
rect 468916 699610 468972 699612
rect 468996 699610 469052 699612
rect 469076 699610 469132 699612
rect 469156 699610 469212 699612
rect 469236 699610 469292 699612
rect 469316 699610 469372 699612
rect 468836 699558 468874 699610
rect 468874 699558 468886 699610
rect 468886 699558 468892 699610
rect 468916 699558 468938 699610
rect 468938 699558 468950 699610
rect 468950 699558 468972 699610
rect 468996 699558 469002 699610
rect 469002 699558 469014 699610
rect 469014 699558 469052 699610
rect 469076 699558 469078 699610
rect 469078 699558 469130 699610
rect 469130 699558 469132 699610
rect 469156 699558 469194 699610
rect 469194 699558 469206 699610
rect 469206 699558 469212 699610
rect 469236 699558 469258 699610
rect 469258 699558 469270 699610
rect 469270 699558 469292 699610
rect 469316 699558 469322 699610
rect 469322 699558 469334 699610
rect 469334 699558 469372 699610
rect 468836 699556 468892 699558
rect 468916 699556 468972 699558
rect 468996 699556 469052 699558
rect 469076 699556 469132 699558
rect 469156 699556 469212 699558
rect 469236 699556 469292 699558
rect 469316 699556 469372 699558
rect 504836 699610 504892 699612
rect 504916 699610 504972 699612
rect 504996 699610 505052 699612
rect 505076 699610 505132 699612
rect 505156 699610 505212 699612
rect 505236 699610 505292 699612
rect 505316 699610 505372 699612
rect 504836 699558 504874 699610
rect 504874 699558 504886 699610
rect 504886 699558 504892 699610
rect 504916 699558 504938 699610
rect 504938 699558 504950 699610
rect 504950 699558 504972 699610
rect 504996 699558 505002 699610
rect 505002 699558 505014 699610
rect 505014 699558 505052 699610
rect 505076 699558 505078 699610
rect 505078 699558 505130 699610
rect 505130 699558 505132 699610
rect 505156 699558 505194 699610
rect 505194 699558 505206 699610
rect 505206 699558 505212 699610
rect 505236 699558 505258 699610
rect 505258 699558 505270 699610
rect 505270 699558 505292 699610
rect 505316 699558 505322 699610
rect 505322 699558 505334 699610
rect 505334 699558 505372 699610
rect 504836 699556 504892 699558
rect 504916 699556 504972 699558
rect 504996 699556 505052 699558
rect 505076 699556 505132 699558
rect 505156 699556 505212 699558
rect 505236 699556 505292 699558
rect 505316 699556 505372 699558
rect 540836 699610 540892 699612
rect 540916 699610 540972 699612
rect 540996 699610 541052 699612
rect 541076 699610 541132 699612
rect 541156 699610 541212 699612
rect 541236 699610 541292 699612
rect 541316 699610 541372 699612
rect 540836 699558 540874 699610
rect 540874 699558 540886 699610
rect 540886 699558 540892 699610
rect 540916 699558 540938 699610
rect 540938 699558 540950 699610
rect 540950 699558 540972 699610
rect 540996 699558 541002 699610
rect 541002 699558 541014 699610
rect 541014 699558 541052 699610
rect 541076 699558 541078 699610
rect 541078 699558 541130 699610
rect 541130 699558 541132 699610
rect 541156 699558 541194 699610
rect 541194 699558 541206 699610
rect 541206 699558 541212 699610
rect 541236 699558 541258 699610
rect 541258 699558 541270 699610
rect 541270 699558 541292 699610
rect 541316 699558 541322 699610
rect 541322 699558 541334 699610
rect 541334 699558 541372 699610
rect 540836 699556 540892 699558
rect 540916 699556 540972 699558
rect 540996 699556 541052 699558
rect 541076 699556 541132 699558
rect 541156 699556 541212 699558
rect 541236 699556 541292 699558
rect 541316 699556 541372 699558
rect 576836 699610 576892 699612
rect 576916 699610 576972 699612
rect 576996 699610 577052 699612
rect 577076 699610 577132 699612
rect 577156 699610 577212 699612
rect 577236 699610 577292 699612
rect 577316 699610 577372 699612
rect 576836 699558 576874 699610
rect 576874 699558 576886 699610
rect 576886 699558 576892 699610
rect 576916 699558 576938 699610
rect 576938 699558 576950 699610
rect 576950 699558 576972 699610
rect 576996 699558 577002 699610
rect 577002 699558 577014 699610
rect 577014 699558 577052 699610
rect 577076 699558 577078 699610
rect 577078 699558 577130 699610
rect 577130 699558 577132 699610
rect 577156 699558 577194 699610
rect 577194 699558 577206 699610
rect 577206 699558 577212 699610
rect 577236 699558 577258 699610
rect 577258 699558 577270 699610
rect 577270 699558 577292 699610
rect 577316 699558 577322 699610
rect 577322 699558 577334 699610
rect 577334 699558 577372 699610
rect 576836 699556 576892 699558
rect 576916 699556 576972 699558
rect 576996 699556 577052 699558
rect 577076 699556 577132 699558
rect 577156 699556 577212 699558
rect 577236 699556 577292 699558
rect 577316 699556 577372 699558
rect 378836 699066 378892 699068
rect 378916 699066 378972 699068
rect 378996 699066 379052 699068
rect 379076 699066 379132 699068
rect 379156 699066 379212 699068
rect 379236 699066 379292 699068
rect 379316 699066 379372 699068
rect 378836 699014 378874 699066
rect 378874 699014 378886 699066
rect 378886 699014 378892 699066
rect 378916 699014 378938 699066
rect 378938 699014 378950 699066
rect 378950 699014 378972 699066
rect 378996 699014 379002 699066
rect 379002 699014 379014 699066
rect 379014 699014 379052 699066
rect 379076 699014 379078 699066
rect 379078 699014 379130 699066
rect 379130 699014 379132 699066
rect 379156 699014 379194 699066
rect 379194 699014 379206 699066
rect 379206 699014 379212 699066
rect 379236 699014 379258 699066
rect 379258 699014 379270 699066
rect 379270 699014 379292 699066
rect 379316 699014 379322 699066
rect 379322 699014 379334 699066
rect 379334 699014 379372 699066
rect 378836 699012 378892 699014
rect 378916 699012 378972 699014
rect 378996 699012 379052 699014
rect 379076 699012 379132 699014
rect 379156 699012 379212 699014
rect 379236 699012 379292 699014
rect 379316 699012 379372 699014
rect 396836 698522 396892 698524
rect 396916 698522 396972 698524
rect 396996 698522 397052 698524
rect 397076 698522 397132 698524
rect 397156 698522 397212 698524
rect 397236 698522 397292 698524
rect 397316 698522 397372 698524
rect 396836 698470 396874 698522
rect 396874 698470 396886 698522
rect 396886 698470 396892 698522
rect 396916 698470 396938 698522
rect 396938 698470 396950 698522
rect 396950 698470 396972 698522
rect 396996 698470 397002 698522
rect 397002 698470 397014 698522
rect 397014 698470 397052 698522
rect 397076 698470 397078 698522
rect 397078 698470 397130 698522
rect 397130 698470 397132 698522
rect 397156 698470 397194 698522
rect 397194 698470 397206 698522
rect 397206 698470 397212 698522
rect 397236 698470 397258 698522
rect 397258 698470 397270 698522
rect 397270 698470 397292 698522
rect 397316 698470 397322 698522
rect 397322 698470 397334 698522
rect 397334 698470 397372 698522
rect 396836 698468 396892 698470
rect 396916 698468 396972 698470
rect 396996 698468 397052 698470
rect 397076 698468 397132 698470
rect 397156 698468 397212 698470
rect 397236 698468 397292 698470
rect 397316 698468 397372 698470
rect 414836 699066 414892 699068
rect 414916 699066 414972 699068
rect 414996 699066 415052 699068
rect 415076 699066 415132 699068
rect 415156 699066 415212 699068
rect 415236 699066 415292 699068
rect 415316 699066 415372 699068
rect 414836 699014 414874 699066
rect 414874 699014 414886 699066
rect 414886 699014 414892 699066
rect 414916 699014 414938 699066
rect 414938 699014 414950 699066
rect 414950 699014 414972 699066
rect 414996 699014 415002 699066
rect 415002 699014 415014 699066
rect 415014 699014 415052 699066
rect 415076 699014 415078 699066
rect 415078 699014 415130 699066
rect 415130 699014 415132 699066
rect 415156 699014 415194 699066
rect 415194 699014 415206 699066
rect 415206 699014 415212 699066
rect 415236 699014 415258 699066
rect 415258 699014 415270 699066
rect 415270 699014 415292 699066
rect 415316 699014 415322 699066
rect 415322 699014 415334 699066
rect 415334 699014 415372 699066
rect 414836 699012 414892 699014
rect 414916 699012 414972 699014
rect 414996 699012 415052 699014
rect 415076 699012 415132 699014
rect 415156 699012 415212 699014
rect 415236 699012 415292 699014
rect 415316 699012 415372 699014
rect 530950 699216 531006 699272
rect 432836 698522 432892 698524
rect 432916 698522 432972 698524
rect 432996 698522 433052 698524
rect 433076 698522 433132 698524
rect 433156 698522 433212 698524
rect 433236 698522 433292 698524
rect 433316 698522 433372 698524
rect 432836 698470 432874 698522
rect 432874 698470 432886 698522
rect 432886 698470 432892 698522
rect 432916 698470 432938 698522
rect 432938 698470 432950 698522
rect 432950 698470 432972 698522
rect 432996 698470 433002 698522
rect 433002 698470 433014 698522
rect 433014 698470 433052 698522
rect 433076 698470 433078 698522
rect 433078 698470 433130 698522
rect 433130 698470 433132 698522
rect 433156 698470 433194 698522
rect 433194 698470 433206 698522
rect 433206 698470 433212 698522
rect 433236 698470 433258 698522
rect 433258 698470 433270 698522
rect 433270 698470 433292 698522
rect 433316 698470 433322 698522
rect 433322 698470 433334 698522
rect 433334 698470 433372 698522
rect 432836 698468 432892 698470
rect 432916 698468 432972 698470
rect 432996 698468 433052 698470
rect 433076 698468 433132 698470
rect 433156 698468 433212 698470
rect 433236 698468 433292 698470
rect 433316 698468 433372 698470
rect 450836 699066 450892 699068
rect 450916 699066 450972 699068
rect 450996 699066 451052 699068
rect 451076 699066 451132 699068
rect 451156 699066 451212 699068
rect 451236 699066 451292 699068
rect 451316 699066 451372 699068
rect 450836 699014 450874 699066
rect 450874 699014 450886 699066
rect 450886 699014 450892 699066
rect 450916 699014 450938 699066
rect 450938 699014 450950 699066
rect 450950 699014 450972 699066
rect 450996 699014 451002 699066
rect 451002 699014 451014 699066
rect 451014 699014 451052 699066
rect 451076 699014 451078 699066
rect 451078 699014 451130 699066
rect 451130 699014 451132 699066
rect 451156 699014 451194 699066
rect 451194 699014 451206 699066
rect 451206 699014 451212 699066
rect 451236 699014 451258 699066
rect 451258 699014 451270 699066
rect 451270 699014 451292 699066
rect 451316 699014 451322 699066
rect 451322 699014 451334 699066
rect 451334 699014 451372 699066
rect 450836 699012 450892 699014
rect 450916 699012 450972 699014
rect 450996 699012 451052 699014
rect 451076 699012 451132 699014
rect 451156 699012 451212 699014
rect 451236 699012 451292 699014
rect 451316 699012 451372 699014
rect 486836 699066 486892 699068
rect 486916 699066 486972 699068
rect 486996 699066 487052 699068
rect 487076 699066 487132 699068
rect 487156 699066 487212 699068
rect 487236 699066 487292 699068
rect 487316 699066 487372 699068
rect 486836 699014 486874 699066
rect 486874 699014 486886 699066
rect 486886 699014 486892 699066
rect 486916 699014 486938 699066
rect 486938 699014 486950 699066
rect 486950 699014 486972 699066
rect 486996 699014 487002 699066
rect 487002 699014 487014 699066
rect 487014 699014 487052 699066
rect 487076 699014 487078 699066
rect 487078 699014 487130 699066
rect 487130 699014 487132 699066
rect 487156 699014 487194 699066
rect 487194 699014 487206 699066
rect 487206 699014 487212 699066
rect 487236 699014 487258 699066
rect 487258 699014 487270 699066
rect 487270 699014 487292 699066
rect 487316 699014 487322 699066
rect 487322 699014 487334 699066
rect 487334 699014 487372 699066
rect 486836 699012 486892 699014
rect 486916 699012 486972 699014
rect 486996 699012 487052 699014
rect 487076 699012 487132 699014
rect 487156 699012 487212 699014
rect 487236 699012 487292 699014
rect 487316 699012 487372 699014
rect 522836 699066 522892 699068
rect 522916 699066 522972 699068
rect 522996 699066 523052 699068
rect 523076 699066 523132 699068
rect 523156 699066 523212 699068
rect 523236 699066 523292 699068
rect 523316 699066 523372 699068
rect 522836 699014 522874 699066
rect 522874 699014 522886 699066
rect 522886 699014 522892 699066
rect 522916 699014 522938 699066
rect 522938 699014 522950 699066
rect 522950 699014 522972 699066
rect 522996 699014 523002 699066
rect 523002 699014 523014 699066
rect 523014 699014 523052 699066
rect 523076 699014 523078 699066
rect 523078 699014 523130 699066
rect 523130 699014 523132 699066
rect 523156 699014 523194 699066
rect 523194 699014 523206 699066
rect 523206 699014 523212 699066
rect 523236 699014 523258 699066
rect 523258 699014 523270 699066
rect 523270 699014 523292 699066
rect 523316 699014 523322 699066
rect 523322 699014 523334 699066
rect 523334 699014 523372 699066
rect 522836 699012 522892 699014
rect 522916 699012 522972 699014
rect 522996 699012 523052 699014
rect 523076 699012 523132 699014
rect 523156 699012 523212 699014
rect 523236 699012 523292 699014
rect 523316 699012 523372 699014
rect 526258 698808 526314 698864
rect 468836 698522 468892 698524
rect 468916 698522 468972 698524
rect 468996 698522 469052 698524
rect 469076 698522 469132 698524
rect 469156 698522 469212 698524
rect 469236 698522 469292 698524
rect 469316 698522 469372 698524
rect 468836 698470 468874 698522
rect 468874 698470 468886 698522
rect 468886 698470 468892 698522
rect 468916 698470 468938 698522
rect 468938 698470 468950 698522
rect 468950 698470 468972 698522
rect 468996 698470 469002 698522
rect 469002 698470 469014 698522
rect 469014 698470 469052 698522
rect 469076 698470 469078 698522
rect 469078 698470 469130 698522
rect 469130 698470 469132 698522
rect 469156 698470 469194 698522
rect 469194 698470 469206 698522
rect 469206 698470 469212 698522
rect 469236 698470 469258 698522
rect 469258 698470 469270 698522
rect 469270 698470 469292 698522
rect 469316 698470 469322 698522
rect 469322 698470 469334 698522
rect 469334 698470 469372 698522
rect 468836 698468 468892 698470
rect 468916 698468 468972 698470
rect 468996 698468 469052 698470
rect 469076 698468 469132 698470
rect 469156 698468 469212 698470
rect 469236 698468 469292 698470
rect 469316 698468 469372 698470
rect 516782 698672 516838 698728
rect 504836 698522 504892 698524
rect 504916 698522 504972 698524
rect 504996 698522 505052 698524
rect 505076 698522 505132 698524
rect 505156 698522 505212 698524
rect 505236 698522 505292 698524
rect 505316 698522 505372 698524
rect 504836 698470 504874 698522
rect 504874 698470 504886 698522
rect 504886 698470 504892 698522
rect 504916 698470 504938 698522
rect 504938 698470 504950 698522
rect 504950 698470 504972 698522
rect 504996 698470 505002 698522
rect 505002 698470 505014 698522
rect 505014 698470 505052 698522
rect 505076 698470 505078 698522
rect 505078 698470 505130 698522
rect 505130 698470 505132 698522
rect 505156 698470 505194 698522
rect 505194 698470 505206 698522
rect 505206 698470 505212 698522
rect 505236 698470 505258 698522
rect 505258 698470 505270 698522
rect 505270 698470 505292 698522
rect 505316 698470 505322 698522
rect 505322 698470 505334 698522
rect 505334 698470 505372 698522
rect 504836 698468 504892 698470
rect 504916 698468 504972 698470
rect 504996 698468 505052 698470
rect 505076 698468 505132 698470
rect 505156 698468 505212 698470
rect 505236 698468 505292 698470
rect 505316 698468 505372 698470
rect 558836 699066 558892 699068
rect 558916 699066 558972 699068
rect 558996 699066 559052 699068
rect 559076 699066 559132 699068
rect 559156 699066 559212 699068
rect 559236 699066 559292 699068
rect 559316 699066 559372 699068
rect 558836 699014 558874 699066
rect 558874 699014 558886 699066
rect 558886 699014 558892 699066
rect 558916 699014 558938 699066
rect 558938 699014 558950 699066
rect 558950 699014 558972 699066
rect 558996 699014 559002 699066
rect 559002 699014 559014 699066
rect 559014 699014 559052 699066
rect 559076 699014 559078 699066
rect 559078 699014 559130 699066
rect 559130 699014 559132 699066
rect 559156 699014 559194 699066
rect 559194 699014 559206 699066
rect 559206 699014 559212 699066
rect 559236 699014 559258 699066
rect 559258 699014 559270 699066
rect 559270 699014 559292 699066
rect 559316 699014 559322 699066
rect 559322 699014 559334 699066
rect 559334 699014 559372 699066
rect 558836 699012 558892 699014
rect 558916 699012 558972 699014
rect 558996 699012 559052 699014
rect 559076 699012 559132 699014
rect 559156 699012 559212 699014
rect 559236 699012 559292 699014
rect 559316 699012 559372 699014
rect 540836 698522 540892 698524
rect 540916 698522 540972 698524
rect 540996 698522 541052 698524
rect 541076 698522 541132 698524
rect 541156 698522 541212 698524
rect 541236 698522 541292 698524
rect 541316 698522 541372 698524
rect 540836 698470 540874 698522
rect 540874 698470 540886 698522
rect 540886 698470 540892 698522
rect 540916 698470 540938 698522
rect 540938 698470 540950 698522
rect 540950 698470 540972 698522
rect 540996 698470 541002 698522
rect 541002 698470 541014 698522
rect 541014 698470 541052 698522
rect 541076 698470 541078 698522
rect 541078 698470 541130 698522
rect 541130 698470 541132 698522
rect 541156 698470 541194 698522
rect 541194 698470 541206 698522
rect 541206 698470 541212 698522
rect 541236 698470 541258 698522
rect 541258 698470 541270 698522
rect 541270 698470 541292 698522
rect 541316 698470 541322 698522
rect 541322 698470 541334 698522
rect 541334 698470 541372 698522
rect 540836 698468 540892 698470
rect 540916 698468 540972 698470
rect 540996 698468 541052 698470
rect 541076 698468 541132 698470
rect 541156 698468 541212 698470
rect 541236 698468 541292 698470
rect 541316 698468 541372 698470
rect 540426 697040 540482 697096
rect 509514 695816 509570 695872
rect 518070 695816 518126 695872
rect 545026 695680 545082 695736
rect 509514 695544 509570 695600
rect 518070 695544 518126 695600
rect 521382 695272 521438 695328
rect 569866 694048 569922 694104
rect 569866 693640 569922 693696
rect 574558 674872 574614 674928
rect 574742 696904 574798 696960
rect 574650 627952 574706 628008
rect 574834 694184 574890 694240
rect 576122 695544 576178 695600
rect 575478 674872 575534 674928
rect 575478 627952 575534 628008
rect 576836 698522 576892 698524
rect 576916 698522 576972 698524
rect 576996 698522 577052 698524
rect 577076 698522 577132 698524
rect 577156 698522 577212 698524
rect 577236 698522 577292 698524
rect 577316 698522 577372 698524
rect 576836 698470 576874 698522
rect 576874 698470 576886 698522
rect 576886 698470 576892 698522
rect 576916 698470 576938 698522
rect 576938 698470 576950 698522
rect 576950 698470 576972 698522
rect 576996 698470 577002 698522
rect 577002 698470 577014 698522
rect 577014 698470 577052 698522
rect 577076 698470 577078 698522
rect 577078 698470 577130 698522
rect 577130 698470 577132 698522
rect 577156 698470 577194 698522
rect 577194 698470 577206 698522
rect 577206 698470 577212 698522
rect 577236 698470 577258 698522
rect 577258 698470 577270 698522
rect 577270 698470 577292 698522
rect 577316 698470 577322 698522
rect 577322 698470 577334 698522
rect 577334 698470 577372 698522
rect 576836 698468 576892 698470
rect 576916 698468 576972 698470
rect 576996 698468 577052 698470
rect 577076 698468 577132 698470
rect 577156 698468 577212 698470
rect 577236 698468 577292 698470
rect 577316 698468 577372 698470
rect 579618 698028 579620 698048
rect 579620 698028 579672 698048
rect 579672 698028 579674 698048
rect 579618 697992 579674 698028
rect 579342 694048 579398 694104
rect 579802 674600 579858 674656
rect 579618 651072 579674 651128
rect 579526 639376 579582 639432
rect 579802 627680 579858 627736
rect 579618 604152 579674 604208
rect 579434 592456 579490 592512
rect 580170 580760 580226 580816
rect 579618 557232 579674 557288
rect 579342 545536 579398 545592
rect 579710 533840 579766 533896
rect 580170 510312 580226 510368
rect 580170 498616 580226 498672
rect 579986 486784 580042 486840
rect 579618 463392 579674 463448
rect 579250 451696 579306 451752
rect 579986 439864 580042 439920
rect 580170 416472 580226 416528
rect 579158 404776 579214 404832
rect 579066 392944 579122 393000
rect 579986 346024 580042 346080
rect 578974 322632 579030 322688
rect 579618 299104 579674 299160
rect 580170 263880 580226 263936
rect 580170 252184 580226 252240
rect 578882 216960 578938 217016
rect 580170 205264 580226 205320
rect 580170 181872 580226 181928
rect 579618 170040 579674 170096
rect 579618 111424 579674 111480
rect 580354 693776 580410 693832
rect 580538 693912 580594 693968
rect 580906 686296 580962 686352
rect 580814 369552 580870 369608
rect 580814 357856 580870 357912
rect 580814 310800 580870 310856
rect 580722 275712 580778 275768
rect 580630 228792 580686 228848
rect 580630 158344 580686 158400
rect 580538 134816 580594 134872
rect 580446 123120 580502 123176
rect 580354 87896 580410 87952
rect 580262 76200 580318 76256
rect 579802 64504 579858 64560
rect 580170 40976 580226 41032
rect 580170 29280 580226 29336
rect 580170 17584 580226 17640
rect 3146 7148 3148 7168
rect 3148 7148 3200 7168
rect 3200 7148 3202 7168
rect 3146 7112 3202 7148
rect 18836 6010 18892 6012
rect 18916 6010 18972 6012
rect 18996 6010 19052 6012
rect 19076 6010 19132 6012
rect 19156 6010 19212 6012
rect 19236 6010 19292 6012
rect 19316 6010 19372 6012
rect 18836 5958 18874 6010
rect 18874 5958 18886 6010
rect 18886 5958 18892 6010
rect 18916 5958 18938 6010
rect 18938 5958 18950 6010
rect 18950 5958 18972 6010
rect 18996 5958 19002 6010
rect 19002 5958 19014 6010
rect 19014 5958 19052 6010
rect 19076 5958 19078 6010
rect 19078 5958 19130 6010
rect 19130 5958 19132 6010
rect 19156 5958 19194 6010
rect 19194 5958 19206 6010
rect 19206 5958 19212 6010
rect 19236 5958 19258 6010
rect 19258 5958 19270 6010
rect 19270 5958 19292 6010
rect 19316 5958 19322 6010
rect 19322 5958 19334 6010
rect 19334 5958 19372 6010
rect 18836 5956 18892 5958
rect 18916 5956 18972 5958
rect 18996 5956 19052 5958
rect 19076 5956 19132 5958
rect 19156 5956 19212 5958
rect 19236 5956 19292 5958
rect 19316 5956 19372 5958
rect 18836 4922 18892 4924
rect 18916 4922 18972 4924
rect 18996 4922 19052 4924
rect 19076 4922 19132 4924
rect 19156 4922 19212 4924
rect 19236 4922 19292 4924
rect 19316 4922 19372 4924
rect 18836 4870 18874 4922
rect 18874 4870 18886 4922
rect 18886 4870 18892 4922
rect 18916 4870 18938 4922
rect 18938 4870 18950 4922
rect 18950 4870 18972 4922
rect 18996 4870 19002 4922
rect 19002 4870 19014 4922
rect 19014 4870 19052 4922
rect 19076 4870 19078 4922
rect 19078 4870 19130 4922
rect 19130 4870 19132 4922
rect 19156 4870 19194 4922
rect 19194 4870 19206 4922
rect 19206 4870 19212 4922
rect 19236 4870 19258 4922
rect 19258 4870 19270 4922
rect 19270 4870 19292 4922
rect 19316 4870 19322 4922
rect 19322 4870 19334 4922
rect 19334 4870 19372 4922
rect 18836 4868 18892 4870
rect 18916 4868 18972 4870
rect 18996 4868 19052 4870
rect 19076 4868 19132 4870
rect 19156 4868 19212 4870
rect 19236 4868 19292 4870
rect 19316 4868 19372 4870
rect 18836 3834 18892 3836
rect 18916 3834 18972 3836
rect 18996 3834 19052 3836
rect 19076 3834 19132 3836
rect 19156 3834 19212 3836
rect 19236 3834 19292 3836
rect 19316 3834 19372 3836
rect 18836 3782 18874 3834
rect 18874 3782 18886 3834
rect 18886 3782 18892 3834
rect 18916 3782 18938 3834
rect 18938 3782 18950 3834
rect 18950 3782 18972 3834
rect 18996 3782 19002 3834
rect 19002 3782 19014 3834
rect 19014 3782 19052 3834
rect 19076 3782 19078 3834
rect 19078 3782 19130 3834
rect 19130 3782 19132 3834
rect 19156 3782 19194 3834
rect 19194 3782 19206 3834
rect 19206 3782 19212 3834
rect 19236 3782 19258 3834
rect 19258 3782 19270 3834
rect 19270 3782 19292 3834
rect 19316 3782 19322 3834
rect 19322 3782 19334 3834
rect 19334 3782 19372 3834
rect 18836 3780 18892 3782
rect 18916 3780 18972 3782
rect 18996 3780 19052 3782
rect 19076 3780 19132 3782
rect 19156 3780 19212 3782
rect 19236 3780 19292 3782
rect 19316 3780 19372 3782
rect 18836 2746 18892 2748
rect 18916 2746 18972 2748
rect 18996 2746 19052 2748
rect 19076 2746 19132 2748
rect 19156 2746 19212 2748
rect 19236 2746 19292 2748
rect 19316 2746 19372 2748
rect 18836 2694 18874 2746
rect 18874 2694 18886 2746
rect 18886 2694 18892 2746
rect 18916 2694 18938 2746
rect 18938 2694 18950 2746
rect 18950 2694 18972 2746
rect 18996 2694 19002 2746
rect 19002 2694 19014 2746
rect 19014 2694 19052 2746
rect 19076 2694 19078 2746
rect 19078 2694 19130 2746
rect 19130 2694 19132 2746
rect 19156 2694 19194 2746
rect 19194 2694 19206 2746
rect 19206 2694 19212 2746
rect 19236 2694 19258 2746
rect 19258 2694 19270 2746
rect 19270 2694 19292 2746
rect 19316 2694 19322 2746
rect 19322 2694 19334 2746
rect 19334 2694 19372 2746
rect 18836 2692 18892 2694
rect 18916 2692 18972 2694
rect 18996 2692 19052 2694
rect 19076 2692 19132 2694
rect 19156 2692 19212 2694
rect 19236 2692 19292 2694
rect 19316 2692 19372 2694
rect 36836 5466 36892 5468
rect 36916 5466 36972 5468
rect 36996 5466 37052 5468
rect 37076 5466 37132 5468
rect 37156 5466 37212 5468
rect 37236 5466 37292 5468
rect 37316 5466 37372 5468
rect 36836 5414 36874 5466
rect 36874 5414 36886 5466
rect 36886 5414 36892 5466
rect 36916 5414 36938 5466
rect 36938 5414 36950 5466
rect 36950 5414 36972 5466
rect 36996 5414 37002 5466
rect 37002 5414 37014 5466
rect 37014 5414 37052 5466
rect 37076 5414 37078 5466
rect 37078 5414 37130 5466
rect 37130 5414 37132 5466
rect 37156 5414 37194 5466
rect 37194 5414 37206 5466
rect 37206 5414 37212 5466
rect 37236 5414 37258 5466
rect 37258 5414 37270 5466
rect 37270 5414 37292 5466
rect 37316 5414 37322 5466
rect 37322 5414 37334 5466
rect 37334 5414 37372 5466
rect 36836 5412 36892 5414
rect 36916 5412 36972 5414
rect 36996 5412 37052 5414
rect 37076 5412 37132 5414
rect 37156 5412 37212 5414
rect 37236 5412 37292 5414
rect 37316 5412 37372 5414
rect 36836 4378 36892 4380
rect 36916 4378 36972 4380
rect 36996 4378 37052 4380
rect 37076 4378 37132 4380
rect 37156 4378 37212 4380
rect 37236 4378 37292 4380
rect 37316 4378 37372 4380
rect 36836 4326 36874 4378
rect 36874 4326 36886 4378
rect 36886 4326 36892 4378
rect 36916 4326 36938 4378
rect 36938 4326 36950 4378
rect 36950 4326 36972 4378
rect 36996 4326 37002 4378
rect 37002 4326 37014 4378
rect 37014 4326 37052 4378
rect 37076 4326 37078 4378
rect 37078 4326 37130 4378
rect 37130 4326 37132 4378
rect 37156 4326 37194 4378
rect 37194 4326 37206 4378
rect 37206 4326 37212 4378
rect 37236 4326 37258 4378
rect 37258 4326 37270 4378
rect 37270 4326 37292 4378
rect 37316 4326 37322 4378
rect 37322 4326 37334 4378
rect 37334 4326 37372 4378
rect 36836 4324 36892 4326
rect 36916 4324 36972 4326
rect 36996 4324 37052 4326
rect 37076 4324 37132 4326
rect 37156 4324 37212 4326
rect 37236 4324 37292 4326
rect 37316 4324 37372 4326
rect 36836 3290 36892 3292
rect 36916 3290 36972 3292
rect 36996 3290 37052 3292
rect 37076 3290 37132 3292
rect 37156 3290 37212 3292
rect 37236 3290 37292 3292
rect 37316 3290 37372 3292
rect 36836 3238 36874 3290
rect 36874 3238 36886 3290
rect 36886 3238 36892 3290
rect 36916 3238 36938 3290
rect 36938 3238 36950 3290
rect 36950 3238 36972 3290
rect 36996 3238 37002 3290
rect 37002 3238 37014 3290
rect 37014 3238 37052 3290
rect 37076 3238 37078 3290
rect 37078 3238 37130 3290
rect 37130 3238 37132 3290
rect 37156 3238 37194 3290
rect 37194 3238 37206 3290
rect 37206 3238 37212 3290
rect 37236 3238 37258 3290
rect 37258 3238 37270 3290
rect 37270 3238 37292 3290
rect 37316 3238 37322 3290
rect 37322 3238 37334 3290
rect 37334 3238 37372 3290
rect 36836 3236 36892 3238
rect 36916 3236 36972 3238
rect 36996 3236 37052 3238
rect 37076 3236 37132 3238
rect 37156 3236 37212 3238
rect 37236 3236 37292 3238
rect 37316 3236 37372 3238
rect 36836 2202 36892 2204
rect 36916 2202 36972 2204
rect 36996 2202 37052 2204
rect 37076 2202 37132 2204
rect 37156 2202 37212 2204
rect 37236 2202 37292 2204
rect 37316 2202 37372 2204
rect 36836 2150 36874 2202
rect 36874 2150 36886 2202
rect 36886 2150 36892 2202
rect 36916 2150 36938 2202
rect 36938 2150 36950 2202
rect 36950 2150 36972 2202
rect 36996 2150 37002 2202
rect 37002 2150 37014 2202
rect 37014 2150 37052 2202
rect 37076 2150 37078 2202
rect 37078 2150 37130 2202
rect 37130 2150 37132 2202
rect 37156 2150 37194 2202
rect 37194 2150 37206 2202
rect 37206 2150 37212 2202
rect 37236 2150 37258 2202
rect 37258 2150 37270 2202
rect 37270 2150 37292 2202
rect 37316 2150 37322 2202
rect 37322 2150 37334 2202
rect 37334 2150 37372 2202
rect 36836 2148 36892 2150
rect 36916 2148 36972 2150
rect 36996 2148 37052 2150
rect 37076 2148 37132 2150
rect 37156 2148 37212 2150
rect 37236 2148 37292 2150
rect 37316 2148 37372 2150
rect 54836 6010 54892 6012
rect 54916 6010 54972 6012
rect 54996 6010 55052 6012
rect 55076 6010 55132 6012
rect 55156 6010 55212 6012
rect 55236 6010 55292 6012
rect 55316 6010 55372 6012
rect 54836 5958 54874 6010
rect 54874 5958 54886 6010
rect 54886 5958 54892 6010
rect 54916 5958 54938 6010
rect 54938 5958 54950 6010
rect 54950 5958 54972 6010
rect 54996 5958 55002 6010
rect 55002 5958 55014 6010
rect 55014 5958 55052 6010
rect 55076 5958 55078 6010
rect 55078 5958 55130 6010
rect 55130 5958 55132 6010
rect 55156 5958 55194 6010
rect 55194 5958 55206 6010
rect 55206 5958 55212 6010
rect 55236 5958 55258 6010
rect 55258 5958 55270 6010
rect 55270 5958 55292 6010
rect 55316 5958 55322 6010
rect 55322 5958 55334 6010
rect 55334 5958 55372 6010
rect 54836 5956 54892 5958
rect 54916 5956 54972 5958
rect 54996 5956 55052 5958
rect 55076 5956 55132 5958
rect 55156 5956 55212 5958
rect 55236 5956 55292 5958
rect 55316 5956 55372 5958
rect 54836 4922 54892 4924
rect 54916 4922 54972 4924
rect 54996 4922 55052 4924
rect 55076 4922 55132 4924
rect 55156 4922 55212 4924
rect 55236 4922 55292 4924
rect 55316 4922 55372 4924
rect 54836 4870 54874 4922
rect 54874 4870 54886 4922
rect 54886 4870 54892 4922
rect 54916 4870 54938 4922
rect 54938 4870 54950 4922
rect 54950 4870 54972 4922
rect 54996 4870 55002 4922
rect 55002 4870 55014 4922
rect 55014 4870 55052 4922
rect 55076 4870 55078 4922
rect 55078 4870 55130 4922
rect 55130 4870 55132 4922
rect 55156 4870 55194 4922
rect 55194 4870 55206 4922
rect 55206 4870 55212 4922
rect 55236 4870 55258 4922
rect 55258 4870 55270 4922
rect 55270 4870 55292 4922
rect 55316 4870 55322 4922
rect 55322 4870 55334 4922
rect 55334 4870 55372 4922
rect 54836 4868 54892 4870
rect 54916 4868 54972 4870
rect 54996 4868 55052 4870
rect 55076 4868 55132 4870
rect 55156 4868 55212 4870
rect 55236 4868 55292 4870
rect 55316 4868 55372 4870
rect 54836 3834 54892 3836
rect 54916 3834 54972 3836
rect 54996 3834 55052 3836
rect 55076 3834 55132 3836
rect 55156 3834 55212 3836
rect 55236 3834 55292 3836
rect 55316 3834 55372 3836
rect 54836 3782 54874 3834
rect 54874 3782 54886 3834
rect 54886 3782 54892 3834
rect 54916 3782 54938 3834
rect 54938 3782 54950 3834
rect 54950 3782 54972 3834
rect 54996 3782 55002 3834
rect 55002 3782 55014 3834
rect 55014 3782 55052 3834
rect 55076 3782 55078 3834
rect 55078 3782 55130 3834
rect 55130 3782 55132 3834
rect 55156 3782 55194 3834
rect 55194 3782 55206 3834
rect 55206 3782 55212 3834
rect 55236 3782 55258 3834
rect 55258 3782 55270 3834
rect 55270 3782 55292 3834
rect 55316 3782 55322 3834
rect 55322 3782 55334 3834
rect 55334 3782 55372 3834
rect 54836 3780 54892 3782
rect 54916 3780 54972 3782
rect 54996 3780 55052 3782
rect 55076 3780 55132 3782
rect 55156 3780 55212 3782
rect 55236 3780 55292 3782
rect 55316 3780 55372 3782
rect 54836 2746 54892 2748
rect 54916 2746 54972 2748
rect 54996 2746 55052 2748
rect 55076 2746 55132 2748
rect 55156 2746 55212 2748
rect 55236 2746 55292 2748
rect 55316 2746 55372 2748
rect 54836 2694 54874 2746
rect 54874 2694 54886 2746
rect 54886 2694 54892 2746
rect 54916 2694 54938 2746
rect 54938 2694 54950 2746
rect 54950 2694 54972 2746
rect 54996 2694 55002 2746
rect 55002 2694 55014 2746
rect 55014 2694 55052 2746
rect 55076 2694 55078 2746
rect 55078 2694 55130 2746
rect 55130 2694 55132 2746
rect 55156 2694 55194 2746
rect 55194 2694 55206 2746
rect 55206 2694 55212 2746
rect 55236 2694 55258 2746
rect 55258 2694 55270 2746
rect 55270 2694 55292 2746
rect 55316 2694 55322 2746
rect 55322 2694 55334 2746
rect 55334 2694 55372 2746
rect 54836 2692 54892 2694
rect 54916 2692 54972 2694
rect 54996 2692 55052 2694
rect 55076 2692 55132 2694
rect 55156 2692 55212 2694
rect 55236 2692 55292 2694
rect 55316 2692 55372 2694
rect 72836 5466 72892 5468
rect 72916 5466 72972 5468
rect 72996 5466 73052 5468
rect 73076 5466 73132 5468
rect 73156 5466 73212 5468
rect 73236 5466 73292 5468
rect 73316 5466 73372 5468
rect 72836 5414 72874 5466
rect 72874 5414 72886 5466
rect 72886 5414 72892 5466
rect 72916 5414 72938 5466
rect 72938 5414 72950 5466
rect 72950 5414 72972 5466
rect 72996 5414 73002 5466
rect 73002 5414 73014 5466
rect 73014 5414 73052 5466
rect 73076 5414 73078 5466
rect 73078 5414 73130 5466
rect 73130 5414 73132 5466
rect 73156 5414 73194 5466
rect 73194 5414 73206 5466
rect 73206 5414 73212 5466
rect 73236 5414 73258 5466
rect 73258 5414 73270 5466
rect 73270 5414 73292 5466
rect 73316 5414 73322 5466
rect 73322 5414 73334 5466
rect 73334 5414 73372 5466
rect 72836 5412 72892 5414
rect 72916 5412 72972 5414
rect 72996 5412 73052 5414
rect 73076 5412 73132 5414
rect 73156 5412 73212 5414
rect 73236 5412 73292 5414
rect 73316 5412 73372 5414
rect 72836 4378 72892 4380
rect 72916 4378 72972 4380
rect 72996 4378 73052 4380
rect 73076 4378 73132 4380
rect 73156 4378 73212 4380
rect 73236 4378 73292 4380
rect 73316 4378 73372 4380
rect 72836 4326 72874 4378
rect 72874 4326 72886 4378
rect 72886 4326 72892 4378
rect 72916 4326 72938 4378
rect 72938 4326 72950 4378
rect 72950 4326 72972 4378
rect 72996 4326 73002 4378
rect 73002 4326 73014 4378
rect 73014 4326 73052 4378
rect 73076 4326 73078 4378
rect 73078 4326 73130 4378
rect 73130 4326 73132 4378
rect 73156 4326 73194 4378
rect 73194 4326 73206 4378
rect 73206 4326 73212 4378
rect 73236 4326 73258 4378
rect 73258 4326 73270 4378
rect 73270 4326 73292 4378
rect 73316 4326 73322 4378
rect 73322 4326 73334 4378
rect 73334 4326 73372 4378
rect 72836 4324 72892 4326
rect 72916 4324 72972 4326
rect 72996 4324 73052 4326
rect 73076 4324 73132 4326
rect 73156 4324 73212 4326
rect 73236 4324 73292 4326
rect 73316 4324 73372 4326
rect 72836 3290 72892 3292
rect 72916 3290 72972 3292
rect 72996 3290 73052 3292
rect 73076 3290 73132 3292
rect 73156 3290 73212 3292
rect 73236 3290 73292 3292
rect 73316 3290 73372 3292
rect 72836 3238 72874 3290
rect 72874 3238 72886 3290
rect 72886 3238 72892 3290
rect 72916 3238 72938 3290
rect 72938 3238 72950 3290
rect 72950 3238 72972 3290
rect 72996 3238 73002 3290
rect 73002 3238 73014 3290
rect 73014 3238 73052 3290
rect 73076 3238 73078 3290
rect 73078 3238 73130 3290
rect 73130 3238 73132 3290
rect 73156 3238 73194 3290
rect 73194 3238 73206 3290
rect 73206 3238 73212 3290
rect 73236 3238 73258 3290
rect 73258 3238 73270 3290
rect 73270 3238 73292 3290
rect 73316 3238 73322 3290
rect 73322 3238 73334 3290
rect 73334 3238 73372 3290
rect 72836 3236 72892 3238
rect 72916 3236 72972 3238
rect 72996 3236 73052 3238
rect 73076 3236 73132 3238
rect 73156 3236 73212 3238
rect 73236 3236 73292 3238
rect 73316 3236 73372 3238
rect 72836 2202 72892 2204
rect 72916 2202 72972 2204
rect 72996 2202 73052 2204
rect 73076 2202 73132 2204
rect 73156 2202 73212 2204
rect 73236 2202 73292 2204
rect 73316 2202 73372 2204
rect 72836 2150 72874 2202
rect 72874 2150 72886 2202
rect 72886 2150 72892 2202
rect 72916 2150 72938 2202
rect 72938 2150 72950 2202
rect 72950 2150 72972 2202
rect 72996 2150 73002 2202
rect 73002 2150 73014 2202
rect 73014 2150 73052 2202
rect 73076 2150 73078 2202
rect 73078 2150 73130 2202
rect 73130 2150 73132 2202
rect 73156 2150 73194 2202
rect 73194 2150 73206 2202
rect 73206 2150 73212 2202
rect 73236 2150 73258 2202
rect 73258 2150 73270 2202
rect 73270 2150 73292 2202
rect 73316 2150 73322 2202
rect 73322 2150 73334 2202
rect 73334 2150 73372 2202
rect 72836 2148 72892 2150
rect 72916 2148 72972 2150
rect 72996 2148 73052 2150
rect 73076 2148 73132 2150
rect 73156 2148 73212 2150
rect 73236 2148 73292 2150
rect 73316 2148 73372 2150
rect 90836 6010 90892 6012
rect 90916 6010 90972 6012
rect 90996 6010 91052 6012
rect 91076 6010 91132 6012
rect 91156 6010 91212 6012
rect 91236 6010 91292 6012
rect 91316 6010 91372 6012
rect 90836 5958 90874 6010
rect 90874 5958 90886 6010
rect 90886 5958 90892 6010
rect 90916 5958 90938 6010
rect 90938 5958 90950 6010
rect 90950 5958 90972 6010
rect 90996 5958 91002 6010
rect 91002 5958 91014 6010
rect 91014 5958 91052 6010
rect 91076 5958 91078 6010
rect 91078 5958 91130 6010
rect 91130 5958 91132 6010
rect 91156 5958 91194 6010
rect 91194 5958 91206 6010
rect 91206 5958 91212 6010
rect 91236 5958 91258 6010
rect 91258 5958 91270 6010
rect 91270 5958 91292 6010
rect 91316 5958 91322 6010
rect 91322 5958 91334 6010
rect 91334 5958 91372 6010
rect 90836 5956 90892 5958
rect 90916 5956 90972 5958
rect 90996 5956 91052 5958
rect 91076 5956 91132 5958
rect 91156 5956 91212 5958
rect 91236 5956 91292 5958
rect 91316 5956 91372 5958
rect 90836 4922 90892 4924
rect 90916 4922 90972 4924
rect 90996 4922 91052 4924
rect 91076 4922 91132 4924
rect 91156 4922 91212 4924
rect 91236 4922 91292 4924
rect 91316 4922 91372 4924
rect 90836 4870 90874 4922
rect 90874 4870 90886 4922
rect 90886 4870 90892 4922
rect 90916 4870 90938 4922
rect 90938 4870 90950 4922
rect 90950 4870 90972 4922
rect 90996 4870 91002 4922
rect 91002 4870 91014 4922
rect 91014 4870 91052 4922
rect 91076 4870 91078 4922
rect 91078 4870 91130 4922
rect 91130 4870 91132 4922
rect 91156 4870 91194 4922
rect 91194 4870 91206 4922
rect 91206 4870 91212 4922
rect 91236 4870 91258 4922
rect 91258 4870 91270 4922
rect 91270 4870 91292 4922
rect 91316 4870 91322 4922
rect 91322 4870 91334 4922
rect 91334 4870 91372 4922
rect 90836 4868 90892 4870
rect 90916 4868 90972 4870
rect 90996 4868 91052 4870
rect 91076 4868 91132 4870
rect 91156 4868 91212 4870
rect 91236 4868 91292 4870
rect 91316 4868 91372 4870
rect 90836 3834 90892 3836
rect 90916 3834 90972 3836
rect 90996 3834 91052 3836
rect 91076 3834 91132 3836
rect 91156 3834 91212 3836
rect 91236 3834 91292 3836
rect 91316 3834 91372 3836
rect 90836 3782 90874 3834
rect 90874 3782 90886 3834
rect 90886 3782 90892 3834
rect 90916 3782 90938 3834
rect 90938 3782 90950 3834
rect 90950 3782 90972 3834
rect 90996 3782 91002 3834
rect 91002 3782 91014 3834
rect 91014 3782 91052 3834
rect 91076 3782 91078 3834
rect 91078 3782 91130 3834
rect 91130 3782 91132 3834
rect 91156 3782 91194 3834
rect 91194 3782 91206 3834
rect 91206 3782 91212 3834
rect 91236 3782 91258 3834
rect 91258 3782 91270 3834
rect 91270 3782 91292 3834
rect 91316 3782 91322 3834
rect 91322 3782 91334 3834
rect 91334 3782 91372 3834
rect 90836 3780 90892 3782
rect 90916 3780 90972 3782
rect 90996 3780 91052 3782
rect 91076 3780 91132 3782
rect 91156 3780 91212 3782
rect 91236 3780 91292 3782
rect 91316 3780 91372 3782
rect 90836 2746 90892 2748
rect 90916 2746 90972 2748
rect 90996 2746 91052 2748
rect 91076 2746 91132 2748
rect 91156 2746 91212 2748
rect 91236 2746 91292 2748
rect 91316 2746 91372 2748
rect 90836 2694 90874 2746
rect 90874 2694 90886 2746
rect 90886 2694 90892 2746
rect 90916 2694 90938 2746
rect 90938 2694 90950 2746
rect 90950 2694 90972 2746
rect 90996 2694 91002 2746
rect 91002 2694 91014 2746
rect 91014 2694 91052 2746
rect 91076 2694 91078 2746
rect 91078 2694 91130 2746
rect 91130 2694 91132 2746
rect 91156 2694 91194 2746
rect 91194 2694 91206 2746
rect 91206 2694 91212 2746
rect 91236 2694 91258 2746
rect 91258 2694 91270 2746
rect 91270 2694 91292 2746
rect 91316 2694 91322 2746
rect 91322 2694 91334 2746
rect 91334 2694 91372 2746
rect 90836 2692 90892 2694
rect 90916 2692 90972 2694
rect 90996 2692 91052 2694
rect 91076 2692 91132 2694
rect 91156 2692 91212 2694
rect 91236 2692 91292 2694
rect 91316 2692 91372 2694
rect 108836 5466 108892 5468
rect 108916 5466 108972 5468
rect 108996 5466 109052 5468
rect 109076 5466 109132 5468
rect 109156 5466 109212 5468
rect 109236 5466 109292 5468
rect 109316 5466 109372 5468
rect 108836 5414 108874 5466
rect 108874 5414 108886 5466
rect 108886 5414 108892 5466
rect 108916 5414 108938 5466
rect 108938 5414 108950 5466
rect 108950 5414 108972 5466
rect 108996 5414 109002 5466
rect 109002 5414 109014 5466
rect 109014 5414 109052 5466
rect 109076 5414 109078 5466
rect 109078 5414 109130 5466
rect 109130 5414 109132 5466
rect 109156 5414 109194 5466
rect 109194 5414 109206 5466
rect 109206 5414 109212 5466
rect 109236 5414 109258 5466
rect 109258 5414 109270 5466
rect 109270 5414 109292 5466
rect 109316 5414 109322 5466
rect 109322 5414 109334 5466
rect 109334 5414 109372 5466
rect 108836 5412 108892 5414
rect 108916 5412 108972 5414
rect 108996 5412 109052 5414
rect 109076 5412 109132 5414
rect 109156 5412 109212 5414
rect 109236 5412 109292 5414
rect 109316 5412 109372 5414
rect 108836 4378 108892 4380
rect 108916 4378 108972 4380
rect 108996 4378 109052 4380
rect 109076 4378 109132 4380
rect 109156 4378 109212 4380
rect 109236 4378 109292 4380
rect 109316 4378 109372 4380
rect 108836 4326 108874 4378
rect 108874 4326 108886 4378
rect 108886 4326 108892 4378
rect 108916 4326 108938 4378
rect 108938 4326 108950 4378
rect 108950 4326 108972 4378
rect 108996 4326 109002 4378
rect 109002 4326 109014 4378
rect 109014 4326 109052 4378
rect 109076 4326 109078 4378
rect 109078 4326 109130 4378
rect 109130 4326 109132 4378
rect 109156 4326 109194 4378
rect 109194 4326 109206 4378
rect 109206 4326 109212 4378
rect 109236 4326 109258 4378
rect 109258 4326 109270 4378
rect 109270 4326 109292 4378
rect 109316 4326 109322 4378
rect 109322 4326 109334 4378
rect 109334 4326 109372 4378
rect 108836 4324 108892 4326
rect 108916 4324 108972 4326
rect 108996 4324 109052 4326
rect 109076 4324 109132 4326
rect 109156 4324 109212 4326
rect 109236 4324 109292 4326
rect 109316 4324 109372 4326
rect 108836 3290 108892 3292
rect 108916 3290 108972 3292
rect 108996 3290 109052 3292
rect 109076 3290 109132 3292
rect 109156 3290 109212 3292
rect 109236 3290 109292 3292
rect 109316 3290 109372 3292
rect 108836 3238 108874 3290
rect 108874 3238 108886 3290
rect 108886 3238 108892 3290
rect 108916 3238 108938 3290
rect 108938 3238 108950 3290
rect 108950 3238 108972 3290
rect 108996 3238 109002 3290
rect 109002 3238 109014 3290
rect 109014 3238 109052 3290
rect 109076 3238 109078 3290
rect 109078 3238 109130 3290
rect 109130 3238 109132 3290
rect 109156 3238 109194 3290
rect 109194 3238 109206 3290
rect 109206 3238 109212 3290
rect 109236 3238 109258 3290
rect 109258 3238 109270 3290
rect 109270 3238 109292 3290
rect 109316 3238 109322 3290
rect 109322 3238 109334 3290
rect 109334 3238 109372 3290
rect 108836 3236 108892 3238
rect 108916 3236 108972 3238
rect 108996 3236 109052 3238
rect 109076 3236 109132 3238
rect 109156 3236 109212 3238
rect 109236 3236 109292 3238
rect 109316 3236 109372 3238
rect 108836 2202 108892 2204
rect 108916 2202 108972 2204
rect 108996 2202 109052 2204
rect 109076 2202 109132 2204
rect 109156 2202 109212 2204
rect 109236 2202 109292 2204
rect 109316 2202 109372 2204
rect 108836 2150 108874 2202
rect 108874 2150 108886 2202
rect 108886 2150 108892 2202
rect 108916 2150 108938 2202
rect 108938 2150 108950 2202
rect 108950 2150 108972 2202
rect 108996 2150 109002 2202
rect 109002 2150 109014 2202
rect 109014 2150 109052 2202
rect 109076 2150 109078 2202
rect 109078 2150 109130 2202
rect 109130 2150 109132 2202
rect 109156 2150 109194 2202
rect 109194 2150 109206 2202
rect 109206 2150 109212 2202
rect 109236 2150 109258 2202
rect 109258 2150 109270 2202
rect 109270 2150 109292 2202
rect 109316 2150 109322 2202
rect 109322 2150 109334 2202
rect 109334 2150 109372 2202
rect 108836 2148 108892 2150
rect 108916 2148 108972 2150
rect 108996 2148 109052 2150
rect 109076 2148 109132 2150
rect 109156 2148 109212 2150
rect 109236 2148 109292 2150
rect 109316 2148 109372 2150
rect 126836 6010 126892 6012
rect 126916 6010 126972 6012
rect 126996 6010 127052 6012
rect 127076 6010 127132 6012
rect 127156 6010 127212 6012
rect 127236 6010 127292 6012
rect 127316 6010 127372 6012
rect 126836 5958 126874 6010
rect 126874 5958 126886 6010
rect 126886 5958 126892 6010
rect 126916 5958 126938 6010
rect 126938 5958 126950 6010
rect 126950 5958 126972 6010
rect 126996 5958 127002 6010
rect 127002 5958 127014 6010
rect 127014 5958 127052 6010
rect 127076 5958 127078 6010
rect 127078 5958 127130 6010
rect 127130 5958 127132 6010
rect 127156 5958 127194 6010
rect 127194 5958 127206 6010
rect 127206 5958 127212 6010
rect 127236 5958 127258 6010
rect 127258 5958 127270 6010
rect 127270 5958 127292 6010
rect 127316 5958 127322 6010
rect 127322 5958 127334 6010
rect 127334 5958 127372 6010
rect 126836 5956 126892 5958
rect 126916 5956 126972 5958
rect 126996 5956 127052 5958
rect 127076 5956 127132 5958
rect 127156 5956 127212 5958
rect 127236 5956 127292 5958
rect 127316 5956 127372 5958
rect 126836 4922 126892 4924
rect 126916 4922 126972 4924
rect 126996 4922 127052 4924
rect 127076 4922 127132 4924
rect 127156 4922 127212 4924
rect 127236 4922 127292 4924
rect 127316 4922 127372 4924
rect 126836 4870 126874 4922
rect 126874 4870 126886 4922
rect 126886 4870 126892 4922
rect 126916 4870 126938 4922
rect 126938 4870 126950 4922
rect 126950 4870 126972 4922
rect 126996 4870 127002 4922
rect 127002 4870 127014 4922
rect 127014 4870 127052 4922
rect 127076 4870 127078 4922
rect 127078 4870 127130 4922
rect 127130 4870 127132 4922
rect 127156 4870 127194 4922
rect 127194 4870 127206 4922
rect 127206 4870 127212 4922
rect 127236 4870 127258 4922
rect 127258 4870 127270 4922
rect 127270 4870 127292 4922
rect 127316 4870 127322 4922
rect 127322 4870 127334 4922
rect 127334 4870 127372 4922
rect 126836 4868 126892 4870
rect 126916 4868 126972 4870
rect 126996 4868 127052 4870
rect 127076 4868 127132 4870
rect 127156 4868 127212 4870
rect 127236 4868 127292 4870
rect 127316 4868 127372 4870
rect 126836 3834 126892 3836
rect 126916 3834 126972 3836
rect 126996 3834 127052 3836
rect 127076 3834 127132 3836
rect 127156 3834 127212 3836
rect 127236 3834 127292 3836
rect 127316 3834 127372 3836
rect 126836 3782 126874 3834
rect 126874 3782 126886 3834
rect 126886 3782 126892 3834
rect 126916 3782 126938 3834
rect 126938 3782 126950 3834
rect 126950 3782 126972 3834
rect 126996 3782 127002 3834
rect 127002 3782 127014 3834
rect 127014 3782 127052 3834
rect 127076 3782 127078 3834
rect 127078 3782 127130 3834
rect 127130 3782 127132 3834
rect 127156 3782 127194 3834
rect 127194 3782 127206 3834
rect 127206 3782 127212 3834
rect 127236 3782 127258 3834
rect 127258 3782 127270 3834
rect 127270 3782 127292 3834
rect 127316 3782 127322 3834
rect 127322 3782 127334 3834
rect 127334 3782 127372 3834
rect 126836 3780 126892 3782
rect 126916 3780 126972 3782
rect 126996 3780 127052 3782
rect 127076 3780 127132 3782
rect 127156 3780 127212 3782
rect 127236 3780 127292 3782
rect 127316 3780 127372 3782
rect 126836 2746 126892 2748
rect 126916 2746 126972 2748
rect 126996 2746 127052 2748
rect 127076 2746 127132 2748
rect 127156 2746 127212 2748
rect 127236 2746 127292 2748
rect 127316 2746 127372 2748
rect 126836 2694 126874 2746
rect 126874 2694 126886 2746
rect 126886 2694 126892 2746
rect 126916 2694 126938 2746
rect 126938 2694 126950 2746
rect 126950 2694 126972 2746
rect 126996 2694 127002 2746
rect 127002 2694 127014 2746
rect 127014 2694 127052 2746
rect 127076 2694 127078 2746
rect 127078 2694 127130 2746
rect 127130 2694 127132 2746
rect 127156 2694 127194 2746
rect 127194 2694 127206 2746
rect 127206 2694 127212 2746
rect 127236 2694 127258 2746
rect 127258 2694 127270 2746
rect 127270 2694 127292 2746
rect 127316 2694 127322 2746
rect 127322 2694 127334 2746
rect 127334 2694 127372 2746
rect 126836 2692 126892 2694
rect 126916 2692 126972 2694
rect 126996 2692 127052 2694
rect 127076 2692 127132 2694
rect 127156 2692 127212 2694
rect 127236 2692 127292 2694
rect 127316 2692 127372 2694
rect 144836 5466 144892 5468
rect 144916 5466 144972 5468
rect 144996 5466 145052 5468
rect 145076 5466 145132 5468
rect 145156 5466 145212 5468
rect 145236 5466 145292 5468
rect 145316 5466 145372 5468
rect 144836 5414 144874 5466
rect 144874 5414 144886 5466
rect 144886 5414 144892 5466
rect 144916 5414 144938 5466
rect 144938 5414 144950 5466
rect 144950 5414 144972 5466
rect 144996 5414 145002 5466
rect 145002 5414 145014 5466
rect 145014 5414 145052 5466
rect 145076 5414 145078 5466
rect 145078 5414 145130 5466
rect 145130 5414 145132 5466
rect 145156 5414 145194 5466
rect 145194 5414 145206 5466
rect 145206 5414 145212 5466
rect 145236 5414 145258 5466
rect 145258 5414 145270 5466
rect 145270 5414 145292 5466
rect 145316 5414 145322 5466
rect 145322 5414 145334 5466
rect 145334 5414 145372 5466
rect 144836 5412 144892 5414
rect 144916 5412 144972 5414
rect 144996 5412 145052 5414
rect 145076 5412 145132 5414
rect 145156 5412 145212 5414
rect 145236 5412 145292 5414
rect 145316 5412 145372 5414
rect 144836 4378 144892 4380
rect 144916 4378 144972 4380
rect 144996 4378 145052 4380
rect 145076 4378 145132 4380
rect 145156 4378 145212 4380
rect 145236 4378 145292 4380
rect 145316 4378 145372 4380
rect 144836 4326 144874 4378
rect 144874 4326 144886 4378
rect 144886 4326 144892 4378
rect 144916 4326 144938 4378
rect 144938 4326 144950 4378
rect 144950 4326 144972 4378
rect 144996 4326 145002 4378
rect 145002 4326 145014 4378
rect 145014 4326 145052 4378
rect 145076 4326 145078 4378
rect 145078 4326 145130 4378
rect 145130 4326 145132 4378
rect 145156 4326 145194 4378
rect 145194 4326 145206 4378
rect 145206 4326 145212 4378
rect 145236 4326 145258 4378
rect 145258 4326 145270 4378
rect 145270 4326 145292 4378
rect 145316 4326 145322 4378
rect 145322 4326 145334 4378
rect 145334 4326 145372 4378
rect 144836 4324 144892 4326
rect 144916 4324 144972 4326
rect 144996 4324 145052 4326
rect 145076 4324 145132 4326
rect 145156 4324 145212 4326
rect 145236 4324 145292 4326
rect 145316 4324 145372 4326
rect 144836 3290 144892 3292
rect 144916 3290 144972 3292
rect 144996 3290 145052 3292
rect 145076 3290 145132 3292
rect 145156 3290 145212 3292
rect 145236 3290 145292 3292
rect 145316 3290 145372 3292
rect 144836 3238 144874 3290
rect 144874 3238 144886 3290
rect 144886 3238 144892 3290
rect 144916 3238 144938 3290
rect 144938 3238 144950 3290
rect 144950 3238 144972 3290
rect 144996 3238 145002 3290
rect 145002 3238 145014 3290
rect 145014 3238 145052 3290
rect 145076 3238 145078 3290
rect 145078 3238 145130 3290
rect 145130 3238 145132 3290
rect 145156 3238 145194 3290
rect 145194 3238 145206 3290
rect 145206 3238 145212 3290
rect 145236 3238 145258 3290
rect 145258 3238 145270 3290
rect 145270 3238 145292 3290
rect 145316 3238 145322 3290
rect 145322 3238 145334 3290
rect 145334 3238 145372 3290
rect 144836 3236 144892 3238
rect 144916 3236 144972 3238
rect 144996 3236 145052 3238
rect 145076 3236 145132 3238
rect 145156 3236 145212 3238
rect 145236 3236 145292 3238
rect 145316 3236 145372 3238
rect 144836 2202 144892 2204
rect 144916 2202 144972 2204
rect 144996 2202 145052 2204
rect 145076 2202 145132 2204
rect 145156 2202 145212 2204
rect 145236 2202 145292 2204
rect 145316 2202 145372 2204
rect 144836 2150 144874 2202
rect 144874 2150 144886 2202
rect 144886 2150 144892 2202
rect 144916 2150 144938 2202
rect 144938 2150 144950 2202
rect 144950 2150 144972 2202
rect 144996 2150 145002 2202
rect 145002 2150 145014 2202
rect 145014 2150 145052 2202
rect 145076 2150 145078 2202
rect 145078 2150 145130 2202
rect 145130 2150 145132 2202
rect 145156 2150 145194 2202
rect 145194 2150 145206 2202
rect 145206 2150 145212 2202
rect 145236 2150 145258 2202
rect 145258 2150 145270 2202
rect 145270 2150 145292 2202
rect 145316 2150 145322 2202
rect 145322 2150 145334 2202
rect 145334 2150 145372 2202
rect 144836 2148 144892 2150
rect 144916 2148 144972 2150
rect 144996 2148 145052 2150
rect 145076 2148 145132 2150
rect 145156 2148 145212 2150
rect 145236 2148 145292 2150
rect 145316 2148 145372 2150
rect 162836 6010 162892 6012
rect 162916 6010 162972 6012
rect 162996 6010 163052 6012
rect 163076 6010 163132 6012
rect 163156 6010 163212 6012
rect 163236 6010 163292 6012
rect 163316 6010 163372 6012
rect 162836 5958 162874 6010
rect 162874 5958 162886 6010
rect 162886 5958 162892 6010
rect 162916 5958 162938 6010
rect 162938 5958 162950 6010
rect 162950 5958 162972 6010
rect 162996 5958 163002 6010
rect 163002 5958 163014 6010
rect 163014 5958 163052 6010
rect 163076 5958 163078 6010
rect 163078 5958 163130 6010
rect 163130 5958 163132 6010
rect 163156 5958 163194 6010
rect 163194 5958 163206 6010
rect 163206 5958 163212 6010
rect 163236 5958 163258 6010
rect 163258 5958 163270 6010
rect 163270 5958 163292 6010
rect 163316 5958 163322 6010
rect 163322 5958 163334 6010
rect 163334 5958 163372 6010
rect 162836 5956 162892 5958
rect 162916 5956 162972 5958
rect 162996 5956 163052 5958
rect 163076 5956 163132 5958
rect 163156 5956 163212 5958
rect 163236 5956 163292 5958
rect 163316 5956 163372 5958
rect 162836 4922 162892 4924
rect 162916 4922 162972 4924
rect 162996 4922 163052 4924
rect 163076 4922 163132 4924
rect 163156 4922 163212 4924
rect 163236 4922 163292 4924
rect 163316 4922 163372 4924
rect 162836 4870 162874 4922
rect 162874 4870 162886 4922
rect 162886 4870 162892 4922
rect 162916 4870 162938 4922
rect 162938 4870 162950 4922
rect 162950 4870 162972 4922
rect 162996 4870 163002 4922
rect 163002 4870 163014 4922
rect 163014 4870 163052 4922
rect 163076 4870 163078 4922
rect 163078 4870 163130 4922
rect 163130 4870 163132 4922
rect 163156 4870 163194 4922
rect 163194 4870 163206 4922
rect 163206 4870 163212 4922
rect 163236 4870 163258 4922
rect 163258 4870 163270 4922
rect 163270 4870 163292 4922
rect 163316 4870 163322 4922
rect 163322 4870 163334 4922
rect 163334 4870 163372 4922
rect 162836 4868 162892 4870
rect 162916 4868 162972 4870
rect 162996 4868 163052 4870
rect 163076 4868 163132 4870
rect 163156 4868 163212 4870
rect 163236 4868 163292 4870
rect 163316 4868 163372 4870
rect 162836 3834 162892 3836
rect 162916 3834 162972 3836
rect 162996 3834 163052 3836
rect 163076 3834 163132 3836
rect 163156 3834 163212 3836
rect 163236 3834 163292 3836
rect 163316 3834 163372 3836
rect 162836 3782 162874 3834
rect 162874 3782 162886 3834
rect 162886 3782 162892 3834
rect 162916 3782 162938 3834
rect 162938 3782 162950 3834
rect 162950 3782 162972 3834
rect 162996 3782 163002 3834
rect 163002 3782 163014 3834
rect 163014 3782 163052 3834
rect 163076 3782 163078 3834
rect 163078 3782 163130 3834
rect 163130 3782 163132 3834
rect 163156 3782 163194 3834
rect 163194 3782 163206 3834
rect 163206 3782 163212 3834
rect 163236 3782 163258 3834
rect 163258 3782 163270 3834
rect 163270 3782 163292 3834
rect 163316 3782 163322 3834
rect 163322 3782 163334 3834
rect 163334 3782 163372 3834
rect 162836 3780 162892 3782
rect 162916 3780 162972 3782
rect 162996 3780 163052 3782
rect 163076 3780 163132 3782
rect 163156 3780 163212 3782
rect 163236 3780 163292 3782
rect 163316 3780 163372 3782
rect 162836 2746 162892 2748
rect 162916 2746 162972 2748
rect 162996 2746 163052 2748
rect 163076 2746 163132 2748
rect 163156 2746 163212 2748
rect 163236 2746 163292 2748
rect 163316 2746 163372 2748
rect 162836 2694 162874 2746
rect 162874 2694 162886 2746
rect 162886 2694 162892 2746
rect 162916 2694 162938 2746
rect 162938 2694 162950 2746
rect 162950 2694 162972 2746
rect 162996 2694 163002 2746
rect 163002 2694 163014 2746
rect 163014 2694 163052 2746
rect 163076 2694 163078 2746
rect 163078 2694 163130 2746
rect 163130 2694 163132 2746
rect 163156 2694 163194 2746
rect 163194 2694 163206 2746
rect 163206 2694 163212 2746
rect 163236 2694 163258 2746
rect 163258 2694 163270 2746
rect 163270 2694 163292 2746
rect 163316 2694 163322 2746
rect 163322 2694 163334 2746
rect 163334 2694 163372 2746
rect 162836 2692 162892 2694
rect 162916 2692 162972 2694
rect 162996 2692 163052 2694
rect 163076 2692 163132 2694
rect 163156 2692 163212 2694
rect 163236 2692 163292 2694
rect 163316 2692 163372 2694
rect 180836 5466 180892 5468
rect 180916 5466 180972 5468
rect 180996 5466 181052 5468
rect 181076 5466 181132 5468
rect 181156 5466 181212 5468
rect 181236 5466 181292 5468
rect 181316 5466 181372 5468
rect 180836 5414 180874 5466
rect 180874 5414 180886 5466
rect 180886 5414 180892 5466
rect 180916 5414 180938 5466
rect 180938 5414 180950 5466
rect 180950 5414 180972 5466
rect 180996 5414 181002 5466
rect 181002 5414 181014 5466
rect 181014 5414 181052 5466
rect 181076 5414 181078 5466
rect 181078 5414 181130 5466
rect 181130 5414 181132 5466
rect 181156 5414 181194 5466
rect 181194 5414 181206 5466
rect 181206 5414 181212 5466
rect 181236 5414 181258 5466
rect 181258 5414 181270 5466
rect 181270 5414 181292 5466
rect 181316 5414 181322 5466
rect 181322 5414 181334 5466
rect 181334 5414 181372 5466
rect 180836 5412 180892 5414
rect 180916 5412 180972 5414
rect 180996 5412 181052 5414
rect 181076 5412 181132 5414
rect 181156 5412 181212 5414
rect 181236 5412 181292 5414
rect 181316 5412 181372 5414
rect 180836 4378 180892 4380
rect 180916 4378 180972 4380
rect 180996 4378 181052 4380
rect 181076 4378 181132 4380
rect 181156 4378 181212 4380
rect 181236 4378 181292 4380
rect 181316 4378 181372 4380
rect 180836 4326 180874 4378
rect 180874 4326 180886 4378
rect 180886 4326 180892 4378
rect 180916 4326 180938 4378
rect 180938 4326 180950 4378
rect 180950 4326 180972 4378
rect 180996 4326 181002 4378
rect 181002 4326 181014 4378
rect 181014 4326 181052 4378
rect 181076 4326 181078 4378
rect 181078 4326 181130 4378
rect 181130 4326 181132 4378
rect 181156 4326 181194 4378
rect 181194 4326 181206 4378
rect 181206 4326 181212 4378
rect 181236 4326 181258 4378
rect 181258 4326 181270 4378
rect 181270 4326 181292 4378
rect 181316 4326 181322 4378
rect 181322 4326 181334 4378
rect 181334 4326 181372 4378
rect 180836 4324 180892 4326
rect 180916 4324 180972 4326
rect 180996 4324 181052 4326
rect 181076 4324 181132 4326
rect 181156 4324 181212 4326
rect 181236 4324 181292 4326
rect 181316 4324 181372 4326
rect 180836 3290 180892 3292
rect 180916 3290 180972 3292
rect 180996 3290 181052 3292
rect 181076 3290 181132 3292
rect 181156 3290 181212 3292
rect 181236 3290 181292 3292
rect 181316 3290 181372 3292
rect 180836 3238 180874 3290
rect 180874 3238 180886 3290
rect 180886 3238 180892 3290
rect 180916 3238 180938 3290
rect 180938 3238 180950 3290
rect 180950 3238 180972 3290
rect 180996 3238 181002 3290
rect 181002 3238 181014 3290
rect 181014 3238 181052 3290
rect 181076 3238 181078 3290
rect 181078 3238 181130 3290
rect 181130 3238 181132 3290
rect 181156 3238 181194 3290
rect 181194 3238 181206 3290
rect 181206 3238 181212 3290
rect 181236 3238 181258 3290
rect 181258 3238 181270 3290
rect 181270 3238 181292 3290
rect 181316 3238 181322 3290
rect 181322 3238 181334 3290
rect 181334 3238 181372 3290
rect 180836 3236 180892 3238
rect 180916 3236 180972 3238
rect 180996 3236 181052 3238
rect 181076 3236 181132 3238
rect 181156 3236 181212 3238
rect 181236 3236 181292 3238
rect 181316 3236 181372 3238
rect 180836 2202 180892 2204
rect 180916 2202 180972 2204
rect 180996 2202 181052 2204
rect 181076 2202 181132 2204
rect 181156 2202 181212 2204
rect 181236 2202 181292 2204
rect 181316 2202 181372 2204
rect 180836 2150 180874 2202
rect 180874 2150 180886 2202
rect 180886 2150 180892 2202
rect 180916 2150 180938 2202
rect 180938 2150 180950 2202
rect 180950 2150 180972 2202
rect 180996 2150 181002 2202
rect 181002 2150 181014 2202
rect 181014 2150 181052 2202
rect 181076 2150 181078 2202
rect 181078 2150 181130 2202
rect 181130 2150 181132 2202
rect 181156 2150 181194 2202
rect 181194 2150 181206 2202
rect 181206 2150 181212 2202
rect 181236 2150 181258 2202
rect 181258 2150 181270 2202
rect 181270 2150 181292 2202
rect 181316 2150 181322 2202
rect 181322 2150 181334 2202
rect 181334 2150 181372 2202
rect 180836 2148 180892 2150
rect 180916 2148 180972 2150
rect 180996 2148 181052 2150
rect 181076 2148 181132 2150
rect 181156 2148 181212 2150
rect 181236 2148 181292 2150
rect 181316 2148 181372 2150
rect 198836 6010 198892 6012
rect 198916 6010 198972 6012
rect 198996 6010 199052 6012
rect 199076 6010 199132 6012
rect 199156 6010 199212 6012
rect 199236 6010 199292 6012
rect 199316 6010 199372 6012
rect 198836 5958 198874 6010
rect 198874 5958 198886 6010
rect 198886 5958 198892 6010
rect 198916 5958 198938 6010
rect 198938 5958 198950 6010
rect 198950 5958 198972 6010
rect 198996 5958 199002 6010
rect 199002 5958 199014 6010
rect 199014 5958 199052 6010
rect 199076 5958 199078 6010
rect 199078 5958 199130 6010
rect 199130 5958 199132 6010
rect 199156 5958 199194 6010
rect 199194 5958 199206 6010
rect 199206 5958 199212 6010
rect 199236 5958 199258 6010
rect 199258 5958 199270 6010
rect 199270 5958 199292 6010
rect 199316 5958 199322 6010
rect 199322 5958 199334 6010
rect 199334 5958 199372 6010
rect 198836 5956 198892 5958
rect 198916 5956 198972 5958
rect 198996 5956 199052 5958
rect 199076 5956 199132 5958
rect 199156 5956 199212 5958
rect 199236 5956 199292 5958
rect 199316 5956 199372 5958
rect 198836 4922 198892 4924
rect 198916 4922 198972 4924
rect 198996 4922 199052 4924
rect 199076 4922 199132 4924
rect 199156 4922 199212 4924
rect 199236 4922 199292 4924
rect 199316 4922 199372 4924
rect 198836 4870 198874 4922
rect 198874 4870 198886 4922
rect 198886 4870 198892 4922
rect 198916 4870 198938 4922
rect 198938 4870 198950 4922
rect 198950 4870 198972 4922
rect 198996 4870 199002 4922
rect 199002 4870 199014 4922
rect 199014 4870 199052 4922
rect 199076 4870 199078 4922
rect 199078 4870 199130 4922
rect 199130 4870 199132 4922
rect 199156 4870 199194 4922
rect 199194 4870 199206 4922
rect 199206 4870 199212 4922
rect 199236 4870 199258 4922
rect 199258 4870 199270 4922
rect 199270 4870 199292 4922
rect 199316 4870 199322 4922
rect 199322 4870 199334 4922
rect 199334 4870 199372 4922
rect 198836 4868 198892 4870
rect 198916 4868 198972 4870
rect 198996 4868 199052 4870
rect 199076 4868 199132 4870
rect 199156 4868 199212 4870
rect 199236 4868 199292 4870
rect 199316 4868 199372 4870
rect 198836 3834 198892 3836
rect 198916 3834 198972 3836
rect 198996 3834 199052 3836
rect 199076 3834 199132 3836
rect 199156 3834 199212 3836
rect 199236 3834 199292 3836
rect 199316 3834 199372 3836
rect 198836 3782 198874 3834
rect 198874 3782 198886 3834
rect 198886 3782 198892 3834
rect 198916 3782 198938 3834
rect 198938 3782 198950 3834
rect 198950 3782 198972 3834
rect 198996 3782 199002 3834
rect 199002 3782 199014 3834
rect 199014 3782 199052 3834
rect 199076 3782 199078 3834
rect 199078 3782 199130 3834
rect 199130 3782 199132 3834
rect 199156 3782 199194 3834
rect 199194 3782 199206 3834
rect 199206 3782 199212 3834
rect 199236 3782 199258 3834
rect 199258 3782 199270 3834
rect 199270 3782 199292 3834
rect 199316 3782 199322 3834
rect 199322 3782 199334 3834
rect 199334 3782 199372 3834
rect 198836 3780 198892 3782
rect 198916 3780 198972 3782
rect 198996 3780 199052 3782
rect 199076 3780 199132 3782
rect 199156 3780 199212 3782
rect 199236 3780 199292 3782
rect 199316 3780 199372 3782
rect 198836 2746 198892 2748
rect 198916 2746 198972 2748
rect 198996 2746 199052 2748
rect 199076 2746 199132 2748
rect 199156 2746 199212 2748
rect 199236 2746 199292 2748
rect 199316 2746 199372 2748
rect 198836 2694 198874 2746
rect 198874 2694 198886 2746
rect 198886 2694 198892 2746
rect 198916 2694 198938 2746
rect 198938 2694 198950 2746
rect 198950 2694 198972 2746
rect 198996 2694 199002 2746
rect 199002 2694 199014 2746
rect 199014 2694 199052 2746
rect 199076 2694 199078 2746
rect 199078 2694 199130 2746
rect 199130 2694 199132 2746
rect 199156 2694 199194 2746
rect 199194 2694 199206 2746
rect 199206 2694 199212 2746
rect 199236 2694 199258 2746
rect 199258 2694 199270 2746
rect 199270 2694 199292 2746
rect 199316 2694 199322 2746
rect 199322 2694 199334 2746
rect 199334 2694 199372 2746
rect 198836 2692 198892 2694
rect 198916 2692 198972 2694
rect 198996 2692 199052 2694
rect 199076 2692 199132 2694
rect 199156 2692 199212 2694
rect 199236 2692 199292 2694
rect 199316 2692 199372 2694
rect 216836 5466 216892 5468
rect 216916 5466 216972 5468
rect 216996 5466 217052 5468
rect 217076 5466 217132 5468
rect 217156 5466 217212 5468
rect 217236 5466 217292 5468
rect 217316 5466 217372 5468
rect 216836 5414 216874 5466
rect 216874 5414 216886 5466
rect 216886 5414 216892 5466
rect 216916 5414 216938 5466
rect 216938 5414 216950 5466
rect 216950 5414 216972 5466
rect 216996 5414 217002 5466
rect 217002 5414 217014 5466
rect 217014 5414 217052 5466
rect 217076 5414 217078 5466
rect 217078 5414 217130 5466
rect 217130 5414 217132 5466
rect 217156 5414 217194 5466
rect 217194 5414 217206 5466
rect 217206 5414 217212 5466
rect 217236 5414 217258 5466
rect 217258 5414 217270 5466
rect 217270 5414 217292 5466
rect 217316 5414 217322 5466
rect 217322 5414 217334 5466
rect 217334 5414 217372 5466
rect 216836 5412 216892 5414
rect 216916 5412 216972 5414
rect 216996 5412 217052 5414
rect 217076 5412 217132 5414
rect 217156 5412 217212 5414
rect 217236 5412 217292 5414
rect 217316 5412 217372 5414
rect 216836 4378 216892 4380
rect 216916 4378 216972 4380
rect 216996 4378 217052 4380
rect 217076 4378 217132 4380
rect 217156 4378 217212 4380
rect 217236 4378 217292 4380
rect 217316 4378 217372 4380
rect 216836 4326 216874 4378
rect 216874 4326 216886 4378
rect 216886 4326 216892 4378
rect 216916 4326 216938 4378
rect 216938 4326 216950 4378
rect 216950 4326 216972 4378
rect 216996 4326 217002 4378
rect 217002 4326 217014 4378
rect 217014 4326 217052 4378
rect 217076 4326 217078 4378
rect 217078 4326 217130 4378
rect 217130 4326 217132 4378
rect 217156 4326 217194 4378
rect 217194 4326 217206 4378
rect 217206 4326 217212 4378
rect 217236 4326 217258 4378
rect 217258 4326 217270 4378
rect 217270 4326 217292 4378
rect 217316 4326 217322 4378
rect 217322 4326 217334 4378
rect 217334 4326 217372 4378
rect 216836 4324 216892 4326
rect 216916 4324 216972 4326
rect 216996 4324 217052 4326
rect 217076 4324 217132 4326
rect 217156 4324 217212 4326
rect 217236 4324 217292 4326
rect 217316 4324 217372 4326
rect 216836 3290 216892 3292
rect 216916 3290 216972 3292
rect 216996 3290 217052 3292
rect 217076 3290 217132 3292
rect 217156 3290 217212 3292
rect 217236 3290 217292 3292
rect 217316 3290 217372 3292
rect 216836 3238 216874 3290
rect 216874 3238 216886 3290
rect 216886 3238 216892 3290
rect 216916 3238 216938 3290
rect 216938 3238 216950 3290
rect 216950 3238 216972 3290
rect 216996 3238 217002 3290
rect 217002 3238 217014 3290
rect 217014 3238 217052 3290
rect 217076 3238 217078 3290
rect 217078 3238 217130 3290
rect 217130 3238 217132 3290
rect 217156 3238 217194 3290
rect 217194 3238 217206 3290
rect 217206 3238 217212 3290
rect 217236 3238 217258 3290
rect 217258 3238 217270 3290
rect 217270 3238 217292 3290
rect 217316 3238 217322 3290
rect 217322 3238 217334 3290
rect 217334 3238 217372 3290
rect 216836 3236 216892 3238
rect 216916 3236 216972 3238
rect 216996 3236 217052 3238
rect 217076 3236 217132 3238
rect 217156 3236 217212 3238
rect 217236 3236 217292 3238
rect 217316 3236 217372 3238
rect 216836 2202 216892 2204
rect 216916 2202 216972 2204
rect 216996 2202 217052 2204
rect 217076 2202 217132 2204
rect 217156 2202 217212 2204
rect 217236 2202 217292 2204
rect 217316 2202 217372 2204
rect 216836 2150 216874 2202
rect 216874 2150 216886 2202
rect 216886 2150 216892 2202
rect 216916 2150 216938 2202
rect 216938 2150 216950 2202
rect 216950 2150 216972 2202
rect 216996 2150 217002 2202
rect 217002 2150 217014 2202
rect 217014 2150 217052 2202
rect 217076 2150 217078 2202
rect 217078 2150 217130 2202
rect 217130 2150 217132 2202
rect 217156 2150 217194 2202
rect 217194 2150 217206 2202
rect 217206 2150 217212 2202
rect 217236 2150 217258 2202
rect 217258 2150 217270 2202
rect 217270 2150 217292 2202
rect 217316 2150 217322 2202
rect 217322 2150 217334 2202
rect 217334 2150 217372 2202
rect 216836 2148 216892 2150
rect 216916 2148 216972 2150
rect 216996 2148 217052 2150
rect 217076 2148 217132 2150
rect 217156 2148 217212 2150
rect 217236 2148 217292 2150
rect 217316 2148 217372 2150
rect 234836 6010 234892 6012
rect 234916 6010 234972 6012
rect 234996 6010 235052 6012
rect 235076 6010 235132 6012
rect 235156 6010 235212 6012
rect 235236 6010 235292 6012
rect 235316 6010 235372 6012
rect 234836 5958 234874 6010
rect 234874 5958 234886 6010
rect 234886 5958 234892 6010
rect 234916 5958 234938 6010
rect 234938 5958 234950 6010
rect 234950 5958 234972 6010
rect 234996 5958 235002 6010
rect 235002 5958 235014 6010
rect 235014 5958 235052 6010
rect 235076 5958 235078 6010
rect 235078 5958 235130 6010
rect 235130 5958 235132 6010
rect 235156 5958 235194 6010
rect 235194 5958 235206 6010
rect 235206 5958 235212 6010
rect 235236 5958 235258 6010
rect 235258 5958 235270 6010
rect 235270 5958 235292 6010
rect 235316 5958 235322 6010
rect 235322 5958 235334 6010
rect 235334 5958 235372 6010
rect 234836 5956 234892 5958
rect 234916 5956 234972 5958
rect 234996 5956 235052 5958
rect 235076 5956 235132 5958
rect 235156 5956 235212 5958
rect 235236 5956 235292 5958
rect 235316 5956 235372 5958
rect 234836 4922 234892 4924
rect 234916 4922 234972 4924
rect 234996 4922 235052 4924
rect 235076 4922 235132 4924
rect 235156 4922 235212 4924
rect 235236 4922 235292 4924
rect 235316 4922 235372 4924
rect 234836 4870 234874 4922
rect 234874 4870 234886 4922
rect 234886 4870 234892 4922
rect 234916 4870 234938 4922
rect 234938 4870 234950 4922
rect 234950 4870 234972 4922
rect 234996 4870 235002 4922
rect 235002 4870 235014 4922
rect 235014 4870 235052 4922
rect 235076 4870 235078 4922
rect 235078 4870 235130 4922
rect 235130 4870 235132 4922
rect 235156 4870 235194 4922
rect 235194 4870 235206 4922
rect 235206 4870 235212 4922
rect 235236 4870 235258 4922
rect 235258 4870 235270 4922
rect 235270 4870 235292 4922
rect 235316 4870 235322 4922
rect 235322 4870 235334 4922
rect 235334 4870 235372 4922
rect 234836 4868 234892 4870
rect 234916 4868 234972 4870
rect 234996 4868 235052 4870
rect 235076 4868 235132 4870
rect 235156 4868 235212 4870
rect 235236 4868 235292 4870
rect 235316 4868 235372 4870
rect 234836 3834 234892 3836
rect 234916 3834 234972 3836
rect 234996 3834 235052 3836
rect 235076 3834 235132 3836
rect 235156 3834 235212 3836
rect 235236 3834 235292 3836
rect 235316 3834 235372 3836
rect 234836 3782 234874 3834
rect 234874 3782 234886 3834
rect 234886 3782 234892 3834
rect 234916 3782 234938 3834
rect 234938 3782 234950 3834
rect 234950 3782 234972 3834
rect 234996 3782 235002 3834
rect 235002 3782 235014 3834
rect 235014 3782 235052 3834
rect 235076 3782 235078 3834
rect 235078 3782 235130 3834
rect 235130 3782 235132 3834
rect 235156 3782 235194 3834
rect 235194 3782 235206 3834
rect 235206 3782 235212 3834
rect 235236 3782 235258 3834
rect 235258 3782 235270 3834
rect 235270 3782 235292 3834
rect 235316 3782 235322 3834
rect 235322 3782 235334 3834
rect 235334 3782 235372 3834
rect 234836 3780 234892 3782
rect 234916 3780 234972 3782
rect 234996 3780 235052 3782
rect 235076 3780 235132 3782
rect 235156 3780 235212 3782
rect 235236 3780 235292 3782
rect 235316 3780 235372 3782
rect 234836 2746 234892 2748
rect 234916 2746 234972 2748
rect 234996 2746 235052 2748
rect 235076 2746 235132 2748
rect 235156 2746 235212 2748
rect 235236 2746 235292 2748
rect 235316 2746 235372 2748
rect 234836 2694 234874 2746
rect 234874 2694 234886 2746
rect 234886 2694 234892 2746
rect 234916 2694 234938 2746
rect 234938 2694 234950 2746
rect 234950 2694 234972 2746
rect 234996 2694 235002 2746
rect 235002 2694 235014 2746
rect 235014 2694 235052 2746
rect 235076 2694 235078 2746
rect 235078 2694 235130 2746
rect 235130 2694 235132 2746
rect 235156 2694 235194 2746
rect 235194 2694 235206 2746
rect 235206 2694 235212 2746
rect 235236 2694 235258 2746
rect 235258 2694 235270 2746
rect 235270 2694 235292 2746
rect 235316 2694 235322 2746
rect 235322 2694 235334 2746
rect 235334 2694 235372 2746
rect 234836 2692 234892 2694
rect 234916 2692 234972 2694
rect 234996 2692 235052 2694
rect 235076 2692 235132 2694
rect 235156 2692 235212 2694
rect 235236 2692 235292 2694
rect 235316 2692 235372 2694
rect 252836 5466 252892 5468
rect 252916 5466 252972 5468
rect 252996 5466 253052 5468
rect 253076 5466 253132 5468
rect 253156 5466 253212 5468
rect 253236 5466 253292 5468
rect 253316 5466 253372 5468
rect 252836 5414 252874 5466
rect 252874 5414 252886 5466
rect 252886 5414 252892 5466
rect 252916 5414 252938 5466
rect 252938 5414 252950 5466
rect 252950 5414 252972 5466
rect 252996 5414 253002 5466
rect 253002 5414 253014 5466
rect 253014 5414 253052 5466
rect 253076 5414 253078 5466
rect 253078 5414 253130 5466
rect 253130 5414 253132 5466
rect 253156 5414 253194 5466
rect 253194 5414 253206 5466
rect 253206 5414 253212 5466
rect 253236 5414 253258 5466
rect 253258 5414 253270 5466
rect 253270 5414 253292 5466
rect 253316 5414 253322 5466
rect 253322 5414 253334 5466
rect 253334 5414 253372 5466
rect 252836 5412 252892 5414
rect 252916 5412 252972 5414
rect 252996 5412 253052 5414
rect 253076 5412 253132 5414
rect 253156 5412 253212 5414
rect 253236 5412 253292 5414
rect 253316 5412 253372 5414
rect 252836 4378 252892 4380
rect 252916 4378 252972 4380
rect 252996 4378 253052 4380
rect 253076 4378 253132 4380
rect 253156 4378 253212 4380
rect 253236 4378 253292 4380
rect 253316 4378 253372 4380
rect 252836 4326 252874 4378
rect 252874 4326 252886 4378
rect 252886 4326 252892 4378
rect 252916 4326 252938 4378
rect 252938 4326 252950 4378
rect 252950 4326 252972 4378
rect 252996 4326 253002 4378
rect 253002 4326 253014 4378
rect 253014 4326 253052 4378
rect 253076 4326 253078 4378
rect 253078 4326 253130 4378
rect 253130 4326 253132 4378
rect 253156 4326 253194 4378
rect 253194 4326 253206 4378
rect 253206 4326 253212 4378
rect 253236 4326 253258 4378
rect 253258 4326 253270 4378
rect 253270 4326 253292 4378
rect 253316 4326 253322 4378
rect 253322 4326 253334 4378
rect 253334 4326 253372 4378
rect 252836 4324 252892 4326
rect 252916 4324 252972 4326
rect 252996 4324 253052 4326
rect 253076 4324 253132 4326
rect 253156 4324 253212 4326
rect 253236 4324 253292 4326
rect 253316 4324 253372 4326
rect 252836 3290 252892 3292
rect 252916 3290 252972 3292
rect 252996 3290 253052 3292
rect 253076 3290 253132 3292
rect 253156 3290 253212 3292
rect 253236 3290 253292 3292
rect 253316 3290 253372 3292
rect 252836 3238 252874 3290
rect 252874 3238 252886 3290
rect 252886 3238 252892 3290
rect 252916 3238 252938 3290
rect 252938 3238 252950 3290
rect 252950 3238 252972 3290
rect 252996 3238 253002 3290
rect 253002 3238 253014 3290
rect 253014 3238 253052 3290
rect 253076 3238 253078 3290
rect 253078 3238 253130 3290
rect 253130 3238 253132 3290
rect 253156 3238 253194 3290
rect 253194 3238 253206 3290
rect 253206 3238 253212 3290
rect 253236 3238 253258 3290
rect 253258 3238 253270 3290
rect 253270 3238 253292 3290
rect 253316 3238 253322 3290
rect 253322 3238 253334 3290
rect 253334 3238 253372 3290
rect 252836 3236 252892 3238
rect 252916 3236 252972 3238
rect 252996 3236 253052 3238
rect 253076 3236 253132 3238
rect 253156 3236 253212 3238
rect 253236 3236 253292 3238
rect 253316 3236 253372 3238
rect 252836 2202 252892 2204
rect 252916 2202 252972 2204
rect 252996 2202 253052 2204
rect 253076 2202 253132 2204
rect 253156 2202 253212 2204
rect 253236 2202 253292 2204
rect 253316 2202 253372 2204
rect 252836 2150 252874 2202
rect 252874 2150 252886 2202
rect 252886 2150 252892 2202
rect 252916 2150 252938 2202
rect 252938 2150 252950 2202
rect 252950 2150 252972 2202
rect 252996 2150 253002 2202
rect 253002 2150 253014 2202
rect 253014 2150 253052 2202
rect 253076 2150 253078 2202
rect 253078 2150 253130 2202
rect 253130 2150 253132 2202
rect 253156 2150 253194 2202
rect 253194 2150 253206 2202
rect 253206 2150 253212 2202
rect 253236 2150 253258 2202
rect 253258 2150 253270 2202
rect 253270 2150 253292 2202
rect 253316 2150 253322 2202
rect 253322 2150 253334 2202
rect 253334 2150 253372 2202
rect 252836 2148 252892 2150
rect 252916 2148 252972 2150
rect 252996 2148 253052 2150
rect 253076 2148 253132 2150
rect 253156 2148 253212 2150
rect 253236 2148 253292 2150
rect 253316 2148 253372 2150
rect 270836 6010 270892 6012
rect 270916 6010 270972 6012
rect 270996 6010 271052 6012
rect 271076 6010 271132 6012
rect 271156 6010 271212 6012
rect 271236 6010 271292 6012
rect 271316 6010 271372 6012
rect 270836 5958 270874 6010
rect 270874 5958 270886 6010
rect 270886 5958 270892 6010
rect 270916 5958 270938 6010
rect 270938 5958 270950 6010
rect 270950 5958 270972 6010
rect 270996 5958 271002 6010
rect 271002 5958 271014 6010
rect 271014 5958 271052 6010
rect 271076 5958 271078 6010
rect 271078 5958 271130 6010
rect 271130 5958 271132 6010
rect 271156 5958 271194 6010
rect 271194 5958 271206 6010
rect 271206 5958 271212 6010
rect 271236 5958 271258 6010
rect 271258 5958 271270 6010
rect 271270 5958 271292 6010
rect 271316 5958 271322 6010
rect 271322 5958 271334 6010
rect 271334 5958 271372 6010
rect 270836 5956 270892 5958
rect 270916 5956 270972 5958
rect 270996 5956 271052 5958
rect 271076 5956 271132 5958
rect 271156 5956 271212 5958
rect 271236 5956 271292 5958
rect 271316 5956 271372 5958
rect 270836 4922 270892 4924
rect 270916 4922 270972 4924
rect 270996 4922 271052 4924
rect 271076 4922 271132 4924
rect 271156 4922 271212 4924
rect 271236 4922 271292 4924
rect 271316 4922 271372 4924
rect 270836 4870 270874 4922
rect 270874 4870 270886 4922
rect 270886 4870 270892 4922
rect 270916 4870 270938 4922
rect 270938 4870 270950 4922
rect 270950 4870 270972 4922
rect 270996 4870 271002 4922
rect 271002 4870 271014 4922
rect 271014 4870 271052 4922
rect 271076 4870 271078 4922
rect 271078 4870 271130 4922
rect 271130 4870 271132 4922
rect 271156 4870 271194 4922
rect 271194 4870 271206 4922
rect 271206 4870 271212 4922
rect 271236 4870 271258 4922
rect 271258 4870 271270 4922
rect 271270 4870 271292 4922
rect 271316 4870 271322 4922
rect 271322 4870 271334 4922
rect 271334 4870 271372 4922
rect 270836 4868 270892 4870
rect 270916 4868 270972 4870
rect 270996 4868 271052 4870
rect 271076 4868 271132 4870
rect 271156 4868 271212 4870
rect 271236 4868 271292 4870
rect 271316 4868 271372 4870
rect 270836 3834 270892 3836
rect 270916 3834 270972 3836
rect 270996 3834 271052 3836
rect 271076 3834 271132 3836
rect 271156 3834 271212 3836
rect 271236 3834 271292 3836
rect 271316 3834 271372 3836
rect 270836 3782 270874 3834
rect 270874 3782 270886 3834
rect 270886 3782 270892 3834
rect 270916 3782 270938 3834
rect 270938 3782 270950 3834
rect 270950 3782 270972 3834
rect 270996 3782 271002 3834
rect 271002 3782 271014 3834
rect 271014 3782 271052 3834
rect 271076 3782 271078 3834
rect 271078 3782 271130 3834
rect 271130 3782 271132 3834
rect 271156 3782 271194 3834
rect 271194 3782 271206 3834
rect 271206 3782 271212 3834
rect 271236 3782 271258 3834
rect 271258 3782 271270 3834
rect 271270 3782 271292 3834
rect 271316 3782 271322 3834
rect 271322 3782 271334 3834
rect 271334 3782 271372 3834
rect 270836 3780 270892 3782
rect 270916 3780 270972 3782
rect 270996 3780 271052 3782
rect 271076 3780 271132 3782
rect 271156 3780 271212 3782
rect 271236 3780 271292 3782
rect 271316 3780 271372 3782
rect 270836 2746 270892 2748
rect 270916 2746 270972 2748
rect 270996 2746 271052 2748
rect 271076 2746 271132 2748
rect 271156 2746 271212 2748
rect 271236 2746 271292 2748
rect 271316 2746 271372 2748
rect 270836 2694 270874 2746
rect 270874 2694 270886 2746
rect 270886 2694 270892 2746
rect 270916 2694 270938 2746
rect 270938 2694 270950 2746
rect 270950 2694 270972 2746
rect 270996 2694 271002 2746
rect 271002 2694 271014 2746
rect 271014 2694 271052 2746
rect 271076 2694 271078 2746
rect 271078 2694 271130 2746
rect 271130 2694 271132 2746
rect 271156 2694 271194 2746
rect 271194 2694 271206 2746
rect 271206 2694 271212 2746
rect 271236 2694 271258 2746
rect 271258 2694 271270 2746
rect 271270 2694 271292 2746
rect 271316 2694 271322 2746
rect 271322 2694 271334 2746
rect 271334 2694 271372 2746
rect 270836 2692 270892 2694
rect 270916 2692 270972 2694
rect 270996 2692 271052 2694
rect 271076 2692 271132 2694
rect 271156 2692 271212 2694
rect 271236 2692 271292 2694
rect 271316 2692 271372 2694
rect 288836 5466 288892 5468
rect 288916 5466 288972 5468
rect 288996 5466 289052 5468
rect 289076 5466 289132 5468
rect 289156 5466 289212 5468
rect 289236 5466 289292 5468
rect 289316 5466 289372 5468
rect 288836 5414 288874 5466
rect 288874 5414 288886 5466
rect 288886 5414 288892 5466
rect 288916 5414 288938 5466
rect 288938 5414 288950 5466
rect 288950 5414 288972 5466
rect 288996 5414 289002 5466
rect 289002 5414 289014 5466
rect 289014 5414 289052 5466
rect 289076 5414 289078 5466
rect 289078 5414 289130 5466
rect 289130 5414 289132 5466
rect 289156 5414 289194 5466
rect 289194 5414 289206 5466
rect 289206 5414 289212 5466
rect 289236 5414 289258 5466
rect 289258 5414 289270 5466
rect 289270 5414 289292 5466
rect 289316 5414 289322 5466
rect 289322 5414 289334 5466
rect 289334 5414 289372 5466
rect 288836 5412 288892 5414
rect 288916 5412 288972 5414
rect 288996 5412 289052 5414
rect 289076 5412 289132 5414
rect 289156 5412 289212 5414
rect 289236 5412 289292 5414
rect 289316 5412 289372 5414
rect 288836 4378 288892 4380
rect 288916 4378 288972 4380
rect 288996 4378 289052 4380
rect 289076 4378 289132 4380
rect 289156 4378 289212 4380
rect 289236 4378 289292 4380
rect 289316 4378 289372 4380
rect 288836 4326 288874 4378
rect 288874 4326 288886 4378
rect 288886 4326 288892 4378
rect 288916 4326 288938 4378
rect 288938 4326 288950 4378
rect 288950 4326 288972 4378
rect 288996 4326 289002 4378
rect 289002 4326 289014 4378
rect 289014 4326 289052 4378
rect 289076 4326 289078 4378
rect 289078 4326 289130 4378
rect 289130 4326 289132 4378
rect 289156 4326 289194 4378
rect 289194 4326 289206 4378
rect 289206 4326 289212 4378
rect 289236 4326 289258 4378
rect 289258 4326 289270 4378
rect 289270 4326 289292 4378
rect 289316 4326 289322 4378
rect 289322 4326 289334 4378
rect 289334 4326 289372 4378
rect 288836 4324 288892 4326
rect 288916 4324 288972 4326
rect 288996 4324 289052 4326
rect 289076 4324 289132 4326
rect 289156 4324 289212 4326
rect 289236 4324 289292 4326
rect 289316 4324 289372 4326
rect 288836 3290 288892 3292
rect 288916 3290 288972 3292
rect 288996 3290 289052 3292
rect 289076 3290 289132 3292
rect 289156 3290 289212 3292
rect 289236 3290 289292 3292
rect 289316 3290 289372 3292
rect 288836 3238 288874 3290
rect 288874 3238 288886 3290
rect 288886 3238 288892 3290
rect 288916 3238 288938 3290
rect 288938 3238 288950 3290
rect 288950 3238 288972 3290
rect 288996 3238 289002 3290
rect 289002 3238 289014 3290
rect 289014 3238 289052 3290
rect 289076 3238 289078 3290
rect 289078 3238 289130 3290
rect 289130 3238 289132 3290
rect 289156 3238 289194 3290
rect 289194 3238 289206 3290
rect 289206 3238 289212 3290
rect 289236 3238 289258 3290
rect 289258 3238 289270 3290
rect 289270 3238 289292 3290
rect 289316 3238 289322 3290
rect 289322 3238 289334 3290
rect 289334 3238 289372 3290
rect 288836 3236 288892 3238
rect 288916 3236 288972 3238
rect 288996 3236 289052 3238
rect 289076 3236 289132 3238
rect 289156 3236 289212 3238
rect 289236 3236 289292 3238
rect 289316 3236 289372 3238
rect 288836 2202 288892 2204
rect 288916 2202 288972 2204
rect 288996 2202 289052 2204
rect 289076 2202 289132 2204
rect 289156 2202 289212 2204
rect 289236 2202 289292 2204
rect 289316 2202 289372 2204
rect 288836 2150 288874 2202
rect 288874 2150 288886 2202
rect 288886 2150 288892 2202
rect 288916 2150 288938 2202
rect 288938 2150 288950 2202
rect 288950 2150 288972 2202
rect 288996 2150 289002 2202
rect 289002 2150 289014 2202
rect 289014 2150 289052 2202
rect 289076 2150 289078 2202
rect 289078 2150 289130 2202
rect 289130 2150 289132 2202
rect 289156 2150 289194 2202
rect 289194 2150 289206 2202
rect 289206 2150 289212 2202
rect 289236 2150 289258 2202
rect 289258 2150 289270 2202
rect 289270 2150 289292 2202
rect 289316 2150 289322 2202
rect 289322 2150 289334 2202
rect 289334 2150 289372 2202
rect 288836 2148 288892 2150
rect 288916 2148 288972 2150
rect 288996 2148 289052 2150
rect 289076 2148 289132 2150
rect 289156 2148 289212 2150
rect 289236 2148 289292 2150
rect 289316 2148 289372 2150
rect 306836 6010 306892 6012
rect 306916 6010 306972 6012
rect 306996 6010 307052 6012
rect 307076 6010 307132 6012
rect 307156 6010 307212 6012
rect 307236 6010 307292 6012
rect 307316 6010 307372 6012
rect 306836 5958 306874 6010
rect 306874 5958 306886 6010
rect 306886 5958 306892 6010
rect 306916 5958 306938 6010
rect 306938 5958 306950 6010
rect 306950 5958 306972 6010
rect 306996 5958 307002 6010
rect 307002 5958 307014 6010
rect 307014 5958 307052 6010
rect 307076 5958 307078 6010
rect 307078 5958 307130 6010
rect 307130 5958 307132 6010
rect 307156 5958 307194 6010
rect 307194 5958 307206 6010
rect 307206 5958 307212 6010
rect 307236 5958 307258 6010
rect 307258 5958 307270 6010
rect 307270 5958 307292 6010
rect 307316 5958 307322 6010
rect 307322 5958 307334 6010
rect 307334 5958 307372 6010
rect 306836 5956 306892 5958
rect 306916 5956 306972 5958
rect 306996 5956 307052 5958
rect 307076 5956 307132 5958
rect 307156 5956 307212 5958
rect 307236 5956 307292 5958
rect 307316 5956 307372 5958
rect 306836 4922 306892 4924
rect 306916 4922 306972 4924
rect 306996 4922 307052 4924
rect 307076 4922 307132 4924
rect 307156 4922 307212 4924
rect 307236 4922 307292 4924
rect 307316 4922 307372 4924
rect 306836 4870 306874 4922
rect 306874 4870 306886 4922
rect 306886 4870 306892 4922
rect 306916 4870 306938 4922
rect 306938 4870 306950 4922
rect 306950 4870 306972 4922
rect 306996 4870 307002 4922
rect 307002 4870 307014 4922
rect 307014 4870 307052 4922
rect 307076 4870 307078 4922
rect 307078 4870 307130 4922
rect 307130 4870 307132 4922
rect 307156 4870 307194 4922
rect 307194 4870 307206 4922
rect 307206 4870 307212 4922
rect 307236 4870 307258 4922
rect 307258 4870 307270 4922
rect 307270 4870 307292 4922
rect 307316 4870 307322 4922
rect 307322 4870 307334 4922
rect 307334 4870 307372 4922
rect 306836 4868 306892 4870
rect 306916 4868 306972 4870
rect 306996 4868 307052 4870
rect 307076 4868 307132 4870
rect 307156 4868 307212 4870
rect 307236 4868 307292 4870
rect 307316 4868 307372 4870
rect 306836 3834 306892 3836
rect 306916 3834 306972 3836
rect 306996 3834 307052 3836
rect 307076 3834 307132 3836
rect 307156 3834 307212 3836
rect 307236 3834 307292 3836
rect 307316 3834 307372 3836
rect 306836 3782 306874 3834
rect 306874 3782 306886 3834
rect 306886 3782 306892 3834
rect 306916 3782 306938 3834
rect 306938 3782 306950 3834
rect 306950 3782 306972 3834
rect 306996 3782 307002 3834
rect 307002 3782 307014 3834
rect 307014 3782 307052 3834
rect 307076 3782 307078 3834
rect 307078 3782 307130 3834
rect 307130 3782 307132 3834
rect 307156 3782 307194 3834
rect 307194 3782 307206 3834
rect 307206 3782 307212 3834
rect 307236 3782 307258 3834
rect 307258 3782 307270 3834
rect 307270 3782 307292 3834
rect 307316 3782 307322 3834
rect 307322 3782 307334 3834
rect 307334 3782 307372 3834
rect 306836 3780 306892 3782
rect 306916 3780 306972 3782
rect 306996 3780 307052 3782
rect 307076 3780 307132 3782
rect 307156 3780 307212 3782
rect 307236 3780 307292 3782
rect 307316 3780 307372 3782
rect 306836 2746 306892 2748
rect 306916 2746 306972 2748
rect 306996 2746 307052 2748
rect 307076 2746 307132 2748
rect 307156 2746 307212 2748
rect 307236 2746 307292 2748
rect 307316 2746 307372 2748
rect 306836 2694 306874 2746
rect 306874 2694 306886 2746
rect 306886 2694 306892 2746
rect 306916 2694 306938 2746
rect 306938 2694 306950 2746
rect 306950 2694 306972 2746
rect 306996 2694 307002 2746
rect 307002 2694 307014 2746
rect 307014 2694 307052 2746
rect 307076 2694 307078 2746
rect 307078 2694 307130 2746
rect 307130 2694 307132 2746
rect 307156 2694 307194 2746
rect 307194 2694 307206 2746
rect 307206 2694 307212 2746
rect 307236 2694 307258 2746
rect 307258 2694 307270 2746
rect 307270 2694 307292 2746
rect 307316 2694 307322 2746
rect 307322 2694 307334 2746
rect 307334 2694 307372 2746
rect 306836 2692 306892 2694
rect 306916 2692 306972 2694
rect 306996 2692 307052 2694
rect 307076 2692 307132 2694
rect 307156 2692 307212 2694
rect 307236 2692 307292 2694
rect 307316 2692 307372 2694
rect 324836 5466 324892 5468
rect 324916 5466 324972 5468
rect 324996 5466 325052 5468
rect 325076 5466 325132 5468
rect 325156 5466 325212 5468
rect 325236 5466 325292 5468
rect 325316 5466 325372 5468
rect 324836 5414 324874 5466
rect 324874 5414 324886 5466
rect 324886 5414 324892 5466
rect 324916 5414 324938 5466
rect 324938 5414 324950 5466
rect 324950 5414 324972 5466
rect 324996 5414 325002 5466
rect 325002 5414 325014 5466
rect 325014 5414 325052 5466
rect 325076 5414 325078 5466
rect 325078 5414 325130 5466
rect 325130 5414 325132 5466
rect 325156 5414 325194 5466
rect 325194 5414 325206 5466
rect 325206 5414 325212 5466
rect 325236 5414 325258 5466
rect 325258 5414 325270 5466
rect 325270 5414 325292 5466
rect 325316 5414 325322 5466
rect 325322 5414 325334 5466
rect 325334 5414 325372 5466
rect 324836 5412 324892 5414
rect 324916 5412 324972 5414
rect 324996 5412 325052 5414
rect 325076 5412 325132 5414
rect 325156 5412 325212 5414
rect 325236 5412 325292 5414
rect 325316 5412 325372 5414
rect 324836 4378 324892 4380
rect 324916 4378 324972 4380
rect 324996 4378 325052 4380
rect 325076 4378 325132 4380
rect 325156 4378 325212 4380
rect 325236 4378 325292 4380
rect 325316 4378 325372 4380
rect 324836 4326 324874 4378
rect 324874 4326 324886 4378
rect 324886 4326 324892 4378
rect 324916 4326 324938 4378
rect 324938 4326 324950 4378
rect 324950 4326 324972 4378
rect 324996 4326 325002 4378
rect 325002 4326 325014 4378
rect 325014 4326 325052 4378
rect 325076 4326 325078 4378
rect 325078 4326 325130 4378
rect 325130 4326 325132 4378
rect 325156 4326 325194 4378
rect 325194 4326 325206 4378
rect 325206 4326 325212 4378
rect 325236 4326 325258 4378
rect 325258 4326 325270 4378
rect 325270 4326 325292 4378
rect 325316 4326 325322 4378
rect 325322 4326 325334 4378
rect 325334 4326 325372 4378
rect 324836 4324 324892 4326
rect 324916 4324 324972 4326
rect 324996 4324 325052 4326
rect 325076 4324 325132 4326
rect 325156 4324 325212 4326
rect 325236 4324 325292 4326
rect 325316 4324 325372 4326
rect 324836 3290 324892 3292
rect 324916 3290 324972 3292
rect 324996 3290 325052 3292
rect 325076 3290 325132 3292
rect 325156 3290 325212 3292
rect 325236 3290 325292 3292
rect 325316 3290 325372 3292
rect 324836 3238 324874 3290
rect 324874 3238 324886 3290
rect 324886 3238 324892 3290
rect 324916 3238 324938 3290
rect 324938 3238 324950 3290
rect 324950 3238 324972 3290
rect 324996 3238 325002 3290
rect 325002 3238 325014 3290
rect 325014 3238 325052 3290
rect 325076 3238 325078 3290
rect 325078 3238 325130 3290
rect 325130 3238 325132 3290
rect 325156 3238 325194 3290
rect 325194 3238 325206 3290
rect 325206 3238 325212 3290
rect 325236 3238 325258 3290
rect 325258 3238 325270 3290
rect 325270 3238 325292 3290
rect 325316 3238 325322 3290
rect 325322 3238 325334 3290
rect 325334 3238 325372 3290
rect 324836 3236 324892 3238
rect 324916 3236 324972 3238
rect 324996 3236 325052 3238
rect 325076 3236 325132 3238
rect 325156 3236 325212 3238
rect 325236 3236 325292 3238
rect 325316 3236 325372 3238
rect 324836 2202 324892 2204
rect 324916 2202 324972 2204
rect 324996 2202 325052 2204
rect 325076 2202 325132 2204
rect 325156 2202 325212 2204
rect 325236 2202 325292 2204
rect 325316 2202 325372 2204
rect 324836 2150 324874 2202
rect 324874 2150 324886 2202
rect 324886 2150 324892 2202
rect 324916 2150 324938 2202
rect 324938 2150 324950 2202
rect 324950 2150 324972 2202
rect 324996 2150 325002 2202
rect 325002 2150 325014 2202
rect 325014 2150 325052 2202
rect 325076 2150 325078 2202
rect 325078 2150 325130 2202
rect 325130 2150 325132 2202
rect 325156 2150 325194 2202
rect 325194 2150 325206 2202
rect 325206 2150 325212 2202
rect 325236 2150 325258 2202
rect 325258 2150 325270 2202
rect 325270 2150 325292 2202
rect 325316 2150 325322 2202
rect 325322 2150 325334 2202
rect 325334 2150 325372 2202
rect 324836 2148 324892 2150
rect 324916 2148 324972 2150
rect 324996 2148 325052 2150
rect 325076 2148 325132 2150
rect 325156 2148 325212 2150
rect 325236 2148 325292 2150
rect 325316 2148 325372 2150
rect 342836 6010 342892 6012
rect 342916 6010 342972 6012
rect 342996 6010 343052 6012
rect 343076 6010 343132 6012
rect 343156 6010 343212 6012
rect 343236 6010 343292 6012
rect 343316 6010 343372 6012
rect 342836 5958 342874 6010
rect 342874 5958 342886 6010
rect 342886 5958 342892 6010
rect 342916 5958 342938 6010
rect 342938 5958 342950 6010
rect 342950 5958 342972 6010
rect 342996 5958 343002 6010
rect 343002 5958 343014 6010
rect 343014 5958 343052 6010
rect 343076 5958 343078 6010
rect 343078 5958 343130 6010
rect 343130 5958 343132 6010
rect 343156 5958 343194 6010
rect 343194 5958 343206 6010
rect 343206 5958 343212 6010
rect 343236 5958 343258 6010
rect 343258 5958 343270 6010
rect 343270 5958 343292 6010
rect 343316 5958 343322 6010
rect 343322 5958 343334 6010
rect 343334 5958 343372 6010
rect 342836 5956 342892 5958
rect 342916 5956 342972 5958
rect 342996 5956 343052 5958
rect 343076 5956 343132 5958
rect 343156 5956 343212 5958
rect 343236 5956 343292 5958
rect 343316 5956 343372 5958
rect 342836 4922 342892 4924
rect 342916 4922 342972 4924
rect 342996 4922 343052 4924
rect 343076 4922 343132 4924
rect 343156 4922 343212 4924
rect 343236 4922 343292 4924
rect 343316 4922 343372 4924
rect 342836 4870 342874 4922
rect 342874 4870 342886 4922
rect 342886 4870 342892 4922
rect 342916 4870 342938 4922
rect 342938 4870 342950 4922
rect 342950 4870 342972 4922
rect 342996 4870 343002 4922
rect 343002 4870 343014 4922
rect 343014 4870 343052 4922
rect 343076 4870 343078 4922
rect 343078 4870 343130 4922
rect 343130 4870 343132 4922
rect 343156 4870 343194 4922
rect 343194 4870 343206 4922
rect 343206 4870 343212 4922
rect 343236 4870 343258 4922
rect 343258 4870 343270 4922
rect 343270 4870 343292 4922
rect 343316 4870 343322 4922
rect 343322 4870 343334 4922
rect 343334 4870 343372 4922
rect 342836 4868 342892 4870
rect 342916 4868 342972 4870
rect 342996 4868 343052 4870
rect 343076 4868 343132 4870
rect 343156 4868 343212 4870
rect 343236 4868 343292 4870
rect 343316 4868 343372 4870
rect 342836 3834 342892 3836
rect 342916 3834 342972 3836
rect 342996 3834 343052 3836
rect 343076 3834 343132 3836
rect 343156 3834 343212 3836
rect 343236 3834 343292 3836
rect 343316 3834 343372 3836
rect 342836 3782 342874 3834
rect 342874 3782 342886 3834
rect 342886 3782 342892 3834
rect 342916 3782 342938 3834
rect 342938 3782 342950 3834
rect 342950 3782 342972 3834
rect 342996 3782 343002 3834
rect 343002 3782 343014 3834
rect 343014 3782 343052 3834
rect 343076 3782 343078 3834
rect 343078 3782 343130 3834
rect 343130 3782 343132 3834
rect 343156 3782 343194 3834
rect 343194 3782 343206 3834
rect 343206 3782 343212 3834
rect 343236 3782 343258 3834
rect 343258 3782 343270 3834
rect 343270 3782 343292 3834
rect 343316 3782 343322 3834
rect 343322 3782 343334 3834
rect 343334 3782 343372 3834
rect 342836 3780 342892 3782
rect 342916 3780 342972 3782
rect 342996 3780 343052 3782
rect 343076 3780 343132 3782
rect 343156 3780 343212 3782
rect 343236 3780 343292 3782
rect 343316 3780 343372 3782
rect 342836 2746 342892 2748
rect 342916 2746 342972 2748
rect 342996 2746 343052 2748
rect 343076 2746 343132 2748
rect 343156 2746 343212 2748
rect 343236 2746 343292 2748
rect 343316 2746 343372 2748
rect 342836 2694 342874 2746
rect 342874 2694 342886 2746
rect 342886 2694 342892 2746
rect 342916 2694 342938 2746
rect 342938 2694 342950 2746
rect 342950 2694 342972 2746
rect 342996 2694 343002 2746
rect 343002 2694 343014 2746
rect 343014 2694 343052 2746
rect 343076 2694 343078 2746
rect 343078 2694 343130 2746
rect 343130 2694 343132 2746
rect 343156 2694 343194 2746
rect 343194 2694 343206 2746
rect 343206 2694 343212 2746
rect 343236 2694 343258 2746
rect 343258 2694 343270 2746
rect 343270 2694 343292 2746
rect 343316 2694 343322 2746
rect 343322 2694 343334 2746
rect 343334 2694 343372 2746
rect 342836 2692 342892 2694
rect 342916 2692 342972 2694
rect 342996 2692 343052 2694
rect 343076 2692 343132 2694
rect 343156 2692 343212 2694
rect 343236 2692 343292 2694
rect 343316 2692 343372 2694
rect 360836 5466 360892 5468
rect 360916 5466 360972 5468
rect 360996 5466 361052 5468
rect 361076 5466 361132 5468
rect 361156 5466 361212 5468
rect 361236 5466 361292 5468
rect 361316 5466 361372 5468
rect 360836 5414 360874 5466
rect 360874 5414 360886 5466
rect 360886 5414 360892 5466
rect 360916 5414 360938 5466
rect 360938 5414 360950 5466
rect 360950 5414 360972 5466
rect 360996 5414 361002 5466
rect 361002 5414 361014 5466
rect 361014 5414 361052 5466
rect 361076 5414 361078 5466
rect 361078 5414 361130 5466
rect 361130 5414 361132 5466
rect 361156 5414 361194 5466
rect 361194 5414 361206 5466
rect 361206 5414 361212 5466
rect 361236 5414 361258 5466
rect 361258 5414 361270 5466
rect 361270 5414 361292 5466
rect 361316 5414 361322 5466
rect 361322 5414 361334 5466
rect 361334 5414 361372 5466
rect 360836 5412 360892 5414
rect 360916 5412 360972 5414
rect 360996 5412 361052 5414
rect 361076 5412 361132 5414
rect 361156 5412 361212 5414
rect 361236 5412 361292 5414
rect 361316 5412 361372 5414
rect 360836 4378 360892 4380
rect 360916 4378 360972 4380
rect 360996 4378 361052 4380
rect 361076 4378 361132 4380
rect 361156 4378 361212 4380
rect 361236 4378 361292 4380
rect 361316 4378 361372 4380
rect 360836 4326 360874 4378
rect 360874 4326 360886 4378
rect 360886 4326 360892 4378
rect 360916 4326 360938 4378
rect 360938 4326 360950 4378
rect 360950 4326 360972 4378
rect 360996 4326 361002 4378
rect 361002 4326 361014 4378
rect 361014 4326 361052 4378
rect 361076 4326 361078 4378
rect 361078 4326 361130 4378
rect 361130 4326 361132 4378
rect 361156 4326 361194 4378
rect 361194 4326 361206 4378
rect 361206 4326 361212 4378
rect 361236 4326 361258 4378
rect 361258 4326 361270 4378
rect 361270 4326 361292 4378
rect 361316 4326 361322 4378
rect 361322 4326 361334 4378
rect 361334 4326 361372 4378
rect 360836 4324 360892 4326
rect 360916 4324 360972 4326
rect 360996 4324 361052 4326
rect 361076 4324 361132 4326
rect 361156 4324 361212 4326
rect 361236 4324 361292 4326
rect 361316 4324 361372 4326
rect 360836 3290 360892 3292
rect 360916 3290 360972 3292
rect 360996 3290 361052 3292
rect 361076 3290 361132 3292
rect 361156 3290 361212 3292
rect 361236 3290 361292 3292
rect 361316 3290 361372 3292
rect 360836 3238 360874 3290
rect 360874 3238 360886 3290
rect 360886 3238 360892 3290
rect 360916 3238 360938 3290
rect 360938 3238 360950 3290
rect 360950 3238 360972 3290
rect 360996 3238 361002 3290
rect 361002 3238 361014 3290
rect 361014 3238 361052 3290
rect 361076 3238 361078 3290
rect 361078 3238 361130 3290
rect 361130 3238 361132 3290
rect 361156 3238 361194 3290
rect 361194 3238 361206 3290
rect 361206 3238 361212 3290
rect 361236 3238 361258 3290
rect 361258 3238 361270 3290
rect 361270 3238 361292 3290
rect 361316 3238 361322 3290
rect 361322 3238 361334 3290
rect 361334 3238 361372 3290
rect 360836 3236 360892 3238
rect 360916 3236 360972 3238
rect 360996 3236 361052 3238
rect 361076 3236 361132 3238
rect 361156 3236 361212 3238
rect 361236 3236 361292 3238
rect 361316 3236 361372 3238
rect 360836 2202 360892 2204
rect 360916 2202 360972 2204
rect 360996 2202 361052 2204
rect 361076 2202 361132 2204
rect 361156 2202 361212 2204
rect 361236 2202 361292 2204
rect 361316 2202 361372 2204
rect 360836 2150 360874 2202
rect 360874 2150 360886 2202
rect 360886 2150 360892 2202
rect 360916 2150 360938 2202
rect 360938 2150 360950 2202
rect 360950 2150 360972 2202
rect 360996 2150 361002 2202
rect 361002 2150 361014 2202
rect 361014 2150 361052 2202
rect 361076 2150 361078 2202
rect 361078 2150 361130 2202
rect 361130 2150 361132 2202
rect 361156 2150 361194 2202
rect 361194 2150 361206 2202
rect 361206 2150 361212 2202
rect 361236 2150 361258 2202
rect 361258 2150 361270 2202
rect 361270 2150 361292 2202
rect 361316 2150 361322 2202
rect 361322 2150 361334 2202
rect 361334 2150 361372 2202
rect 360836 2148 360892 2150
rect 360916 2148 360972 2150
rect 360996 2148 361052 2150
rect 361076 2148 361132 2150
rect 361156 2148 361212 2150
rect 361236 2148 361292 2150
rect 361316 2148 361372 2150
rect 378836 6010 378892 6012
rect 378916 6010 378972 6012
rect 378996 6010 379052 6012
rect 379076 6010 379132 6012
rect 379156 6010 379212 6012
rect 379236 6010 379292 6012
rect 379316 6010 379372 6012
rect 378836 5958 378874 6010
rect 378874 5958 378886 6010
rect 378886 5958 378892 6010
rect 378916 5958 378938 6010
rect 378938 5958 378950 6010
rect 378950 5958 378972 6010
rect 378996 5958 379002 6010
rect 379002 5958 379014 6010
rect 379014 5958 379052 6010
rect 379076 5958 379078 6010
rect 379078 5958 379130 6010
rect 379130 5958 379132 6010
rect 379156 5958 379194 6010
rect 379194 5958 379206 6010
rect 379206 5958 379212 6010
rect 379236 5958 379258 6010
rect 379258 5958 379270 6010
rect 379270 5958 379292 6010
rect 379316 5958 379322 6010
rect 379322 5958 379334 6010
rect 379334 5958 379372 6010
rect 378836 5956 378892 5958
rect 378916 5956 378972 5958
rect 378996 5956 379052 5958
rect 379076 5956 379132 5958
rect 379156 5956 379212 5958
rect 379236 5956 379292 5958
rect 379316 5956 379372 5958
rect 378836 4922 378892 4924
rect 378916 4922 378972 4924
rect 378996 4922 379052 4924
rect 379076 4922 379132 4924
rect 379156 4922 379212 4924
rect 379236 4922 379292 4924
rect 379316 4922 379372 4924
rect 378836 4870 378874 4922
rect 378874 4870 378886 4922
rect 378886 4870 378892 4922
rect 378916 4870 378938 4922
rect 378938 4870 378950 4922
rect 378950 4870 378972 4922
rect 378996 4870 379002 4922
rect 379002 4870 379014 4922
rect 379014 4870 379052 4922
rect 379076 4870 379078 4922
rect 379078 4870 379130 4922
rect 379130 4870 379132 4922
rect 379156 4870 379194 4922
rect 379194 4870 379206 4922
rect 379206 4870 379212 4922
rect 379236 4870 379258 4922
rect 379258 4870 379270 4922
rect 379270 4870 379292 4922
rect 379316 4870 379322 4922
rect 379322 4870 379334 4922
rect 379334 4870 379372 4922
rect 378836 4868 378892 4870
rect 378916 4868 378972 4870
rect 378996 4868 379052 4870
rect 379076 4868 379132 4870
rect 379156 4868 379212 4870
rect 379236 4868 379292 4870
rect 379316 4868 379372 4870
rect 378836 3834 378892 3836
rect 378916 3834 378972 3836
rect 378996 3834 379052 3836
rect 379076 3834 379132 3836
rect 379156 3834 379212 3836
rect 379236 3834 379292 3836
rect 379316 3834 379372 3836
rect 378836 3782 378874 3834
rect 378874 3782 378886 3834
rect 378886 3782 378892 3834
rect 378916 3782 378938 3834
rect 378938 3782 378950 3834
rect 378950 3782 378972 3834
rect 378996 3782 379002 3834
rect 379002 3782 379014 3834
rect 379014 3782 379052 3834
rect 379076 3782 379078 3834
rect 379078 3782 379130 3834
rect 379130 3782 379132 3834
rect 379156 3782 379194 3834
rect 379194 3782 379206 3834
rect 379206 3782 379212 3834
rect 379236 3782 379258 3834
rect 379258 3782 379270 3834
rect 379270 3782 379292 3834
rect 379316 3782 379322 3834
rect 379322 3782 379334 3834
rect 379334 3782 379372 3834
rect 378836 3780 378892 3782
rect 378916 3780 378972 3782
rect 378996 3780 379052 3782
rect 379076 3780 379132 3782
rect 379156 3780 379212 3782
rect 379236 3780 379292 3782
rect 379316 3780 379372 3782
rect 378836 2746 378892 2748
rect 378916 2746 378972 2748
rect 378996 2746 379052 2748
rect 379076 2746 379132 2748
rect 379156 2746 379212 2748
rect 379236 2746 379292 2748
rect 379316 2746 379372 2748
rect 378836 2694 378874 2746
rect 378874 2694 378886 2746
rect 378886 2694 378892 2746
rect 378916 2694 378938 2746
rect 378938 2694 378950 2746
rect 378950 2694 378972 2746
rect 378996 2694 379002 2746
rect 379002 2694 379014 2746
rect 379014 2694 379052 2746
rect 379076 2694 379078 2746
rect 379078 2694 379130 2746
rect 379130 2694 379132 2746
rect 379156 2694 379194 2746
rect 379194 2694 379206 2746
rect 379206 2694 379212 2746
rect 379236 2694 379258 2746
rect 379258 2694 379270 2746
rect 379270 2694 379292 2746
rect 379316 2694 379322 2746
rect 379322 2694 379334 2746
rect 379334 2694 379372 2746
rect 378836 2692 378892 2694
rect 378916 2692 378972 2694
rect 378996 2692 379052 2694
rect 379076 2692 379132 2694
rect 379156 2692 379212 2694
rect 379236 2692 379292 2694
rect 379316 2692 379372 2694
rect 396836 5466 396892 5468
rect 396916 5466 396972 5468
rect 396996 5466 397052 5468
rect 397076 5466 397132 5468
rect 397156 5466 397212 5468
rect 397236 5466 397292 5468
rect 397316 5466 397372 5468
rect 396836 5414 396874 5466
rect 396874 5414 396886 5466
rect 396886 5414 396892 5466
rect 396916 5414 396938 5466
rect 396938 5414 396950 5466
rect 396950 5414 396972 5466
rect 396996 5414 397002 5466
rect 397002 5414 397014 5466
rect 397014 5414 397052 5466
rect 397076 5414 397078 5466
rect 397078 5414 397130 5466
rect 397130 5414 397132 5466
rect 397156 5414 397194 5466
rect 397194 5414 397206 5466
rect 397206 5414 397212 5466
rect 397236 5414 397258 5466
rect 397258 5414 397270 5466
rect 397270 5414 397292 5466
rect 397316 5414 397322 5466
rect 397322 5414 397334 5466
rect 397334 5414 397372 5466
rect 396836 5412 396892 5414
rect 396916 5412 396972 5414
rect 396996 5412 397052 5414
rect 397076 5412 397132 5414
rect 397156 5412 397212 5414
rect 397236 5412 397292 5414
rect 397316 5412 397372 5414
rect 396836 4378 396892 4380
rect 396916 4378 396972 4380
rect 396996 4378 397052 4380
rect 397076 4378 397132 4380
rect 397156 4378 397212 4380
rect 397236 4378 397292 4380
rect 397316 4378 397372 4380
rect 396836 4326 396874 4378
rect 396874 4326 396886 4378
rect 396886 4326 396892 4378
rect 396916 4326 396938 4378
rect 396938 4326 396950 4378
rect 396950 4326 396972 4378
rect 396996 4326 397002 4378
rect 397002 4326 397014 4378
rect 397014 4326 397052 4378
rect 397076 4326 397078 4378
rect 397078 4326 397130 4378
rect 397130 4326 397132 4378
rect 397156 4326 397194 4378
rect 397194 4326 397206 4378
rect 397206 4326 397212 4378
rect 397236 4326 397258 4378
rect 397258 4326 397270 4378
rect 397270 4326 397292 4378
rect 397316 4326 397322 4378
rect 397322 4326 397334 4378
rect 397334 4326 397372 4378
rect 396836 4324 396892 4326
rect 396916 4324 396972 4326
rect 396996 4324 397052 4326
rect 397076 4324 397132 4326
rect 397156 4324 397212 4326
rect 397236 4324 397292 4326
rect 397316 4324 397372 4326
rect 396836 3290 396892 3292
rect 396916 3290 396972 3292
rect 396996 3290 397052 3292
rect 397076 3290 397132 3292
rect 397156 3290 397212 3292
rect 397236 3290 397292 3292
rect 397316 3290 397372 3292
rect 396836 3238 396874 3290
rect 396874 3238 396886 3290
rect 396886 3238 396892 3290
rect 396916 3238 396938 3290
rect 396938 3238 396950 3290
rect 396950 3238 396972 3290
rect 396996 3238 397002 3290
rect 397002 3238 397014 3290
rect 397014 3238 397052 3290
rect 397076 3238 397078 3290
rect 397078 3238 397130 3290
rect 397130 3238 397132 3290
rect 397156 3238 397194 3290
rect 397194 3238 397206 3290
rect 397206 3238 397212 3290
rect 397236 3238 397258 3290
rect 397258 3238 397270 3290
rect 397270 3238 397292 3290
rect 397316 3238 397322 3290
rect 397322 3238 397334 3290
rect 397334 3238 397372 3290
rect 396836 3236 396892 3238
rect 396916 3236 396972 3238
rect 396996 3236 397052 3238
rect 397076 3236 397132 3238
rect 397156 3236 397212 3238
rect 397236 3236 397292 3238
rect 397316 3236 397372 3238
rect 396836 2202 396892 2204
rect 396916 2202 396972 2204
rect 396996 2202 397052 2204
rect 397076 2202 397132 2204
rect 397156 2202 397212 2204
rect 397236 2202 397292 2204
rect 397316 2202 397372 2204
rect 396836 2150 396874 2202
rect 396874 2150 396886 2202
rect 396886 2150 396892 2202
rect 396916 2150 396938 2202
rect 396938 2150 396950 2202
rect 396950 2150 396972 2202
rect 396996 2150 397002 2202
rect 397002 2150 397014 2202
rect 397014 2150 397052 2202
rect 397076 2150 397078 2202
rect 397078 2150 397130 2202
rect 397130 2150 397132 2202
rect 397156 2150 397194 2202
rect 397194 2150 397206 2202
rect 397206 2150 397212 2202
rect 397236 2150 397258 2202
rect 397258 2150 397270 2202
rect 397270 2150 397292 2202
rect 397316 2150 397322 2202
rect 397322 2150 397334 2202
rect 397334 2150 397372 2202
rect 396836 2148 396892 2150
rect 396916 2148 396972 2150
rect 396996 2148 397052 2150
rect 397076 2148 397132 2150
rect 397156 2148 397212 2150
rect 397236 2148 397292 2150
rect 397316 2148 397372 2150
rect 414836 6010 414892 6012
rect 414916 6010 414972 6012
rect 414996 6010 415052 6012
rect 415076 6010 415132 6012
rect 415156 6010 415212 6012
rect 415236 6010 415292 6012
rect 415316 6010 415372 6012
rect 414836 5958 414874 6010
rect 414874 5958 414886 6010
rect 414886 5958 414892 6010
rect 414916 5958 414938 6010
rect 414938 5958 414950 6010
rect 414950 5958 414972 6010
rect 414996 5958 415002 6010
rect 415002 5958 415014 6010
rect 415014 5958 415052 6010
rect 415076 5958 415078 6010
rect 415078 5958 415130 6010
rect 415130 5958 415132 6010
rect 415156 5958 415194 6010
rect 415194 5958 415206 6010
rect 415206 5958 415212 6010
rect 415236 5958 415258 6010
rect 415258 5958 415270 6010
rect 415270 5958 415292 6010
rect 415316 5958 415322 6010
rect 415322 5958 415334 6010
rect 415334 5958 415372 6010
rect 414836 5956 414892 5958
rect 414916 5956 414972 5958
rect 414996 5956 415052 5958
rect 415076 5956 415132 5958
rect 415156 5956 415212 5958
rect 415236 5956 415292 5958
rect 415316 5956 415372 5958
rect 414836 4922 414892 4924
rect 414916 4922 414972 4924
rect 414996 4922 415052 4924
rect 415076 4922 415132 4924
rect 415156 4922 415212 4924
rect 415236 4922 415292 4924
rect 415316 4922 415372 4924
rect 414836 4870 414874 4922
rect 414874 4870 414886 4922
rect 414886 4870 414892 4922
rect 414916 4870 414938 4922
rect 414938 4870 414950 4922
rect 414950 4870 414972 4922
rect 414996 4870 415002 4922
rect 415002 4870 415014 4922
rect 415014 4870 415052 4922
rect 415076 4870 415078 4922
rect 415078 4870 415130 4922
rect 415130 4870 415132 4922
rect 415156 4870 415194 4922
rect 415194 4870 415206 4922
rect 415206 4870 415212 4922
rect 415236 4870 415258 4922
rect 415258 4870 415270 4922
rect 415270 4870 415292 4922
rect 415316 4870 415322 4922
rect 415322 4870 415334 4922
rect 415334 4870 415372 4922
rect 414836 4868 414892 4870
rect 414916 4868 414972 4870
rect 414996 4868 415052 4870
rect 415076 4868 415132 4870
rect 415156 4868 415212 4870
rect 415236 4868 415292 4870
rect 415316 4868 415372 4870
rect 414836 3834 414892 3836
rect 414916 3834 414972 3836
rect 414996 3834 415052 3836
rect 415076 3834 415132 3836
rect 415156 3834 415212 3836
rect 415236 3834 415292 3836
rect 415316 3834 415372 3836
rect 414836 3782 414874 3834
rect 414874 3782 414886 3834
rect 414886 3782 414892 3834
rect 414916 3782 414938 3834
rect 414938 3782 414950 3834
rect 414950 3782 414972 3834
rect 414996 3782 415002 3834
rect 415002 3782 415014 3834
rect 415014 3782 415052 3834
rect 415076 3782 415078 3834
rect 415078 3782 415130 3834
rect 415130 3782 415132 3834
rect 415156 3782 415194 3834
rect 415194 3782 415206 3834
rect 415206 3782 415212 3834
rect 415236 3782 415258 3834
rect 415258 3782 415270 3834
rect 415270 3782 415292 3834
rect 415316 3782 415322 3834
rect 415322 3782 415334 3834
rect 415334 3782 415372 3834
rect 414836 3780 414892 3782
rect 414916 3780 414972 3782
rect 414996 3780 415052 3782
rect 415076 3780 415132 3782
rect 415156 3780 415212 3782
rect 415236 3780 415292 3782
rect 415316 3780 415372 3782
rect 414836 2746 414892 2748
rect 414916 2746 414972 2748
rect 414996 2746 415052 2748
rect 415076 2746 415132 2748
rect 415156 2746 415212 2748
rect 415236 2746 415292 2748
rect 415316 2746 415372 2748
rect 414836 2694 414874 2746
rect 414874 2694 414886 2746
rect 414886 2694 414892 2746
rect 414916 2694 414938 2746
rect 414938 2694 414950 2746
rect 414950 2694 414972 2746
rect 414996 2694 415002 2746
rect 415002 2694 415014 2746
rect 415014 2694 415052 2746
rect 415076 2694 415078 2746
rect 415078 2694 415130 2746
rect 415130 2694 415132 2746
rect 415156 2694 415194 2746
rect 415194 2694 415206 2746
rect 415206 2694 415212 2746
rect 415236 2694 415258 2746
rect 415258 2694 415270 2746
rect 415270 2694 415292 2746
rect 415316 2694 415322 2746
rect 415322 2694 415334 2746
rect 415334 2694 415372 2746
rect 414836 2692 414892 2694
rect 414916 2692 414972 2694
rect 414996 2692 415052 2694
rect 415076 2692 415132 2694
rect 415156 2692 415212 2694
rect 415236 2692 415292 2694
rect 415316 2692 415372 2694
rect 432836 5466 432892 5468
rect 432916 5466 432972 5468
rect 432996 5466 433052 5468
rect 433076 5466 433132 5468
rect 433156 5466 433212 5468
rect 433236 5466 433292 5468
rect 433316 5466 433372 5468
rect 432836 5414 432874 5466
rect 432874 5414 432886 5466
rect 432886 5414 432892 5466
rect 432916 5414 432938 5466
rect 432938 5414 432950 5466
rect 432950 5414 432972 5466
rect 432996 5414 433002 5466
rect 433002 5414 433014 5466
rect 433014 5414 433052 5466
rect 433076 5414 433078 5466
rect 433078 5414 433130 5466
rect 433130 5414 433132 5466
rect 433156 5414 433194 5466
rect 433194 5414 433206 5466
rect 433206 5414 433212 5466
rect 433236 5414 433258 5466
rect 433258 5414 433270 5466
rect 433270 5414 433292 5466
rect 433316 5414 433322 5466
rect 433322 5414 433334 5466
rect 433334 5414 433372 5466
rect 432836 5412 432892 5414
rect 432916 5412 432972 5414
rect 432996 5412 433052 5414
rect 433076 5412 433132 5414
rect 433156 5412 433212 5414
rect 433236 5412 433292 5414
rect 433316 5412 433372 5414
rect 432836 4378 432892 4380
rect 432916 4378 432972 4380
rect 432996 4378 433052 4380
rect 433076 4378 433132 4380
rect 433156 4378 433212 4380
rect 433236 4378 433292 4380
rect 433316 4378 433372 4380
rect 432836 4326 432874 4378
rect 432874 4326 432886 4378
rect 432886 4326 432892 4378
rect 432916 4326 432938 4378
rect 432938 4326 432950 4378
rect 432950 4326 432972 4378
rect 432996 4326 433002 4378
rect 433002 4326 433014 4378
rect 433014 4326 433052 4378
rect 433076 4326 433078 4378
rect 433078 4326 433130 4378
rect 433130 4326 433132 4378
rect 433156 4326 433194 4378
rect 433194 4326 433206 4378
rect 433206 4326 433212 4378
rect 433236 4326 433258 4378
rect 433258 4326 433270 4378
rect 433270 4326 433292 4378
rect 433316 4326 433322 4378
rect 433322 4326 433334 4378
rect 433334 4326 433372 4378
rect 432836 4324 432892 4326
rect 432916 4324 432972 4326
rect 432996 4324 433052 4326
rect 433076 4324 433132 4326
rect 433156 4324 433212 4326
rect 433236 4324 433292 4326
rect 433316 4324 433372 4326
rect 432836 3290 432892 3292
rect 432916 3290 432972 3292
rect 432996 3290 433052 3292
rect 433076 3290 433132 3292
rect 433156 3290 433212 3292
rect 433236 3290 433292 3292
rect 433316 3290 433372 3292
rect 432836 3238 432874 3290
rect 432874 3238 432886 3290
rect 432886 3238 432892 3290
rect 432916 3238 432938 3290
rect 432938 3238 432950 3290
rect 432950 3238 432972 3290
rect 432996 3238 433002 3290
rect 433002 3238 433014 3290
rect 433014 3238 433052 3290
rect 433076 3238 433078 3290
rect 433078 3238 433130 3290
rect 433130 3238 433132 3290
rect 433156 3238 433194 3290
rect 433194 3238 433206 3290
rect 433206 3238 433212 3290
rect 433236 3238 433258 3290
rect 433258 3238 433270 3290
rect 433270 3238 433292 3290
rect 433316 3238 433322 3290
rect 433322 3238 433334 3290
rect 433334 3238 433372 3290
rect 432836 3236 432892 3238
rect 432916 3236 432972 3238
rect 432996 3236 433052 3238
rect 433076 3236 433132 3238
rect 433156 3236 433212 3238
rect 433236 3236 433292 3238
rect 433316 3236 433372 3238
rect 432836 2202 432892 2204
rect 432916 2202 432972 2204
rect 432996 2202 433052 2204
rect 433076 2202 433132 2204
rect 433156 2202 433212 2204
rect 433236 2202 433292 2204
rect 433316 2202 433372 2204
rect 432836 2150 432874 2202
rect 432874 2150 432886 2202
rect 432886 2150 432892 2202
rect 432916 2150 432938 2202
rect 432938 2150 432950 2202
rect 432950 2150 432972 2202
rect 432996 2150 433002 2202
rect 433002 2150 433014 2202
rect 433014 2150 433052 2202
rect 433076 2150 433078 2202
rect 433078 2150 433130 2202
rect 433130 2150 433132 2202
rect 433156 2150 433194 2202
rect 433194 2150 433206 2202
rect 433206 2150 433212 2202
rect 433236 2150 433258 2202
rect 433258 2150 433270 2202
rect 433270 2150 433292 2202
rect 433316 2150 433322 2202
rect 433322 2150 433334 2202
rect 433334 2150 433372 2202
rect 432836 2148 432892 2150
rect 432916 2148 432972 2150
rect 432996 2148 433052 2150
rect 433076 2148 433132 2150
rect 433156 2148 433212 2150
rect 433236 2148 433292 2150
rect 433316 2148 433372 2150
rect 450836 6010 450892 6012
rect 450916 6010 450972 6012
rect 450996 6010 451052 6012
rect 451076 6010 451132 6012
rect 451156 6010 451212 6012
rect 451236 6010 451292 6012
rect 451316 6010 451372 6012
rect 450836 5958 450874 6010
rect 450874 5958 450886 6010
rect 450886 5958 450892 6010
rect 450916 5958 450938 6010
rect 450938 5958 450950 6010
rect 450950 5958 450972 6010
rect 450996 5958 451002 6010
rect 451002 5958 451014 6010
rect 451014 5958 451052 6010
rect 451076 5958 451078 6010
rect 451078 5958 451130 6010
rect 451130 5958 451132 6010
rect 451156 5958 451194 6010
rect 451194 5958 451206 6010
rect 451206 5958 451212 6010
rect 451236 5958 451258 6010
rect 451258 5958 451270 6010
rect 451270 5958 451292 6010
rect 451316 5958 451322 6010
rect 451322 5958 451334 6010
rect 451334 5958 451372 6010
rect 450836 5956 450892 5958
rect 450916 5956 450972 5958
rect 450996 5956 451052 5958
rect 451076 5956 451132 5958
rect 451156 5956 451212 5958
rect 451236 5956 451292 5958
rect 451316 5956 451372 5958
rect 450836 4922 450892 4924
rect 450916 4922 450972 4924
rect 450996 4922 451052 4924
rect 451076 4922 451132 4924
rect 451156 4922 451212 4924
rect 451236 4922 451292 4924
rect 451316 4922 451372 4924
rect 450836 4870 450874 4922
rect 450874 4870 450886 4922
rect 450886 4870 450892 4922
rect 450916 4870 450938 4922
rect 450938 4870 450950 4922
rect 450950 4870 450972 4922
rect 450996 4870 451002 4922
rect 451002 4870 451014 4922
rect 451014 4870 451052 4922
rect 451076 4870 451078 4922
rect 451078 4870 451130 4922
rect 451130 4870 451132 4922
rect 451156 4870 451194 4922
rect 451194 4870 451206 4922
rect 451206 4870 451212 4922
rect 451236 4870 451258 4922
rect 451258 4870 451270 4922
rect 451270 4870 451292 4922
rect 451316 4870 451322 4922
rect 451322 4870 451334 4922
rect 451334 4870 451372 4922
rect 450836 4868 450892 4870
rect 450916 4868 450972 4870
rect 450996 4868 451052 4870
rect 451076 4868 451132 4870
rect 451156 4868 451212 4870
rect 451236 4868 451292 4870
rect 451316 4868 451372 4870
rect 450836 3834 450892 3836
rect 450916 3834 450972 3836
rect 450996 3834 451052 3836
rect 451076 3834 451132 3836
rect 451156 3834 451212 3836
rect 451236 3834 451292 3836
rect 451316 3834 451372 3836
rect 450836 3782 450874 3834
rect 450874 3782 450886 3834
rect 450886 3782 450892 3834
rect 450916 3782 450938 3834
rect 450938 3782 450950 3834
rect 450950 3782 450972 3834
rect 450996 3782 451002 3834
rect 451002 3782 451014 3834
rect 451014 3782 451052 3834
rect 451076 3782 451078 3834
rect 451078 3782 451130 3834
rect 451130 3782 451132 3834
rect 451156 3782 451194 3834
rect 451194 3782 451206 3834
rect 451206 3782 451212 3834
rect 451236 3782 451258 3834
rect 451258 3782 451270 3834
rect 451270 3782 451292 3834
rect 451316 3782 451322 3834
rect 451322 3782 451334 3834
rect 451334 3782 451372 3834
rect 450836 3780 450892 3782
rect 450916 3780 450972 3782
rect 450996 3780 451052 3782
rect 451076 3780 451132 3782
rect 451156 3780 451212 3782
rect 451236 3780 451292 3782
rect 451316 3780 451372 3782
rect 450836 2746 450892 2748
rect 450916 2746 450972 2748
rect 450996 2746 451052 2748
rect 451076 2746 451132 2748
rect 451156 2746 451212 2748
rect 451236 2746 451292 2748
rect 451316 2746 451372 2748
rect 450836 2694 450874 2746
rect 450874 2694 450886 2746
rect 450886 2694 450892 2746
rect 450916 2694 450938 2746
rect 450938 2694 450950 2746
rect 450950 2694 450972 2746
rect 450996 2694 451002 2746
rect 451002 2694 451014 2746
rect 451014 2694 451052 2746
rect 451076 2694 451078 2746
rect 451078 2694 451130 2746
rect 451130 2694 451132 2746
rect 451156 2694 451194 2746
rect 451194 2694 451206 2746
rect 451206 2694 451212 2746
rect 451236 2694 451258 2746
rect 451258 2694 451270 2746
rect 451270 2694 451292 2746
rect 451316 2694 451322 2746
rect 451322 2694 451334 2746
rect 451334 2694 451372 2746
rect 450836 2692 450892 2694
rect 450916 2692 450972 2694
rect 450996 2692 451052 2694
rect 451076 2692 451132 2694
rect 451156 2692 451212 2694
rect 451236 2692 451292 2694
rect 451316 2692 451372 2694
rect 468836 5466 468892 5468
rect 468916 5466 468972 5468
rect 468996 5466 469052 5468
rect 469076 5466 469132 5468
rect 469156 5466 469212 5468
rect 469236 5466 469292 5468
rect 469316 5466 469372 5468
rect 468836 5414 468874 5466
rect 468874 5414 468886 5466
rect 468886 5414 468892 5466
rect 468916 5414 468938 5466
rect 468938 5414 468950 5466
rect 468950 5414 468972 5466
rect 468996 5414 469002 5466
rect 469002 5414 469014 5466
rect 469014 5414 469052 5466
rect 469076 5414 469078 5466
rect 469078 5414 469130 5466
rect 469130 5414 469132 5466
rect 469156 5414 469194 5466
rect 469194 5414 469206 5466
rect 469206 5414 469212 5466
rect 469236 5414 469258 5466
rect 469258 5414 469270 5466
rect 469270 5414 469292 5466
rect 469316 5414 469322 5466
rect 469322 5414 469334 5466
rect 469334 5414 469372 5466
rect 468836 5412 468892 5414
rect 468916 5412 468972 5414
rect 468996 5412 469052 5414
rect 469076 5412 469132 5414
rect 469156 5412 469212 5414
rect 469236 5412 469292 5414
rect 469316 5412 469372 5414
rect 468836 4378 468892 4380
rect 468916 4378 468972 4380
rect 468996 4378 469052 4380
rect 469076 4378 469132 4380
rect 469156 4378 469212 4380
rect 469236 4378 469292 4380
rect 469316 4378 469372 4380
rect 468836 4326 468874 4378
rect 468874 4326 468886 4378
rect 468886 4326 468892 4378
rect 468916 4326 468938 4378
rect 468938 4326 468950 4378
rect 468950 4326 468972 4378
rect 468996 4326 469002 4378
rect 469002 4326 469014 4378
rect 469014 4326 469052 4378
rect 469076 4326 469078 4378
rect 469078 4326 469130 4378
rect 469130 4326 469132 4378
rect 469156 4326 469194 4378
rect 469194 4326 469206 4378
rect 469206 4326 469212 4378
rect 469236 4326 469258 4378
rect 469258 4326 469270 4378
rect 469270 4326 469292 4378
rect 469316 4326 469322 4378
rect 469322 4326 469334 4378
rect 469334 4326 469372 4378
rect 468836 4324 468892 4326
rect 468916 4324 468972 4326
rect 468996 4324 469052 4326
rect 469076 4324 469132 4326
rect 469156 4324 469212 4326
rect 469236 4324 469292 4326
rect 469316 4324 469372 4326
rect 468836 3290 468892 3292
rect 468916 3290 468972 3292
rect 468996 3290 469052 3292
rect 469076 3290 469132 3292
rect 469156 3290 469212 3292
rect 469236 3290 469292 3292
rect 469316 3290 469372 3292
rect 468836 3238 468874 3290
rect 468874 3238 468886 3290
rect 468886 3238 468892 3290
rect 468916 3238 468938 3290
rect 468938 3238 468950 3290
rect 468950 3238 468972 3290
rect 468996 3238 469002 3290
rect 469002 3238 469014 3290
rect 469014 3238 469052 3290
rect 469076 3238 469078 3290
rect 469078 3238 469130 3290
rect 469130 3238 469132 3290
rect 469156 3238 469194 3290
rect 469194 3238 469206 3290
rect 469206 3238 469212 3290
rect 469236 3238 469258 3290
rect 469258 3238 469270 3290
rect 469270 3238 469292 3290
rect 469316 3238 469322 3290
rect 469322 3238 469334 3290
rect 469334 3238 469372 3290
rect 468836 3236 468892 3238
rect 468916 3236 468972 3238
rect 468996 3236 469052 3238
rect 469076 3236 469132 3238
rect 469156 3236 469212 3238
rect 469236 3236 469292 3238
rect 469316 3236 469372 3238
rect 468836 2202 468892 2204
rect 468916 2202 468972 2204
rect 468996 2202 469052 2204
rect 469076 2202 469132 2204
rect 469156 2202 469212 2204
rect 469236 2202 469292 2204
rect 469316 2202 469372 2204
rect 468836 2150 468874 2202
rect 468874 2150 468886 2202
rect 468886 2150 468892 2202
rect 468916 2150 468938 2202
rect 468938 2150 468950 2202
rect 468950 2150 468972 2202
rect 468996 2150 469002 2202
rect 469002 2150 469014 2202
rect 469014 2150 469052 2202
rect 469076 2150 469078 2202
rect 469078 2150 469130 2202
rect 469130 2150 469132 2202
rect 469156 2150 469194 2202
rect 469194 2150 469206 2202
rect 469206 2150 469212 2202
rect 469236 2150 469258 2202
rect 469258 2150 469270 2202
rect 469270 2150 469292 2202
rect 469316 2150 469322 2202
rect 469322 2150 469334 2202
rect 469334 2150 469372 2202
rect 468836 2148 468892 2150
rect 468916 2148 468972 2150
rect 468996 2148 469052 2150
rect 469076 2148 469132 2150
rect 469156 2148 469212 2150
rect 469236 2148 469292 2150
rect 469316 2148 469372 2150
rect 486836 6010 486892 6012
rect 486916 6010 486972 6012
rect 486996 6010 487052 6012
rect 487076 6010 487132 6012
rect 487156 6010 487212 6012
rect 487236 6010 487292 6012
rect 487316 6010 487372 6012
rect 486836 5958 486874 6010
rect 486874 5958 486886 6010
rect 486886 5958 486892 6010
rect 486916 5958 486938 6010
rect 486938 5958 486950 6010
rect 486950 5958 486972 6010
rect 486996 5958 487002 6010
rect 487002 5958 487014 6010
rect 487014 5958 487052 6010
rect 487076 5958 487078 6010
rect 487078 5958 487130 6010
rect 487130 5958 487132 6010
rect 487156 5958 487194 6010
rect 487194 5958 487206 6010
rect 487206 5958 487212 6010
rect 487236 5958 487258 6010
rect 487258 5958 487270 6010
rect 487270 5958 487292 6010
rect 487316 5958 487322 6010
rect 487322 5958 487334 6010
rect 487334 5958 487372 6010
rect 486836 5956 486892 5958
rect 486916 5956 486972 5958
rect 486996 5956 487052 5958
rect 487076 5956 487132 5958
rect 487156 5956 487212 5958
rect 487236 5956 487292 5958
rect 487316 5956 487372 5958
rect 486836 4922 486892 4924
rect 486916 4922 486972 4924
rect 486996 4922 487052 4924
rect 487076 4922 487132 4924
rect 487156 4922 487212 4924
rect 487236 4922 487292 4924
rect 487316 4922 487372 4924
rect 486836 4870 486874 4922
rect 486874 4870 486886 4922
rect 486886 4870 486892 4922
rect 486916 4870 486938 4922
rect 486938 4870 486950 4922
rect 486950 4870 486972 4922
rect 486996 4870 487002 4922
rect 487002 4870 487014 4922
rect 487014 4870 487052 4922
rect 487076 4870 487078 4922
rect 487078 4870 487130 4922
rect 487130 4870 487132 4922
rect 487156 4870 487194 4922
rect 487194 4870 487206 4922
rect 487206 4870 487212 4922
rect 487236 4870 487258 4922
rect 487258 4870 487270 4922
rect 487270 4870 487292 4922
rect 487316 4870 487322 4922
rect 487322 4870 487334 4922
rect 487334 4870 487372 4922
rect 486836 4868 486892 4870
rect 486916 4868 486972 4870
rect 486996 4868 487052 4870
rect 487076 4868 487132 4870
rect 487156 4868 487212 4870
rect 487236 4868 487292 4870
rect 487316 4868 487372 4870
rect 486836 3834 486892 3836
rect 486916 3834 486972 3836
rect 486996 3834 487052 3836
rect 487076 3834 487132 3836
rect 487156 3834 487212 3836
rect 487236 3834 487292 3836
rect 487316 3834 487372 3836
rect 486836 3782 486874 3834
rect 486874 3782 486886 3834
rect 486886 3782 486892 3834
rect 486916 3782 486938 3834
rect 486938 3782 486950 3834
rect 486950 3782 486972 3834
rect 486996 3782 487002 3834
rect 487002 3782 487014 3834
rect 487014 3782 487052 3834
rect 487076 3782 487078 3834
rect 487078 3782 487130 3834
rect 487130 3782 487132 3834
rect 487156 3782 487194 3834
rect 487194 3782 487206 3834
rect 487206 3782 487212 3834
rect 487236 3782 487258 3834
rect 487258 3782 487270 3834
rect 487270 3782 487292 3834
rect 487316 3782 487322 3834
rect 487322 3782 487334 3834
rect 487334 3782 487372 3834
rect 486836 3780 486892 3782
rect 486916 3780 486972 3782
rect 486996 3780 487052 3782
rect 487076 3780 487132 3782
rect 487156 3780 487212 3782
rect 487236 3780 487292 3782
rect 487316 3780 487372 3782
rect 486836 2746 486892 2748
rect 486916 2746 486972 2748
rect 486996 2746 487052 2748
rect 487076 2746 487132 2748
rect 487156 2746 487212 2748
rect 487236 2746 487292 2748
rect 487316 2746 487372 2748
rect 486836 2694 486874 2746
rect 486874 2694 486886 2746
rect 486886 2694 486892 2746
rect 486916 2694 486938 2746
rect 486938 2694 486950 2746
rect 486950 2694 486972 2746
rect 486996 2694 487002 2746
rect 487002 2694 487014 2746
rect 487014 2694 487052 2746
rect 487076 2694 487078 2746
rect 487078 2694 487130 2746
rect 487130 2694 487132 2746
rect 487156 2694 487194 2746
rect 487194 2694 487206 2746
rect 487206 2694 487212 2746
rect 487236 2694 487258 2746
rect 487258 2694 487270 2746
rect 487270 2694 487292 2746
rect 487316 2694 487322 2746
rect 487322 2694 487334 2746
rect 487334 2694 487372 2746
rect 486836 2692 486892 2694
rect 486916 2692 486972 2694
rect 486996 2692 487052 2694
rect 487076 2692 487132 2694
rect 487156 2692 487212 2694
rect 487236 2692 487292 2694
rect 487316 2692 487372 2694
rect 504836 5466 504892 5468
rect 504916 5466 504972 5468
rect 504996 5466 505052 5468
rect 505076 5466 505132 5468
rect 505156 5466 505212 5468
rect 505236 5466 505292 5468
rect 505316 5466 505372 5468
rect 504836 5414 504874 5466
rect 504874 5414 504886 5466
rect 504886 5414 504892 5466
rect 504916 5414 504938 5466
rect 504938 5414 504950 5466
rect 504950 5414 504972 5466
rect 504996 5414 505002 5466
rect 505002 5414 505014 5466
rect 505014 5414 505052 5466
rect 505076 5414 505078 5466
rect 505078 5414 505130 5466
rect 505130 5414 505132 5466
rect 505156 5414 505194 5466
rect 505194 5414 505206 5466
rect 505206 5414 505212 5466
rect 505236 5414 505258 5466
rect 505258 5414 505270 5466
rect 505270 5414 505292 5466
rect 505316 5414 505322 5466
rect 505322 5414 505334 5466
rect 505334 5414 505372 5466
rect 504836 5412 504892 5414
rect 504916 5412 504972 5414
rect 504996 5412 505052 5414
rect 505076 5412 505132 5414
rect 505156 5412 505212 5414
rect 505236 5412 505292 5414
rect 505316 5412 505372 5414
rect 504836 4378 504892 4380
rect 504916 4378 504972 4380
rect 504996 4378 505052 4380
rect 505076 4378 505132 4380
rect 505156 4378 505212 4380
rect 505236 4378 505292 4380
rect 505316 4378 505372 4380
rect 504836 4326 504874 4378
rect 504874 4326 504886 4378
rect 504886 4326 504892 4378
rect 504916 4326 504938 4378
rect 504938 4326 504950 4378
rect 504950 4326 504972 4378
rect 504996 4326 505002 4378
rect 505002 4326 505014 4378
rect 505014 4326 505052 4378
rect 505076 4326 505078 4378
rect 505078 4326 505130 4378
rect 505130 4326 505132 4378
rect 505156 4326 505194 4378
rect 505194 4326 505206 4378
rect 505206 4326 505212 4378
rect 505236 4326 505258 4378
rect 505258 4326 505270 4378
rect 505270 4326 505292 4378
rect 505316 4326 505322 4378
rect 505322 4326 505334 4378
rect 505334 4326 505372 4378
rect 504836 4324 504892 4326
rect 504916 4324 504972 4326
rect 504996 4324 505052 4326
rect 505076 4324 505132 4326
rect 505156 4324 505212 4326
rect 505236 4324 505292 4326
rect 505316 4324 505372 4326
rect 504836 3290 504892 3292
rect 504916 3290 504972 3292
rect 504996 3290 505052 3292
rect 505076 3290 505132 3292
rect 505156 3290 505212 3292
rect 505236 3290 505292 3292
rect 505316 3290 505372 3292
rect 504836 3238 504874 3290
rect 504874 3238 504886 3290
rect 504886 3238 504892 3290
rect 504916 3238 504938 3290
rect 504938 3238 504950 3290
rect 504950 3238 504972 3290
rect 504996 3238 505002 3290
rect 505002 3238 505014 3290
rect 505014 3238 505052 3290
rect 505076 3238 505078 3290
rect 505078 3238 505130 3290
rect 505130 3238 505132 3290
rect 505156 3238 505194 3290
rect 505194 3238 505206 3290
rect 505206 3238 505212 3290
rect 505236 3238 505258 3290
rect 505258 3238 505270 3290
rect 505270 3238 505292 3290
rect 505316 3238 505322 3290
rect 505322 3238 505334 3290
rect 505334 3238 505372 3290
rect 504836 3236 504892 3238
rect 504916 3236 504972 3238
rect 504996 3236 505052 3238
rect 505076 3236 505132 3238
rect 505156 3236 505212 3238
rect 505236 3236 505292 3238
rect 505316 3236 505372 3238
rect 504836 2202 504892 2204
rect 504916 2202 504972 2204
rect 504996 2202 505052 2204
rect 505076 2202 505132 2204
rect 505156 2202 505212 2204
rect 505236 2202 505292 2204
rect 505316 2202 505372 2204
rect 504836 2150 504874 2202
rect 504874 2150 504886 2202
rect 504886 2150 504892 2202
rect 504916 2150 504938 2202
rect 504938 2150 504950 2202
rect 504950 2150 504972 2202
rect 504996 2150 505002 2202
rect 505002 2150 505014 2202
rect 505014 2150 505052 2202
rect 505076 2150 505078 2202
rect 505078 2150 505130 2202
rect 505130 2150 505132 2202
rect 505156 2150 505194 2202
rect 505194 2150 505206 2202
rect 505206 2150 505212 2202
rect 505236 2150 505258 2202
rect 505258 2150 505270 2202
rect 505270 2150 505292 2202
rect 505316 2150 505322 2202
rect 505322 2150 505334 2202
rect 505334 2150 505372 2202
rect 504836 2148 504892 2150
rect 504916 2148 504972 2150
rect 504996 2148 505052 2150
rect 505076 2148 505132 2150
rect 505156 2148 505212 2150
rect 505236 2148 505292 2150
rect 505316 2148 505372 2150
rect 522836 6010 522892 6012
rect 522916 6010 522972 6012
rect 522996 6010 523052 6012
rect 523076 6010 523132 6012
rect 523156 6010 523212 6012
rect 523236 6010 523292 6012
rect 523316 6010 523372 6012
rect 522836 5958 522874 6010
rect 522874 5958 522886 6010
rect 522886 5958 522892 6010
rect 522916 5958 522938 6010
rect 522938 5958 522950 6010
rect 522950 5958 522972 6010
rect 522996 5958 523002 6010
rect 523002 5958 523014 6010
rect 523014 5958 523052 6010
rect 523076 5958 523078 6010
rect 523078 5958 523130 6010
rect 523130 5958 523132 6010
rect 523156 5958 523194 6010
rect 523194 5958 523206 6010
rect 523206 5958 523212 6010
rect 523236 5958 523258 6010
rect 523258 5958 523270 6010
rect 523270 5958 523292 6010
rect 523316 5958 523322 6010
rect 523322 5958 523334 6010
rect 523334 5958 523372 6010
rect 522836 5956 522892 5958
rect 522916 5956 522972 5958
rect 522996 5956 523052 5958
rect 523076 5956 523132 5958
rect 523156 5956 523212 5958
rect 523236 5956 523292 5958
rect 523316 5956 523372 5958
rect 522836 4922 522892 4924
rect 522916 4922 522972 4924
rect 522996 4922 523052 4924
rect 523076 4922 523132 4924
rect 523156 4922 523212 4924
rect 523236 4922 523292 4924
rect 523316 4922 523372 4924
rect 522836 4870 522874 4922
rect 522874 4870 522886 4922
rect 522886 4870 522892 4922
rect 522916 4870 522938 4922
rect 522938 4870 522950 4922
rect 522950 4870 522972 4922
rect 522996 4870 523002 4922
rect 523002 4870 523014 4922
rect 523014 4870 523052 4922
rect 523076 4870 523078 4922
rect 523078 4870 523130 4922
rect 523130 4870 523132 4922
rect 523156 4870 523194 4922
rect 523194 4870 523206 4922
rect 523206 4870 523212 4922
rect 523236 4870 523258 4922
rect 523258 4870 523270 4922
rect 523270 4870 523292 4922
rect 523316 4870 523322 4922
rect 523322 4870 523334 4922
rect 523334 4870 523372 4922
rect 522836 4868 522892 4870
rect 522916 4868 522972 4870
rect 522996 4868 523052 4870
rect 523076 4868 523132 4870
rect 523156 4868 523212 4870
rect 523236 4868 523292 4870
rect 523316 4868 523372 4870
rect 522836 3834 522892 3836
rect 522916 3834 522972 3836
rect 522996 3834 523052 3836
rect 523076 3834 523132 3836
rect 523156 3834 523212 3836
rect 523236 3834 523292 3836
rect 523316 3834 523372 3836
rect 522836 3782 522874 3834
rect 522874 3782 522886 3834
rect 522886 3782 522892 3834
rect 522916 3782 522938 3834
rect 522938 3782 522950 3834
rect 522950 3782 522972 3834
rect 522996 3782 523002 3834
rect 523002 3782 523014 3834
rect 523014 3782 523052 3834
rect 523076 3782 523078 3834
rect 523078 3782 523130 3834
rect 523130 3782 523132 3834
rect 523156 3782 523194 3834
rect 523194 3782 523206 3834
rect 523206 3782 523212 3834
rect 523236 3782 523258 3834
rect 523258 3782 523270 3834
rect 523270 3782 523292 3834
rect 523316 3782 523322 3834
rect 523322 3782 523334 3834
rect 523334 3782 523372 3834
rect 522836 3780 522892 3782
rect 522916 3780 522972 3782
rect 522996 3780 523052 3782
rect 523076 3780 523132 3782
rect 523156 3780 523212 3782
rect 523236 3780 523292 3782
rect 523316 3780 523372 3782
rect 522836 2746 522892 2748
rect 522916 2746 522972 2748
rect 522996 2746 523052 2748
rect 523076 2746 523132 2748
rect 523156 2746 523212 2748
rect 523236 2746 523292 2748
rect 523316 2746 523372 2748
rect 522836 2694 522874 2746
rect 522874 2694 522886 2746
rect 522886 2694 522892 2746
rect 522916 2694 522938 2746
rect 522938 2694 522950 2746
rect 522950 2694 522972 2746
rect 522996 2694 523002 2746
rect 523002 2694 523014 2746
rect 523014 2694 523052 2746
rect 523076 2694 523078 2746
rect 523078 2694 523130 2746
rect 523130 2694 523132 2746
rect 523156 2694 523194 2746
rect 523194 2694 523206 2746
rect 523206 2694 523212 2746
rect 523236 2694 523258 2746
rect 523258 2694 523270 2746
rect 523270 2694 523292 2746
rect 523316 2694 523322 2746
rect 523322 2694 523334 2746
rect 523334 2694 523372 2746
rect 522836 2692 522892 2694
rect 522916 2692 522972 2694
rect 522996 2692 523052 2694
rect 523076 2692 523132 2694
rect 523156 2692 523212 2694
rect 523236 2692 523292 2694
rect 523316 2692 523372 2694
rect 540836 5466 540892 5468
rect 540916 5466 540972 5468
rect 540996 5466 541052 5468
rect 541076 5466 541132 5468
rect 541156 5466 541212 5468
rect 541236 5466 541292 5468
rect 541316 5466 541372 5468
rect 540836 5414 540874 5466
rect 540874 5414 540886 5466
rect 540886 5414 540892 5466
rect 540916 5414 540938 5466
rect 540938 5414 540950 5466
rect 540950 5414 540972 5466
rect 540996 5414 541002 5466
rect 541002 5414 541014 5466
rect 541014 5414 541052 5466
rect 541076 5414 541078 5466
rect 541078 5414 541130 5466
rect 541130 5414 541132 5466
rect 541156 5414 541194 5466
rect 541194 5414 541206 5466
rect 541206 5414 541212 5466
rect 541236 5414 541258 5466
rect 541258 5414 541270 5466
rect 541270 5414 541292 5466
rect 541316 5414 541322 5466
rect 541322 5414 541334 5466
rect 541334 5414 541372 5466
rect 540836 5412 540892 5414
rect 540916 5412 540972 5414
rect 540996 5412 541052 5414
rect 541076 5412 541132 5414
rect 541156 5412 541212 5414
rect 541236 5412 541292 5414
rect 541316 5412 541372 5414
rect 540836 4378 540892 4380
rect 540916 4378 540972 4380
rect 540996 4378 541052 4380
rect 541076 4378 541132 4380
rect 541156 4378 541212 4380
rect 541236 4378 541292 4380
rect 541316 4378 541372 4380
rect 540836 4326 540874 4378
rect 540874 4326 540886 4378
rect 540886 4326 540892 4378
rect 540916 4326 540938 4378
rect 540938 4326 540950 4378
rect 540950 4326 540972 4378
rect 540996 4326 541002 4378
rect 541002 4326 541014 4378
rect 541014 4326 541052 4378
rect 541076 4326 541078 4378
rect 541078 4326 541130 4378
rect 541130 4326 541132 4378
rect 541156 4326 541194 4378
rect 541194 4326 541206 4378
rect 541206 4326 541212 4378
rect 541236 4326 541258 4378
rect 541258 4326 541270 4378
rect 541270 4326 541292 4378
rect 541316 4326 541322 4378
rect 541322 4326 541334 4378
rect 541334 4326 541372 4378
rect 540836 4324 540892 4326
rect 540916 4324 540972 4326
rect 540996 4324 541052 4326
rect 541076 4324 541132 4326
rect 541156 4324 541212 4326
rect 541236 4324 541292 4326
rect 541316 4324 541372 4326
rect 540836 3290 540892 3292
rect 540916 3290 540972 3292
rect 540996 3290 541052 3292
rect 541076 3290 541132 3292
rect 541156 3290 541212 3292
rect 541236 3290 541292 3292
rect 541316 3290 541372 3292
rect 540836 3238 540874 3290
rect 540874 3238 540886 3290
rect 540886 3238 540892 3290
rect 540916 3238 540938 3290
rect 540938 3238 540950 3290
rect 540950 3238 540972 3290
rect 540996 3238 541002 3290
rect 541002 3238 541014 3290
rect 541014 3238 541052 3290
rect 541076 3238 541078 3290
rect 541078 3238 541130 3290
rect 541130 3238 541132 3290
rect 541156 3238 541194 3290
rect 541194 3238 541206 3290
rect 541206 3238 541212 3290
rect 541236 3238 541258 3290
rect 541258 3238 541270 3290
rect 541270 3238 541292 3290
rect 541316 3238 541322 3290
rect 541322 3238 541334 3290
rect 541334 3238 541372 3290
rect 540836 3236 540892 3238
rect 540916 3236 540972 3238
rect 540996 3236 541052 3238
rect 541076 3236 541132 3238
rect 541156 3236 541212 3238
rect 541236 3236 541292 3238
rect 541316 3236 541372 3238
rect 540836 2202 540892 2204
rect 540916 2202 540972 2204
rect 540996 2202 541052 2204
rect 541076 2202 541132 2204
rect 541156 2202 541212 2204
rect 541236 2202 541292 2204
rect 541316 2202 541372 2204
rect 540836 2150 540874 2202
rect 540874 2150 540886 2202
rect 540886 2150 540892 2202
rect 540916 2150 540938 2202
rect 540938 2150 540950 2202
rect 540950 2150 540972 2202
rect 540996 2150 541002 2202
rect 541002 2150 541014 2202
rect 541014 2150 541052 2202
rect 541076 2150 541078 2202
rect 541078 2150 541130 2202
rect 541130 2150 541132 2202
rect 541156 2150 541194 2202
rect 541194 2150 541206 2202
rect 541206 2150 541212 2202
rect 541236 2150 541258 2202
rect 541258 2150 541270 2202
rect 541270 2150 541292 2202
rect 541316 2150 541322 2202
rect 541322 2150 541334 2202
rect 541334 2150 541372 2202
rect 540836 2148 540892 2150
rect 540916 2148 540972 2150
rect 540996 2148 541052 2150
rect 541076 2148 541132 2150
rect 541156 2148 541212 2150
rect 541236 2148 541292 2150
rect 541316 2148 541372 2150
rect 558836 6010 558892 6012
rect 558916 6010 558972 6012
rect 558996 6010 559052 6012
rect 559076 6010 559132 6012
rect 559156 6010 559212 6012
rect 559236 6010 559292 6012
rect 559316 6010 559372 6012
rect 558836 5958 558874 6010
rect 558874 5958 558886 6010
rect 558886 5958 558892 6010
rect 558916 5958 558938 6010
rect 558938 5958 558950 6010
rect 558950 5958 558972 6010
rect 558996 5958 559002 6010
rect 559002 5958 559014 6010
rect 559014 5958 559052 6010
rect 559076 5958 559078 6010
rect 559078 5958 559130 6010
rect 559130 5958 559132 6010
rect 559156 5958 559194 6010
rect 559194 5958 559206 6010
rect 559206 5958 559212 6010
rect 559236 5958 559258 6010
rect 559258 5958 559270 6010
rect 559270 5958 559292 6010
rect 559316 5958 559322 6010
rect 559322 5958 559334 6010
rect 559334 5958 559372 6010
rect 558836 5956 558892 5958
rect 558916 5956 558972 5958
rect 558996 5956 559052 5958
rect 559076 5956 559132 5958
rect 559156 5956 559212 5958
rect 559236 5956 559292 5958
rect 559316 5956 559372 5958
rect 558836 4922 558892 4924
rect 558916 4922 558972 4924
rect 558996 4922 559052 4924
rect 559076 4922 559132 4924
rect 559156 4922 559212 4924
rect 559236 4922 559292 4924
rect 559316 4922 559372 4924
rect 558836 4870 558874 4922
rect 558874 4870 558886 4922
rect 558886 4870 558892 4922
rect 558916 4870 558938 4922
rect 558938 4870 558950 4922
rect 558950 4870 558972 4922
rect 558996 4870 559002 4922
rect 559002 4870 559014 4922
rect 559014 4870 559052 4922
rect 559076 4870 559078 4922
rect 559078 4870 559130 4922
rect 559130 4870 559132 4922
rect 559156 4870 559194 4922
rect 559194 4870 559206 4922
rect 559206 4870 559212 4922
rect 559236 4870 559258 4922
rect 559258 4870 559270 4922
rect 559270 4870 559292 4922
rect 559316 4870 559322 4922
rect 559322 4870 559334 4922
rect 559334 4870 559372 4922
rect 558836 4868 558892 4870
rect 558916 4868 558972 4870
rect 558996 4868 559052 4870
rect 559076 4868 559132 4870
rect 559156 4868 559212 4870
rect 559236 4868 559292 4870
rect 559316 4868 559372 4870
rect 558836 3834 558892 3836
rect 558916 3834 558972 3836
rect 558996 3834 559052 3836
rect 559076 3834 559132 3836
rect 559156 3834 559212 3836
rect 559236 3834 559292 3836
rect 559316 3834 559372 3836
rect 558836 3782 558874 3834
rect 558874 3782 558886 3834
rect 558886 3782 558892 3834
rect 558916 3782 558938 3834
rect 558938 3782 558950 3834
rect 558950 3782 558972 3834
rect 558996 3782 559002 3834
rect 559002 3782 559014 3834
rect 559014 3782 559052 3834
rect 559076 3782 559078 3834
rect 559078 3782 559130 3834
rect 559130 3782 559132 3834
rect 559156 3782 559194 3834
rect 559194 3782 559206 3834
rect 559206 3782 559212 3834
rect 559236 3782 559258 3834
rect 559258 3782 559270 3834
rect 559270 3782 559292 3834
rect 559316 3782 559322 3834
rect 559322 3782 559334 3834
rect 559334 3782 559372 3834
rect 558836 3780 558892 3782
rect 558916 3780 558972 3782
rect 558996 3780 559052 3782
rect 559076 3780 559132 3782
rect 559156 3780 559212 3782
rect 559236 3780 559292 3782
rect 559316 3780 559372 3782
rect 558836 2746 558892 2748
rect 558916 2746 558972 2748
rect 558996 2746 559052 2748
rect 559076 2746 559132 2748
rect 559156 2746 559212 2748
rect 559236 2746 559292 2748
rect 559316 2746 559372 2748
rect 558836 2694 558874 2746
rect 558874 2694 558886 2746
rect 558886 2694 558892 2746
rect 558916 2694 558938 2746
rect 558938 2694 558950 2746
rect 558950 2694 558972 2746
rect 558996 2694 559002 2746
rect 559002 2694 559014 2746
rect 559014 2694 559052 2746
rect 559076 2694 559078 2746
rect 559078 2694 559130 2746
rect 559130 2694 559132 2746
rect 559156 2694 559194 2746
rect 559194 2694 559206 2746
rect 559206 2694 559212 2746
rect 559236 2694 559258 2746
rect 559258 2694 559270 2746
rect 559270 2694 559292 2746
rect 559316 2694 559322 2746
rect 559322 2694 559334 2746
rect 559334 2694 559372 2746
rect 558836 2692 558892 2694
rect 558916 2692 558972 2694
rect 558996 2692 559052 2694
rect 559076 2692 559132 2694
rect 559156 2692 559212 2694
rect 559236 2692 559292 2694
rect 559316 2692 559372 2694
rect 576836 5466 576892 5468
rect 576916 5466 576972 5468
rect 576996 5466 577052 5468
rect 577076 5466 577132 5468
rect 577156 5466 577212 5468
rect 577236 5466 577292 5468
rect 577316 5466 577372 5468
rect 576836 5414 576874 5466
rect 576874 5414 576886 5466
rect 576886 5414 576892 5466
rect 576916 5414 576938 5466
rect 576938 5414 576950 5466
rect 576950 5414 576972 5466
rect 576996 5414 577002 5466
rect 577002 5414 577014 5466
rect 577014 5414 577052 5466
rect 577076 5414 577078 5466
rect 577078 5414 577130 5466
rect 577130 5414 577132 5466
rect 577156 5414 577194 5466
rect 577194 5414 577206 5466
rect 577206 5414 577212 5466
rect 577236 5414 577258 5466
rect 577258 5414 577270 5466
rect 577270 5414 577292 5466
rect 577316 5414 577322 5466
rect 577322 5414 577334 5466
rect 577334 5414 577372 5466
rect 576836 5412 576892 5414
rect 576916 5412 576972 5414
rect 576996 5412 577052 5414
rect 577076 5412 577132 5414
rect 577156 5412 577212 5414
rect 577236 5412 577292 5414
rect 577316 5412 577372 5414
rect 576836 4378 576892 4380
rect 576916 4378 576972 4380
rect 576996 4378 577052 4380
rect 577076 4378 577132 4380
rect 577156 4378 577212 4380
rect 577236 4378 577292 4380
rect 577316 4378 577372 4380
rect 576836 4326 576874 4378
rect 576874 4326 576886 4378
rect 576886 4326 576892 4378
rect 576916 4326 576938 4378
rect 576938 4326 576950 4378
rect 576950 4326 576972 4378
rect 576996 4326 577002 4378
rect 577002 4326 577014 4378
rect 577014 4326 577052 4378
rect 577076 4326 577078 4378
rect 577078 4326 577130 4378
rect 577130 4326 577132 4378
rect 577156 4326 577194 4378
rect 577194 4326 577206 4378
rect 577206 4326 577212 4378
rect 577236 4326 577258 4378
rect 577258 4326 577270 4378
rect 577270 4326 577292 4378
rect 577316 4326 577322 4378
rect 577322 4326 577334 4378
rect 577334 4326 577372 4378
rect 576836 4324 576892 4326
rect 576916 4324 576972 4326
rect 576996 4324 577052 4326
rect 577076 4324 577132 4326
rect 577156 4324 577212 4326
rect 577236 4324 577292 4326
rect 577316 4324 577372 4326
rect 576836 3290 576892 3292
rect 576916 3290 576972 3292
rect 576996 3290 577052 3292
rect 577076 3290 577132 3292
rect 577156 3290 577212 3292
rect 577236 3290 577292 3292
rect 577316 3290 577372 3292
rect 576836 3238 576874 3290
rect 576874 3238 576886 3290
rect 576886 3238 576892 3290
rect 576916 3238 576938 3290
rect 576938 3238 576950 3290
rect 576950 3238 576972 3290
rect 576996 3238 577002 3290
rect 577002 3238 577014 3290
rect 577014 3238 577052 3290
rect 577076 3238 577078 3290
rect 577078 3238 577130 3290
rect 577130 3238 577132 3290
rect 577156 3238 577194 3290
rect 577194 3238 577206 3290
rect 577206 3238 577212 3290
rect 577236 3238 577258 3290
rect 577258 3238 577270 3290
rect 577270 3238 577292 3290
rect 577316 3238 577322 3290
rect 577322 3238 577334 3290
rect 577334 3238 577372 3290
rect 576836 3236 576892 3238
rect 576916 3236 576972 3238
rect 576996 3236 577052 3238
rect 577076 3236 577132 3238
rect 577156 3236 577212 3238
rect 577236 3236 577292 3238
rect 577316 3236 577372 3238
rect 576836 2202 576892 2204
rect 576916 2202 576972 2204
rect 576996 2202 577052 2204
rect 577076 2202 577132 2204
rect 577156 2202 577212 2204
rect 577236 2202 577292 2204
rect 577316 2202 577372 2204
rect 576836 2150 576874 2202
rect 576874 2150 576886 2202
rect 576886 2150 576892 2202
rect 576916 2150 576938 2202
rect 576938 2150 576950 2202
rect 576950 2150 576972 2202
rect 576996 2150 577002 2202
rect 577002 2150 577014 2202
rect 577014 2150 577052 2202
rect 577076 2150 577078 2202
rect 577078 2150 577130 2202
rect 577130 2150 577132 2202
rect 577156 2150 577194 2202
rect 577194 2150 577206 2202
rect 577206 2150 577212 2202
rect 577236 2150 577258 2202
rect 577258 2150 577270 2202
rect 577270 2150 577292 2202
rect 577316 2150 577322 2202
rect 577322 2150 577334 2202
rect 577334 2150 577372 2202
rect 576836 2148 576892 2150
rect 576916 2148 576972 2150
rect 576996 2148 577052 2150
rect 577076 2148 577132 2150
rect 577156 2148 577212 2150
rect 577236 2148 577292 2150
rect 577316 2148 577372 2150
<< metal3 >>
rect 36804 701792 37404 701793
rect 36804 701728 36832 701792
rect 36896 701728 36912 701792
rect 36976 701728 36992 701792
rect 37056 701728 37072 701792
rect 37136 701728 37152 701792
rect 37216 701728 37232 701792
rect 37296 701728 37312 701792
rect 37376 701728 37404 701792
rect 36804 701727 37404 701728
rect 72804 701792 73404 701793
rect 72804 701728 72832 701792
rect 72896 701728 72912 701792
rect 72976 701728 72992 701792
rect 73056 701728 73072 701792
rect 73136 701728 73152 701792
rect 73216 701728 73232 701792
rect 73296 701728 73312 701792
rect 73376 701728 73404 701792
rect 72804 701727 73404 701728
rect 108804 701792 109404 701793
rect 108804 701728 108832 701792
rect 108896 701728 108912 701792
rect 108976 701728 108992 701792
rect 109056 701728 109072 701792
rect 109136 701728 109152 701792
rect 109216 701728 109232 701792
rect 109296 701728 109312 701792
rect 109376 701728 109404 701792
rect 108804 701727 109404 701728
rect 144804 701792 145404 701793
rect 144804 701728 144832 701792
rect 144896 701728 144912 701792
rect 144976 701728 144992 701792
rect 145056 701728 145072 701792
rect 145136 701728 145152 701792
rect 145216 701728 145232 701792
rect 145296 701728 145312 701792
rect 145376 701728 145404 701792
rect 144804 701727 145404 701728
rect 180804 701792 181404 701793
rect 180804 701728 180832 701792
rect 180896 701728 180912 701792
rect 180976 701728 180992 701792
rect 181056 701728 181072 701792
rect 181136 701728 181152 701792
rect 181216 701728 181232 701792
rect 181296 701728 181312 701792
rect 181376 701728 181404 701792
rect 180804 701727 181404 701728
rect 216804 701792 217404 701793
rect 216804 701728 216832 701792
rect 216896 701728 216912 701792
rect 216976 701728 216992 701792
rect 217056 701728 217072 701792
rect 217136 701728 217152 701792
rect 217216 701728 217232 701792
rect 217296 701728 217312 701792
rect 217376 701728 217404 701792
rect 216804 701727 217404 701728
rect 252804 701792 253404 701793
rect 252804 701728 252832 701792
rect 252896 701728 252912 701792
rect 252976 701728 252992 701792
rect 253056 701728 253072 701792
rect 253136 701728 253152 701792
rect 253216 701728 253232 701792
rect 253296 701728 253312 701792
rect 253376 701728 253404 701792
rect 252804 701727 253404 701728
rect 288804 701792 289404 701793
rect 288804 701728 288832 701792
rect 288896 701728 288912 701792
rect 288976 701728 288992 701792
rect 289056 701728 289072 701792
rect 289136 701728 289152 701792
rect 289216 701728 289232 701792
rect 289296 701728 289312 701792
rect 289376 701728 289404 701792
rect 288804 701727 289404 701728
rect 324804 701792 325404 701793
rect 324804 701728 324832 701792
rect 324896 701728 324912 701792
rect 324976 701728 324992 701792
rect 325056 701728 325072 701792
rect 325136 701728 325152 701792
rect 325216 701728 325232 701792
rect 325296 701728 325312 701792
rect 325376 701728 325404 701792
rect 324804 701727 325404 701728
rect 360804 701792 361404 701793
rect 360804 701728 360832 701792
rect 360896 701728 360912 701792
rect 360976 701728 360992 701792
rect 361056 701728 361072 701792
rect 361136 701728 361152 701792
rect 361216 701728 361232 701792
rect 361296 701728 361312 701792
rect 361376 701728 361404 701792
rect 360804 701727 361404 701728
rect 396804 701792 397404 701793
rect 396804 701728 396832 701792
rect 396896 701728 396912 701792
rect 396976 701728 396992 701792
rect 397056 701728 397072 701792
rect 397136 701728 397152 701792
rect 397216 701728 397232 701792
rect 397296 701728 397312 701792
rect 397376 701728 397404 701792
rect 396804 701727 397404 701728
rect 432804 701792 433404 701793
rect 432804 701728 432832 701792
rect 432896 701728 432912 701792
rect 432976 701728 432992 701792
rect 433056 701728 433072 701792
rect 433136 701728 433152 701792
rect 433216 701728 433232 701792
rect 433296 701728 433312 701792
rect 433376 701728 433404 701792
rect 432804 701727 433404 701728
rect 468804 701792 469404 701793
rect 468804 701728 468832 701792
rect 468896 701728 468912 701792
rect 468976 701728 468992 701792
rect 469056 701728 469072 701792
rect 469136 701728 469152 701792
rect 469216 701728 469232 701792
rect 469296 701728 469312 701792
rect 469376 701728 469404 701792
rect 468804 701727 469404 701728
rect 504804 701792 505404 701793
rect 504804 701728 504832 701792
rect 504896 701728 504912 701792
rect 504976 701728 504992 701792
rect 505056 701728 505072 701792
rect 505136 701728 505152 701792
rect 505216 701728 505232 701792
rect 505296 701728 505312 701792
rect 505376 701728 505404 701792
rect 504804 701727 505404 701728
rect 540804 701792 541404 701793
rect 540804 701728 540832 701792
rect 540896 701728 540912 701792
rect 540976 701728 540992 701792
rect 541056 701728 541072 701792
rect 541136 701728 541152 701792
rect 541216 701728 541232 701792
rect 541296 701728 541312 701792
rect 541376 701728 541404 701792
rect 540804 701727 541404 701728
rect 576804 701792 577404 701793
rect 576804 701728 576832 701792
rect 576896 701728 576912 701792
rect 576976 701728 576992 701792
rect 577056 701728 577072 701792
rect 577136 701728 577152 701792
rect 577216 701728 577232 701792
rect 577296 701728 577312 701792
rect 577376 701728 577404 701792
rect 576804 701727 577404 701728
rect 18804 701248 19404 701249
rect 18804 701184 18832 701248
rect 18896 701184 18912 701248
rect 18976 701184 18992 701248
rect 19056 701184 19072 701248
rect 19136 701184 19152 701248
rect 19216 701184 19232 701248
rect 19296 701184 19312 701248
rect 19376 701184 19404 701248
rect 18804 701183 19404 701184
rect 54804 701248 55404 701249
rect 54804 701184 54832 701248
rect 54896 701184 54912 701248
rect 54976 701184 54992 701248
rect 55056 701184 55072 701248
rect 55136 701184 55152 701248
rect 55216 701184 55232 701248
rect 55296 701184 55312 701248
rect 55376 701184 55404 701248
rect 54804 701183 55404 701184
rect 90804 701248 91404 701249
rect 90804 701184 90832 701248
rect 90896 701184 90912 701248
rect 90976 701184 90992 701248
rect 91056 701184 91072 701248
rect 91136 701184 91152 701248
rect 91216 701184 91232 701248
rect 91296 701184 91312 701248
rect 91376 701184 91404 701248
rect 90804 701183 91404 701184
rect 126804 701248 127404 701249
rect 126804 701184 126832 701248
rect 126896 701184 126912 701248
rect 126976 701184 126992 701248
rect 127056 701184 127072 701248
rect 127136 701184 127152 701248
rect 127216 701184 127232 701248
rect 127296 701184 127312 701248
rect 127376 701184 127404 701248
rect 126804 701183 127404 701184
rect 162804 701248 163404 701249
rect 162804 701184 162832 701248
rect 162896 701184 162912 701248
rect 162976 701184 162992 701248
rect 163056 701184 163072 701248
rect 163136 701184 163152 701248
rect 163216 701184 163232 701248
rect 163296 701184 163312 701248
rect 163376 701184 163404 701248
rect 162804 701183 163404 701184
rect 198804 701248 199404 701249
rect 198804 701184 198832 701248
rect 198896 701184 198912 701248
rect 198976 701184 198992 701248
rect 199056 701184 199072 701248
rect 199136 701184 199152 701248
rect 199216 701184 199232 701248
rect 199296 701184 199312 701248
rect 199376 701184 199404 701248
rect 198804 701183 199404 701184
rect 234804 701248 235404 701249
rect 234804 701184 234832 701248
rect 234896 701184 234912 701248
rect 234976 701184 234992 701248
rect 235056 701184 235072 701248
rect 235136 701184 235152 701248
rect 235216 701184 235232 701248
rect 235296 701184 235312 701248
rect 235376 701184 235404 701248
rect 234804 701183 235404 701184
rect 270804 701248 271404 701249
rect 270804 701184 270832 701248
rect 270896 701184 270912 701248
rect 270976 701184 270992 701248
rect 271056 701184 271072 701248
rect 271136 701184 271152 701248
rect 271216 701184 271232 701248
rect 271296 701184 271312 701248
rect 271376 701184 271404 701248
rect 270804 701183 271404 701184
rect 306804 701248 307404 701249
rect 306804 701184 306832 701248
rect 306896 701184 306912 701248
rect 306976 701184 306992 701248
rect 307056 701184 307072 701248
rect 307136 701184 307152 701248
rect 307216 701184 307232 701248
rect 307296 701184 307312 701248
rect 307376 701184 307404 701248
rect 306804 701183 307404 701184
rect 342804 701248 343404 701249
rect 342804 701184 342832 701248
rect 342896 701184 342912 701248
rect 342976 701184 342992 701248
rect 343056 701184 343072 701248
rect 343136 701184 343152 701248
rect 343216 701184 343232 701248
rect 343296 701184 343312 701248
rect 343376 701184 343404 701248
rect 342804 701183 343404 701184
rect 378804 701248 379404 701249
rect 378804 701184 378832 701248
rect 378896 701184 378912 701248
rect 378976 701184 378992 701248
rect 379056 701184 379072 701248
rect 379136 701184 379152 701248
rect 379216 701184 379232 701248
rect 379296 701184 379312 701248
rect 379376 701184 379404 701248
rect 378804 701183 379404 701184
rect 414804 701248 415404 701249
rect 414804 701184 414832 701248
rect 414896 701184 414912 701248
rect 414976 701184 414992 701248
rect 415056 701184 415072 701248
rect 415136 701184 415152 701248
rect 415216 701184 415232 701248
rect 415296 701184 415312 701248
rect 415376 701184 415404 701248
rect 414804 701183 415404 701184
rect 450804 701248 451404 701249
rect 450804 701184 450832 701248
rect 450896 701184 450912 701248
rect 450976 701184 450992 701248
rect 451056 701184 451072 701248
rect 451136 701184 451152 701248
rect 451216 701184 451232 701248
rect 451296 701184 451312 701248
rect 451376 701184 451404 701248
rect 450804 701183 451404 701184
rect 486804 701248 487404 701249
rect 486804 701184 486832 701248
rect 486896 701184 486912 701248
rect 486976 701184 486992 701248
rect 487056 701184 487072 701248
rect 487136 701184 487152 701248
rect 487216 701184 487232 701248
rect 487296 701184 487312 701248
rect 487376 701184 487404 701248
rect 486804 701183 487404 701184
rect 522804 701248 523404 701249
rect 522804 701184 522832 701248
rect 522896 701184 522912 701248
rect 522976 701184 522992 701248
rect 523056 701184 523072 701248
rect 523136 701184 523152 701248
rect 523216 701184 523232 701248
rect 523296 701184 523312 701248
rect 523376 701184 523404 701248
rect 522804 701183 523404 701184
rect 558804 701248 559404 701249
rect 558804 701184 558832 701248
rect 558896 701184 558912 701248
rect 558976 701184 558992 701248
rect 559056 701184 559072 701248
rect 559136 701184 559152 701248
rect 559216 701184 559232 701248
rect 559296 701184 559312 701248
rect 559376 701184 559404 701248
rect 558804 701183 559404 701184
rect 40493 701042 40559 701045
rect 336917 701042 336983 701045
rect 40493 701040 336983 701042
rect 40493 700984 40498 701040
rect 40554 700984 336922 701040
rect 336978 700984 336983 701040
rect 40493 700982 336983 700984
rect 40493 700979 40559 700982
rect 336917 700979 336983 700982
rect 227989 700906 228055 700909
rect 527173 700906 527239 700909
rect 227989 700904 527239 700906
rect 227989 700848 227994 700904
rect 228050 700848 527178 700904
rect 527234 700848 527239 700904
rect 227989 700846 527239 700848
rect 227989 700843 228055 700846
rect 527173 700843 527239 700846
rect 36804 700704 37404 700705
rect 36804 700640 36832 700704
rect 36896 700640 36912 700704
rect 36976 700640 36992 700704
rect 37056 700640 37072 700704
rect 37136 700640 37152 700704
rect 37216 700640 37232 700704
rect 37296 700640 37312 700704
rect 37376 700640 37404 700704
rect 36804 700639 37404 700640
rect 72804 700704 73404 700705
rect 72804 700640 72832 700704
rect 72896 700640 72912 700704
rect 72976 700640 72992 700704
rect 73056 700640 73072 700704
rect 73136 700640 73152 700704
rect 73216 700640 73232 700704
rect 73296 700640 73312 700704
rect 73376 700640 73404 700704
rect 72804 700639 73404 700640
rect 108804 700704 109404 700705
rect 108804 700640 108832 700704
rect 108896 700640 108912 700704
rect 108976 700640 108992 700704
rect 109056 700640 109072 700704
rect 109136 700640 109152 700704
rect 109216 700640 109232 700704
rect 109296 700640 109312 700704
rect 109376 700640 109404 700704
rect 108804 700639 109404 700640
rect 144804 700704 145404 700705
rect 144804 700640 144832 700704
rect 144896 700640 144912 700704
rect 144976 700640 144992 700704
rect 145056 700640 145072 700704
rect 145136 700640 145152 700704
rect 145216 700640 145232 700704
rect 145296 700640 145312 700704
rect 145376 700640 145404 700704
rect 144804 700639 145404 700640
rect 180804 700704 181404 700705
rect 180804 700640 180832 700704
rect 180896 700640 180912 700704
rect 180976 700640 180992 700704
rect 181056 700640 181072 700704
rect 181136 700640 181152 700704
rect 181216 700640 181232 700704
rect 181296 700640 181312 700704
rect 181376 700640 181404 700704
rect 180804 700639 181404 700640
rect 216804 700704 217404 700705
rect 216804 700640 216832 700704
rect 216896 700640 216912 700704
rect 216976 700640 216992 700704
rect 217056 700640 217072 700704
rect 217136 700640 217152 700704
rect 217216 700640 217232 700704
rect 217296 700640 217312 700704
rect 217376 700640 217404 700704
rect 216804 700639 217404 700640
rect 252804 700704 253404 700705
rect 252804 700640 252832 700704
rect 252896 700640 252912 700704
rect 252976 700640 252992 700704
rect 253056 700640 253072 700704
rect 253136 700640 253152 700704
rect 253216 700640 253232 700704
rect 253296 700640 253312 700704
rect 253376 700640 253404 700704
rect 252804 700639 253404 700640
rect 288804 700704 289404 700705
rect 288804 700640 288832 700704
rect 288896 700640 288912 700704
rect 288976 700640 288992 700704
rect 289056 700640 289072 700704
rect 289136 700640 289152 700704
rect 289216 700640 289232 700704
rect 289296 700640 289312 700704
rect 289376 700640 289404 700704
rect 288804 700639 289404 700640
rect 324804 700704 325404 700705
rect 324804 700640 324832 700704
rect 324896 700640 324912 700704
rect 324976 700640 324992 700704
rect 325056 700640 325072 700704
rect 325136 700640 325152 700704
rect 325216 700640 325232 700704
rect 325296 700640 325312 700704
rect 325376 700640 325404 700704
rect 324804 700639 325404 700640
rect 360804 700704 361404 700705
rect 360804 700640 360832 700704
rect 360896 700640 360912 700704
rect 360976 700640 360992 700704
rect 361056 700640 361072 700704
rect 361136 700640 361152 700704
rect 361216 700640 361232 700704
rect 361296 700640 361312 700704
rect 361376 700640 361404 700704
rect 360804 700639 361404 700640
rect 396804 700704 397404 700705
rect 396804 700640 396832 700704
rect 396896 700640 396912 700704
rect 396976 700640 396992 700704
rect 397056 700640 397072 700704
rect 397136 700640 397152 700704
rect 397216 700640 397232 700704
rect 397296 700640 397312 700704
rect 397376 700640 397404 700704
rect 396804 700639 397404 700640
rect 432804 700704 433404 700705
rect 432804 700640 432832 700704
rect 432896 700640 432912 700704
rect 432976 700640 432992 700704
rect 433056 700640 433072 700704
rect 433136 700640 433152 700704
rect 433216 700640 433232 700704
rect 433296 700640 433312 700704
rect 433376 700640 433404 700704
rect 432804 700639 433404 700640
rect 468804 700704 469404 700705
rect 468804 700640 468832 700704
rect 468896 700640 468912 700704
rect 468976 700640 468992 700704
rect 469056 700640 469072 700704
rect 469136 700640 469152 700704
rect 469216 700640 469232 700704
rect 469296 700640 469312 700704
rect 469376 700640 469404 700704
rect 468804 700639 469404 700640
rect 504804 700704 505404 700705
rect 504804 700640 504832 700704
rect 504896 700640 504912 700704
rect 504976 700640 504992 700704
rect 505056 700640 505072 700704
rect 505136 700640 505152 700704
rect 505216 700640 505232 700704
rect 505296 700640 505312 700704
rect 505376 700640 505404 700704
rect 504804 700639 505404 700640
rect 540804 700704 541404 700705
rect 540804 700640 540832 700704
rect 540896 700640 540912 700704
rect 540976 700640 540992 700704
rect 541056 700640 541072 700704
rect 541136 700640 541152 700704
rect 541216 700640 541232 700704
rect 541296 700640 541312 700704
rect 541376 700640 541404 700704
rect 540804 700639 541404 700640
rect 576804 700704 577404 700705
rect 576804 700640 576832 700704
rect 576896 700640 576912 700704
rect 576976 700640 576992 700704
rect 577056 700640 577072 700704
rect 577136 700640 577152 700704
rect 577216 700640 577232 700704
rect 577296 700640 577312 700704
rect 577376 700640 577404 700704
rect 576804 700639 577404 700640
rect 24301 700498 24367 700501
rect 346301 700498 346367 700501
rect 24301 700496 346367 700498
rect 24301 700440 24306 700496
rect 24362 700440 346306 700496
rect 346362 700440 346367 700496
rect 24301 700438 346367 700440
rect 24301 700435 24367 700438
rect 346301 700435 346367 700438
rect 8109 700362 8175 700365
rect 341609 700362 341675 700365
rect 8109 700360 341675 700362
rect 8109 700304 8114 700360
rect 8170 700304 341614 700360
rect 341670 700304 341675 700360
rect 8109 700302 341675 700304
rect 8109 700299 8175 700302
rect 341609 700299 341675 700302
rect 292573 700226 292639 700229
rect 298645 700226 298711 700229
rect 292573 700224 298711 700226
rect 292573 700168 292578 700224
rect 292634 700168 298650 700224
rect 298706 700168 298711 700224
rect 292573 700166 298711 700168
rect 292573 700163 292639 700166
rect 298645 700163 298711 700166
rect 18804 700160 19404 700161
rect 18804 700096 18832 700160
rect 18896 700096 18912 700160
rect 18976 700096 18992 700160
rect 19056 700096 19072 700160
rect 19136 700096 19152 700160
rect 19216 700096 19232 700160
rect 19296 700096 19312 700160
rect 19376 700096 19404 700160
rect 18804 700095 19404 700096
rect 54804 700160 55404 700161
rect 54804 700096 54832 700160
rect 54896 700096 54912 700160
rect 54976 700096 54992 700160
rect 55056 700096 55072 700160
rect 55136 700096 55152 700160
rect 55216 700096 55232 700160
rect 55296 700096 55312 700160
rect 55376 700096 55404 700160
rect 54804 700095 55404 700096
rect 90804 700160 91404 700161
rect 90804 700096 90832 700160
rect 90896 700096 90912 700160
rect 90976 700096 90992 700160
rect 91056 700096 91072 700160
rect 91136 700096 91152 700160
rect 91216 700096 91232 700160
rect 91296 700096 91312 700160
rect 91376 700096 91404 700160
rect 90804 700095 91404 700096
rect 126804 700160 127404 700161
rect 126804 700096 126832 700160
rect 126896 700096 126912 700160
rect 126976 700096 126992 700160
rect 127056 700096 127072 700160
rect 127136 700096 127152 700160
rect 127216 700096 127232 700160
rect 127296 700096 127312 700160
rect 127376 700096 127404 700160
rect 126804 700095 127404 700096
rect 162804 700160 163404 700161
rect 162804 700096 162832 700160
rect 162896 700096 162912 700160
rect 162976 700096 162992 700160
rect 163056 700096 163072 700160
rect 163136 700096 163152 700160
rect 163216 700096 163232 700160
rect 163296 700096 163312 700160
rect 163376 700096 163404 700160
rect 162804 700095 163404 700096
rect 198804 700160 199404 700161
rect 198804 700096 198832 700160
rect 198896 700096 198912 700160
rect 198976 700096 198992 700160
rect 199056 700096 199072 700160
rect 199136 700096 199152 700160
rect 199216 700096 199232 700160
rect 199296 700096 199312 700160
rect 199376 700096 199404 700160
rect 198804 700095 199404 700096
rect 234804 700160 235404 700161
rect 234804 700096 234832 700160
rect 234896 700096 234912 700160
rect 234976 700096 234992 700160
rect 235056 700096 235072 700160
rect 235136 700096 235152 700160
rect 235216 700096 235232 700160
rect 235296 700096 235312 700160
rect 235376 700096 235404 700160
rect 234804 700095 235404 700096
rect 270804 700160 271404 700161
rect 270804 700096 270832 700160
rect 270896 700096 270912 700160
rect 270976 700096 270992 700160
rect 271056 700096 271072 700160
rect 271136 700096 271152 700160
rect 271216 700096 271232 700160
rect 271296 700096 271312 700160
rect 271376 700096 271404 700160
rect 270804 700095 271404 700096
rect 306804 700160 307404 700161
rect 306804 700096 306832 700160
rect 306896 700096 306912 700160
rect 306976 700096 306992 700160
rect 307056 700096 307072 700160
rect 307136 700096 307152 700160
rect 307216 700096 307232 700160
rect 307296 700096 307312 700160
rect 307376 700096 307404 700160
rect 306804 700095 307404 700096
rect 342804 700160 343404 700161
rect 342804 700096 342832 700160
rect 342896 700096 342912 700160
rect 342976 700096 342992 700160
rect 343056 700096 343072 700160
rect 343136 700096 343152 700160
rect 343216 700096 343232 700160
rect 343296 700096 343312 700160
rect 343376 700096 343404 700160
rect 342804 700095 343404 700096
rect 378804 700160 379404 700161
rect 378804 700096 378832 700160
rect 378896 700096 378912 700160
rect 378976 700096 378992 700160
rect 379056 700096 379072 700160
rect 379136 700096 379152 700160
rect 379216 700096 379232 700160
rect 379296 700096 379312 700160
rect 379376 700096 379404 700160
rect 378804 700095 379404 700096
rect 414804 700160 415404 700161
rect 414804 700096 414832 700160
rect 414896 700096 414912 700160
rect 414976 700096 414992 700160
rect 415056 700096 415072 700160
rect 415136 700096 415152 700160
rect 415216 700096 415232 700160
rect 415296 700096 415312 700160
rect 415376 700096 415404 700160
rect 414804 700095 415404 700096
rect 450804 700160 451404 700161
rect 450804 700096 450832 700160
rect 450896 700096 450912 700160
rect 450976 700096 450992 700160
rect 451056 700096 451072 700160
rect 451136 700096 451152 700160
rect 451216 700096 451232 700160
rect 451296 700096 451312 700160
rect 451376 700096 451404 700160
rect 450804 700095 451404 700096
rect 486804 700160 487404 700161
rect 486804 700096 486832 700160
rect 486896 700096 486912 700160
rect 486976 700096 486992 700160
rect 487056 700096 487072 700160
rect 487136 700096 487152 700160
rect 487216 700096 487232 700160
rect 487296 700096 487312 700160
rect 487376 700096 487404 700160
rect 486804 700095 487404 700096
rect 522804 700160 523404 700161
rect 522804 700096 522832 700160
rect 522896 700096 522912 700160
rect 522976 700096 522992 700160
rect 523056 700096 523072 700160
rect 523136 700096 523152 700160
rect 523216 700096 523232 700160
rect 523296 700096 523312 700160
rect 523376 700096 523404 700160
rect 522804 700095 523404 700096
rect 558804 700160 559404 700161
rect 558804 700096 558832 700160
rect 558896 700096 558912 700160
rect 558976 700096 558992 700160
rect 559056 700096 559072 700160
rect 559136 700096 559152 700160
rect 559216 700096 559232 700160
rect 559296 700096 559312 700160
rect 559376 700096 559404 700160
rect 558804 700095 559404 700096
rect 244181 700090 244247 700093
rect 251081 700090 251147 700093
rect 244181 700088 251147 700090
rect 244181 700032 244186 700088
rect 244242 700032 251086 700088
rect 251142 700032 251147 700088
rect 244181 700030 251147 700032
rect 244181 700027 244247 700030
rect 251081 700027 251147 700030
rect 280061 700090 280127 700093
rect 289537 700090 289603 700093
rect 280061 700088 289603 700090
rect 280061 700032 280066 700088
rect 280122 700032 289542 700088
rect 289598 700032 289603 700088
rect 280061 700030 289603 700032
rect 280061 700027 280127 700030
rect 289537 700027 289603 700030
rect 292297 699954 292363 699957
rect 292665 699954 292731 699957
rect 292297 699952 292731 699954
rect 292297 699896 292302 699952
rect 292358 699896 292670 699952
rect 292726 699896 292731 699952
rect 292297 699894 292731 699896
rect 292297 699891 292363 699894
rect 292665 699891 292731 699894
rect 302049 699954 302115 699957
rect 303613 699954 303679 699957
rect 302049 699952 303679 699954
rect 302049 699896 302054 699952
rect 302110 699896 303618 699952
rect 303674 699896 303679 699952
rect 302049 699894 303679 699896
rect 302049 699891 302115 699894
rect 303613 699891 303679 699894
rect 270493 699818 270559 699821
rect 273161 699818 273227 699821
rect 270493 699816 273227 699818
rect 270493 699760 270498 699816
rect 270554 699760 273166 699816
rect 273222 699760 273227 699816
rect 270493 699758 273227 699760
rect 270493 699755 270559 699758
rect 273161 699755 273227 699758
rect 292481 699818 292547 699821
rect 301957 699818 302023 699821
rect 292481 699816 302023 699818
rect 292481 699760 292486 699816
rect 292542 699760 301962 699816
rect 302018 699760 302023 699816
rect 292481 699758 302023 699760
rect 292481 699755 292547 699758
rect 301957 699755 302023 699758
rect 241513 699682 241579 699685
rect 251081 699682 251147 699685
rect 241513 699680 251147 699682
rect 241513 699624 241518 699680
rect 241574 699624 251086 699680
rect 251142 699624 251147 699680
rect 241513 699622 251147 699624
rect 241513 699619 241579 699622
rect 251081 699619 251147 699622
rect 36804 699616 37404 699617
rect 36804 699552 36832 699616
rect 36896 699552 36912 699616
rect 36976 699552 36992 699616
rect 37056 699552 37072 699616
rect 37136 699552 37152 699616
rect 37216 699552 37232 699616
rect 37296 699552 37312 699616
rect 37376 699552 37404 699616
rect 36804 699551 37404 699552
rect 72804 699616 73404 699617
rect 72804 699552 72832 699616
rect 72896 699552 72912 699616
rect 72976 699552 72992 699616
rect 73056 699552 73072 699616
rect 73136 699552 73152 699616
rect 73216 699552 73232 699616
rect 73296 699552 73312 699616
rect 73376 699552 73404 699616
rect 72804 699551 73404 699552
rect 108804 699616 109404 699617
rect 108804 699552 108832 699616
rect 108896 699552 108912 699616
rect 108976 699552 108992 699616
rect 109056 699552 109072 699616
rect 109136 699552 109152 699616
rect 109216 699552 109232 699616
rect 109296 699552 109312 699616
rect 109376 699552 109404 699616
rect 108804 699551 109404 699552
rect 144804 699616 145404 699617
rect 144804 699552 144832 699616
rect 144896 699552 144912 699616
rect 144976 699552 144992 699616
rect 145056 699552 145072 699616
rect 145136 699552 145152 699616
rect 145216 699552 145232 699616
rect 145296 699552 145312 699616
rect 145376 699552 145404 699616
rect 144804 699551 145404 699552
rect 180804 699616 181404 699617
rect 180804 699552 180832 699616
rect 180896 699552 180912 699616
rect 180976 699552 180992 699616
rect 181056 699552 181072 699616
rect 181136 699552 181152 699616
rect 181216 699552 181232 699616
rect 181296 699552 181312 699616
rect 181376 699552 181404 699616
rect 180804 699551 181404 699552
rect 216804 699616 217404 699617
rect 216804 699552 216832 699616
rect 216896 699552 216912 699616
rect 216976 699552 216992 699616
rect 217056 699552 217072 699616
rect 217136 699552 217152 699616
rect 217216 699552 217232 699616
rect 217296 699552 217312 699616
rect 217376 699552 217404 699616
rect 216804 699551 217404 699552
rect 252804 699616 253404 699617
rect 252804 699552 252832 699616
rect 252896 699552 252912 699616
rect 252976 699552 252992 699616
rect 253056 699552 253072 699616
rect 253136 699552 253152 699616
rect 253216 699552 253232 699616
rect 253296 699552 253312 699616
rect 253376 699552 253404 699616
rect 252804 699551 253404 699552
rect 288804 699616 289404 699617
rect 288804 699552 288832 699616
rect 288896 699552 288912 699616
rect 288976 699552 288992 699616
rect 289056 699552 289072 699616
rect 289136 699552 289152 699616
rect 289216 699552 289232 699616
rect 289296 699552 289312 699616
rect 289376 699552 289404 699616
rect 288804 699551 289404 699552
rect 324804 699616 325404 699617
rect 324804 699552 324832 699616
rect 324896 699552 324912 699616
rect 324976 699552 324992 699616
rect 325056 699552 325072 699616
rect 325136 699552 325152 699616
rect 325216 699552 325232 699616
rect 325296 699552 325312 699616
rect 325376 699552 325404 699616
rect 324804 699551 325404 699552
rect 360804 699616 361404 699617
rect 360804 699552 360832 699616
rect 360896 699552 360912 699616
rect 360976 699552 360992 699616
rect 361056 699552 361072 699616
rect 361136 699552 361152 699616
rect 361216 699552 361232 699616
rect 361296 699552 361312 699616
rect 361376 699552 361404 699616
rect 360804 699551 361404 699552
rect 396804 699616 397404 699617
rect 396804 699552 396832 699616
rect 396896 699552 396912 699616
rect 396976 699552 396992 699616
rect 397056 699552 397072 699616
rect 397136 699552 397152 699616
rect 397216 699552 397232 699616
rect 397296 699552 397312 699616
rect 397376 699552 397404 699616
rect 396804 699551 397404 699552
rect 432804 699616 433404 699617
rect 432804 699552 432832 699616
rect 432896 699552 432912 699616
rect 432976 699552 432992 699616
rect 433056 699552 433072 699616
rect 433136 699552 433152 699616
rect 433216 699552 433232 699616
rect 433296 699552 433312 699616
rect 433376 699552 433404 699616
rect 432804 699551 433404 699552
rect 468804 699616 469404 699617
rect 468804 699552 468832 699616
rect 468896 699552 468912 699616
rect 468976 699552 468992 699616
rect 469056 699552 469072 699616
rect 469136 699552 469152 699616
rect 469216 699552 469232 699616
rect 469296 699552 469312 699616
rect 469376 699552 469404 699616
rect 468804 699551 469404 699552
rect 504804 699616 505404 699617
rect 504804 699552 504832 699616
rect 504896 699552 504912 699616
rect 504976 699552 504992 699616
rect 505056 699552 505072 699616
rect 505136 699552 505152 699616
rect 505216 699552 505232 699616
rect 505296 699552 505312 699616
rect 505376 699552 505404 699616
rect 504804 699551 505404 699552
rect 540804 699616 541404 699617
rect 540804 699552 540832 699616
rect 540896 699552 540912 699616
rect 540976 699552 540992 699616
rect 541056 699552 541072 699616
rect 541136 699552 541152 699616
rect 541216 699552 541232 699616
rect 541296 699552 541312 699616
rect 541376 699552 541404 699616
rect 540804 699551 541404 699552
rect 576804 699616 577404 699617
rect 576804 699552 576832 699616
rect 576896 699552 576912 699616
rect 576976 699552 576992 699616
rect 577056 699552 577072 699616
rect 577136 699552 577152 699616
rect 577216 699552 577232 699616
rect 577296 699552 577312 699616
rect 577376 699552 577404 699616
rect 576804 699551 577404 699552
rect 263593 699546 263659 699549
rect 282729 699546 282795 699549
rect 263593 699544 282795 699546
rect 263593 699488 263598 699544
rect 263654 699488 282734 699544
rect 282790 699488 282795 699544
rect 263593 699486 282795 699488
rect 263593 699483 263659 699486
rect 282729 699483 282795 699486
rect 282913 699546 282979 699549
rect 289721 699546 289787 699549
rect 292665 699546 292731 699549
rect 282913 699544 283298 699546
rect 282913 699488 282918 699544
rect 282974 699488 283298 699544
rect 282913 699486 283298 699488
rect 282913 699483 282979 699486
rect 190453 699410 190519 699413
rect 200021 699410 200087 699413
rect 190453 699408 200087 699410
rect 190453 699352 190458 699408
rect 190514 699352 200026 699408
rect 200082 699352 200087 699408
rect 190453 699350 200087 699352
rect 190453 699347 190519 699350
rect 200021 699347 200087 699350
rect 229093 699410 229159 699413
rect 244181 699410 244247 699413
rect 229093 699408 244247 699410
rect 229093 699352 229098 699408
rect 229154 699352 244186 699408
rect 244242 699352 244247 699408
rect 229093 699350 244247 699352
rect 229093 699347 229159 699350
rect 244181 699347 244247 699350
rect 263685 699410 263751 699413
rect 273345 699410 273411 699413
rect 263685 699408 273411 699410
rect 263685 699352 263690 699408
rect 263746 699352 273350 699408
rect 273406 699352 273411 699408
rect 263685 699350 273411 699352
rect 263685 699347 263751 699350
rect 273345 699347 273411 699350
rect 282729 699410 282795 699413
rect 283005 699410 283071 699413
rect 282729 699408 283071 699410
rect 282729 699352 282734 699408
rect 282790 699352 283010 699408
rect 283066 699352 283071 699408
rect 282729 699350 283071 699352
rect 283238 699410 283298 699486
rect 289721 699544 292731 699546
rect 289721 699488 289726 699544
rect 289782 699488 292670 699544
rect 292726 699488 292731 699544
rect 289721 699486 292731 699488
rect 289721 699483 289787 699486
rect 292665 699483 292731 699486
rect 294045 699410 294111 699413
rect 283238 699408 294111 699410
rect 283238 699352 294050 699408
rect 294106 699352 294111 699408
rect 283238 699350 294111 699352
rect 282729 699347 282795 699350
rect 283005 699347 283071 699350
rect 294045 699347 294111 699350
rect 4797 699274 4863 699277
rect 530945 699274 531011 699277
rect 4797 699272 531011 699274
rect 4797 699216 4802 699272
rect 4858 699216 530950 699272
rect 531006 699216 531011 699272
rect 4797 699214 531011 699216
rect 4797 699211 4863 699214
rect 530945 699211 531011 699214
rect 180793 699138 180859 699141
rect 190361 699138 190427 699141
rect 180793 699136 190427 699138
rect 180793 699080 180798 699136
rect 180854 699080 190366 699136
rect 190422 699080 190427 699136
rect 180793 699078 190427 699080
rect 180793 699075 180859 699078
rect 190361 699075 190427 699078
rect 209773 699138 209839 699141
rect 219341 699138 219407 699141
rect 209773 699136 219407 699138
rect 209773 699080 209778 699136
rect 209834 699080 219346 699136
rect 219402 699080 219407 699136
rect 209773 699078 219407 699080
rect 209773 699075 209839 699078
rect 219341 699075 219407 699078
rect 253657 699138 253723 699141
rect 263685 699138 263751 699141
rect 253657 699136 263751 699138
rect 253657 699080 253662 699136
rect 253718 699080 263690 699136
rect 263746 699080 263751 699136
rect 253657 699078 263751 699080
rect 253657 699075 253723 699078
rect 263685 699075 263751 699078
rect 273253 699138 273319 699141
rect 282862 699138 282868 699140
rect 273253 699136 282868 699138
rect 273253 699080 273258 699136
rect 273314 699080 282868 699136
rect 273253 699078 282868 699080
rect 273253 699075 273319 699078
rect 282862 699076 282868 699078
rect 282932 699076 282938 699140
rect 288433 699138 288499 699141
rect 283054 699136 288499 699138
rect 283054 699080 288438 699136
rect 288494 699080 288499 699136
rect 283054 699078 288499 699080
rect 18804 699072 19404 699073
rect 18804 699008 18832 699072
rect 18896 699008 18912 699072
rect 18976 699008 18992 699072
rect 19056 699008 19072 699072
rect 19136 699008 19152 699072
rect 19216 699008 19232 699072
rect 19296 699008 19312 699072
rect 19376 699008 19404 699072
rect 18804 699007 19404 699008
rect 54804 699072 55404 699073
rect 54804 699008 54832 699072
rect 54896 699008 54912 699072
rect 54976 699008 54992 699072
rect 55056 699008 55072 699072
rect 55136 699008 55152 699072
rect 55216 699008 55232 699072
rect 55296 699008 55312 699072
rect 55376 699008 55404 699072
rect 54804 699007 55404 699008
rect 90804 699072 91404 699073
rect 90804 699008 90832 699072
rect 90896 699008 90912 699072
rect 90976 699008 90992 699072
rect 91056 699008 91072 699072
rect 91136 699008 91152 699072
rect 91216 699008 91232 699072
rect 91296 699008 91312 699072
rect 91376 699008 91404 699072
rect 90804 699007 91404 699008
rect 126804 699072 127404 699073
rect 126804 699008 126832 699072
rect 126896 699008 126912 699072
rect 126976 699008 126992 699072
rect 127056 699008 127072 699072
rect 127136 699008 127152 699072
rect 127216 699008 127232 699072
rect 127296 699008 127312 699072
rect 127376 699008 127404 699072
rect 126804 699007 127404 699008
rect 162804 699072 163404 699073
rect 162804 699008 162832 699072
rect 162896 699008 162912 699072
rect 162976 699008 162992 699072
rect 163056 699008 163072 699072
rect 163136 699008 163152 699072
rect 163216 699008 163232 699072
rect 163296 699008 163312 699072
rect 163376 699008 163404 699072
rect 162804 699007 163404 699008
rect 198804 699072 199404 699073
rect 198804 699008 198832 699072
rect 198896 699008 198912 699072
rect 198976 699008 198992 699072
rect 199056 699008 199072 699072
rect 199136 699008 199152 699072
rect 199216 699008 199232 699072
rect 199296 699008 199312 699072
rect 199376 699008 199404 699072
rect 198804 699007 199404 699008
rect 234804 699072 235404 699073
rect 234804 699008 234832 699072
rect 234896 699008 234912 699072
rect 234976 699008 234992 699072
rect 235056 699008 235072 699072
rect 235136 699008 235152 699072
rect 235216 699008 235232 699072
rect 235296 699008 235312 699072
rect 235376 699008 235404 699072
rect 234804 699007 235404 699008
rect 270804 699072 271404 699073
rect 270804 699008 270832 699072
rect 270896 699008 270912 699072
rect 270976 699008 270992 699072
rect 271056 699008 271072 699072
rect 271136 699008 271152 699072
rect 271216 699008 271232 699072
rect 271296 699008 271312 699072
rect 271376 699008 271404 699072
rect 270804 699007 271404 699008
rect 244089 699002 244155 699005
rect 253841 699002 253907 699005
rect 244089 699000 253907 699002
rect 244089 698944 244094 699000
rect 244150 698944 253846 699000
rect 253902 698944 253907 699000
rect 244089 698942 253907 698944
rect 244089 698939 244155 698942
rect 253841 698939 253907 698942
rect 261385 699002 261451 699005
rect 263869 699002 263935 699005
rect 261385 699000 263935 699002
rect 261385 698944 261390 699000
rect 261446 698944 263874 699000
rect 263930 698944 263935 699000
rect 261385 698942 263935 698944
rect 261385 698939 261451 698942
rect 263869 698939 263935 698942
rect 273529 699002 273595 699005
rect 283054 699002 283114 699078
rect 288433 699075 288499 699078
rect 292389 699138 292455 699141
rect 302141 699138 302207 699141
rect 292389 699136 302207 699138
rect 292389 699080 292394 699136
rect 292450 699080 302146 699136
rect 302202 699080 302207 699136
rect 292389 699078 302207 699080
rect 292389 699075 292455 699078
rect 302141 699075 302207 699078
rect 311893 699138 311959 699141
rect 325509 699138 325575 699141
rect 311893 699136 325575 699138
rect 311893 699080 311898 699136
rect 311954 699080 325514 699136
rect 325570 699080 325575 699136
rect 311893 699078 325575 699080
rect 311893 699075 311959 699078
rect 325509 699075 325575 699078
rect 325693 699138 325759 699141
rect 331213 699138 331279 699141
rect 325693 699136 331279 699138
rect 325693 699080 325698 699136
rect 325754 699080 331218 699136
rect 331274 699080 331279 699136
rect 325693 699078 331279 699080
rect 325693 699075 325759 699078
rect 331213 699075 331279 699078
rect 343541 699138 343607 699141
rect 354489 699138 354555 699141
rect 343541 699136 354555 699138
rect 343541 699080 343546 699136
rect 343602 699080 354494 699136
rect 354550 699080 354555 699136
rect 343541 699078 354555 699080
rect 343541 699075 343607 699078
rect 354489 699075 354555 699078
rect 306804 699072 307404 699073
rect 306804 699008 306832 699072
rect 306896 699008 306912 699072
rect 306976 699008 306992 699072
rect 307056 699008 307072 699072
rect 307136 699008 307152 699072
rect 307216 699008 307232 699072
rect 307296 699008 307312 699072
rect 307376 699008 307404 699072
rect 306804 699007 307404 699008
rect 342804 699072 343404 699073
rect 342804 699008 342832 699072
rect 342896 699008 342912 699072
rect 342976 699008 342992 699072
rect 343056 699008 343072 699072
rect 343136 699008 343152 699072
rect 343216 699008 343232 699072
rect 343296 699008 343312 699072
rect 343376 699008 343404 699072
rect 342804 699007 343404 699008
rect 378804 699072 379404 699073
rect 378804 699008 378832 699072
rect 378896 699008 378912 699072
rect 378976 699008 378992 699072
rect 379056 699008 379072 699072
rect 379136 699008 379152 699072
rect 379216 699008 379232 699072
rect 379296 699008 379312 699072
rect 379376 699008 379404 699072
rect 378804 699007 379404 699008
rect 414804 699072 415404 699073
rect 414804 699008 414832 699072
rect 414896 699008 414912 699072
rect 414976 699008 414992 699072
rect 415056 699008 415072 699072
rect 415136 699008 415152 699072
rect 415216 699008 415232 699072
rect 415296 699008 415312 699072
rect 415376 699008 415404 699072
rect 414804 699007 415404 699008
rect 450804 699072 451404 699073
rect 450804 699008 450832 699072
rect 450896 699008 450912 699072
rect 450976 699008 450992 699072
rect 451056 699008 451072 699072
rect 451136 699008 451152 699072
rect 451216 699008 451232 699072
rect 451296 699008 451312 699072
rect 451376 699008 451404 699072
rect 450804 699007 451404 699008
rect 486804 699072 487404 699073
rect 486804 699008 486832 699072
rect 486896 699008 486912 699072
rect 486976 699008 486992 699072
rect 487056 699008 487072 699072
rect 487136 699008 487152 699072
rect 487216 699008 487232 699072
rect 487296 699008 487312 699072
rect 487376 699008 487404 699072
rect 486804 699007 487404 699008
rect 522804 699072 523404 699073
rect 522804 699008 522832 699072
rect 522896 699008 522912 699072
rect 522976 699008 522992 699072
rect 523056 699008 523072 699072
rect 523136 699008 523152 699072
rect 523216 699008 523232 699072
rect 523296 699008 523312 699072
rect 523376 699008 523404 699072
rect 522804 699007 523404 699008
rect 558804 699072 559404 699073
rect 558804 699008 558832 699072
rect 558896 699008 558912 699072
rect 558976 699008 558992 699072
rect 559056 699008 559072 699072
rect 559136 699008 559152 699072
rect 559216 699008 559232 699072
rect 559296 699008 559312 699072
rect 559376 699008 559404 699072
rect 558804 699007 559404 699008
rect 273529 699000 283114 699002
rect 273529 698944 273534 699000
rect 273590 698944 283114 699000
rect 273529 698942 283114 698944
rect 283281 699002 283347 699005
rect 292481 699002 292547 699005
rect 283281 699000 292547 699002
rect 283281 698944 283286 699000
rect 283342 698944 292486 699000
rect 292542 698944 292547 699000
rect 283281 698942 292547 698944
rect 273529 698939 273595 698942
rect 283281 698939 283347 698942
rect 292481 698939 292547 698942
rect 43437 698866 43503 698869
rect 86718 698866 86724 698868
rect 43437 698864 86724 698866
rect 43437 698808 43442 698864
rect 43498 698808 86724 698864
rect 43437 698806 86724 698808
rect 43437 698803 43503 698806
rect 86718 698804 86724 698806
rect 86788 698804 86794 698868
rect 233049 698866 233115 698869
rect 234705 698866 234771 698869
rect 233049 698864 234771 698866
rect 233049 698808 233054 698864
rect 233110 698808 234710 698864
rect 234766 698808 234771 698864
rect 233049 698806 234771 698808
rect 233049 698803 233115 698806
rect 234705 698803 234771 698806
rect 253749 698866 253815 698869
rect 263685 698866 263751 698869
rect 253749 698864 263751 698866
rect 253749 698808 253754 698864
rect 253810 698808 263690 698864
rect 263746 698808 263751 698864
rect 253749 698806 263751 698808
rect 253749 698803 253815 698806
rect 263685 698803 263751 698806
rect 282913 698866 282979 698869
rect 300209 698866 300275 698869
rect 282913 698864 300275 698866
rect 282913 698808 282918 698864
rect 282974 698808 300214 698864
rect 300270 698808 300275 698864
rect 282913 698806 300275 698808
rect 282913 698803 282979 698806
rect 300209 698803 300275 698806
rect 306373 698866 306439 698869
rect 325601 698866 325667 698869
rect 306373 698864 325667 698866
rect 306373 698808 306378 698864
rect 306434 698808 325606 698864
rect 325662 698808 325667 698864
rect 306373 698806 325667 698808
rect 306373 698803 306439 698806
rect 325601 698803 325667 698806
rect 340689 698866 340755 698869
rect 354581 698866 354647 698869
rect 340689 698864 354647 698866
rect 340689 698808 340694 698864
rect 340750 698808 354586 698864
rect 354642 698808 354647 698864
rect 340689 698806 354647 698808
rect 340689 698803 340755 698806
rect 354581 698803 354647 698806
rect 447174 698804 447180 698868
rect 447244 698866 447250 698868
rect 526253 698866 526319 698869
rect 447244 698864 526319 698866
rect 447244 698808 526258 698864
rect 526314 698808 526319 698864
rect 447244 698806 526319 698808
rect 447244 698804 447250 698806
rect 526253 698803 526319 698806
rect 5349 698730 5415 698733
rect 516777 698730 516843 698733
rect 5349 698728 516843 698730
rect 5349 698672 5354 698728
rect 5410 698672 516782 698728
rect 516838 698672 516843 698728
rect 5349 698670 516843 698672
rect 5349 698667 5415 698670
rect 516777 698667 516843 698670
rect 282862 698532 282868 698596
rect 282932 698594 282938 698596
rect 283005 698594 283071 698597
rect 282932 698592 283071 698594
rect 282932 698536 283010 698592
rect 283066 698536 283071 698592
rect 282932 698534 283071 698536
rect 282932 698532 282938 698534
rect 283005 698531 283071 698534
rect 36804 698528 37404 698529
rect 36804 698464 36832 698528
rect 36896 698464 36912 698528
rect 36976 698464 36992 698528
rect 37056 698464 37072 698528
rect 37136 698464 37152 698528
rect 37216 698464 37232 698528
rect 37296 698464 37312 698528
rect 37376 698464 37404 698528
rect 36804 698463 37404 698464
rect 72804 698528 73404 698529
rect 72804 698464 72832 698528
rect 72896 698464 72912 698528
rect 72976 698464 72992 698528
rect 73056 698464 73072 698528
rect 73136 698464 73152 698528
rect 73216 698464 73232 698528
rect 73296 698464 73312 698528
rect 73376 698464 73404 698528
rect 72804 698463 73404 698464
rect 108804 698528 109404 698529
rect 108804 698464 108832 698528
rect 108896 698464 108912 698528
rect 108976 698464 108992 698528
rect 109056 698464 109072 698528
rect 109136 698464 109152 698528
rect 109216 698464 109232 698528
rect 109296 698464 109312 698528
rect 109376 698464 109404 698528
rect 108804 698463 109404 698464
rect 144804 698528 145404 698529
rect 144804 698464 144832 698528
rect 144896 698464 144912 698528
rect 144976 698464 144992 698528
rect 145056 698464 145072 698528
rect 145136 698464 145152 698528
rect 145216 698464 145232 698528
rect 145296 698464 145312 698528
rect 145376 698464 145404 698528
rect 144804 698463 145404 698464
rect 180804 698528 181404 698529
rect 180804 698464 180832 698528
rect 180896 698464 180912 698528
rect 180976 698464 180992 698528
rect 181056 698464 181072 698528
rect 181136 698464 181152 698528
rect 181216 698464 181232 698528
rect 181296 698464 181312 698528
rect 181376 698464 181404 698528
rect 180804 698463 181404 698464
rect 216804 698528 217404 698529
rect 216804 698464 216832 698528
rect 216896 698464 216912 698528
rect 216976 698464 216992 698528
rect 217056 698464 217072 698528
rect 217136 698464 217152 698528
rect 217216 698464 217232 698528
rect 217296 698464 217312 698528
rect 217376 698464 217404 698528
rect 216804 698463 217404 698464
rect 252804 698528 253404 698529
rect 252804 698464 252832 698528
rect 252896 698464 252912 698528
rect 252976 698464 252992 698528
rect 253056 698464 253072 698528
rect 253136 698464 253152 698528
rect 253216 698464 253232 698528
rect 253296 698464 253312 698528
rect 253376 698464 253404 698528
rect 252804 698463 253404 698464
rect 288804 698528 289404 698529
rect 288804 698464 288832 698528
rect 288896 698464 288912 698528
rect 288976 698464 288992 698528
rect 289056 698464 289072 698528
rect 289136 698464 289152 698528
rect 289216 698464 289232 698528
rect 289296 698464 289312 698528
rect 289376 698464 289404 698528
rect 288804 698463 289404 698464
rect 324804 698528 325404 698529
rect 324804 698464 324832 698528
rect 324896 698464 324912 698528
rect 324976 698464 324992 698528
rect 325056 698464 325072 698528
rect 325136 698464 325152 698528
rect 325216 698464 325232 698528
rect 325296 698464 325312 698528
rect 325376 698464 325404 698528
rect 324804 698463 325404 698464
rect 360804 698528 361404 698529
rect 360804 698464 360832 698528
rect 360896 698464 360912 698528
rect 360976 698464 360992 698528
rect 361056 698464 361072 698528
rect 361136 698464 361152 698528
rect 361216 698464 361232 698528
rect 361296 698464 361312 698528
rect 361376 698464 361404 698528
rect 360804 698463 361404 698464
rect 396804 698528 397404 698529
rect 396804 698464 396832 698528
rect 396896 698464 396912 698528
rect 396976 698464 396992 698528
rect 397056 698464 397072 698528
rect 397136 698464 397152 698528
rect 397216 698464 397232 698528
rect 397296 698464 397312 698528
rect 397376 698464 397404 698528
rect 396804 698463 397404 698464
rect 432804 698528 433404 698529
rect 432804 698464 432832 698528
rect 432896 698464 432912 698528
rect 432976 698464 432992 698528
rect 433056 698464 433072 698528
rect 433136 698464 433152 698528
rect 433216 698464 433232 698528
rect 433296 698464 433312 698528
rect 433376 698464 433404 698528
rect 432804 698463 433404 698464
rect 468804 698528 469404 698529
rect 468804 698464 468832 698528
rect 468896 698464 468912 698528
rect 468976 698464 468992 698528
rect 469056 698464 469072 698528
rect 469136 698464 469152 698528
rect 469216 698464 469232 698528
rect 469296 698464 469312 698528
rect 469376 698464 469404 698528
rect 468804 698463 469404 698464
rect 504804 698528 505404 698529
rect 504804 698464 504832 698528
rect 504896 698464 504912 698528
rect 504976 698464 504992 698528
rect 505056 698464 505072 698528
rect 505136 698464 505152 698528
rect 505216 698464 505232 698528
rect 505296 698464 505312 698528
rect 505376 698464 505404 698528
rect 504804 698463 505404 698464
rect 540804 698528 541404 698529
rect 540804 698464 540832 698528
rect 540896 698464 540912 698528
rect 540976 698464 540992 698528
rect 541056 698464 541072 698528
rect 541136 698464 541152 698528
rect 541216 698464 541232 698528
rect 541296 698464 541312 698528
rect 541376 698464 541404 698528
rect 540804 698463 541404 698464
rect 576804 698528 577404 698529
rect 576804 698464 576832 698528
rect 576896 698464 576912 698528
rect 576976 698464 576992 698528
rect 577056 698464 577072 698528
rect 577136 698464 577152 698528
rect 577216 698464 577232 698528
rect 577296 698464 577312 698528
rect 577376 698464 577404 698528
rect 576804 698463 577404 698464
rect 29177 698322 29243 698325
rect 71814 698322 71820 698324
rect 29177 698320 71820 698322
rect 29177 698264 29182 698320
rect 29238 698264 71820 698320
rect 29177 698262 71820 698264
rect 29177 698259 29243 698262
rect 71814 698260 71820 698262
rect 71884 698260 71890 698324
rect 579613 698050 579679 698053
rect 583520 698050 584960 698140
rect 579613 698048 584960 698050
rect 579613 697992 579618 698048
rect 579674 697992 584960 698048
rect 579613 697990 584960 697992
rect 579613 697987 579679 697990
rect 583520 697900 584960 697990
rect 6177 697098 6243 697101
rect 540421 697098 540487 697101
rect 6177 697096 540487 697098
rect 6177 697040 6182 697096
rect 6238 697040 540426 697096
rect 540482 697040 540487 697096
rect 6177 697038 540487 697040
rect 6177 697035 6243 697038
rect 540421 697035 540487 697038
rect 10317 696962 10383 696965
rect 574737 696962 574803 696965
rect 10317 696960 574803 696962
rect 10317 696904 10322 696960
rect 10378 696904 574742 696960
rect 574798 696904 574803 696960
rect 10317 696902 574803 696904
rect 10317 696899 10383 696902
rect 574737 696899 574803 696902
rect -960 696540 480 696780
rect 173893 696010 173959 696013
rect 174261 696010 174327 696013
rect 173893 696008 174327 696010
rect 173893 695952 173898 696008
rect 173954 695952 174266 696008
rect 174322 695952 174327 696008
rect 173893 695950 174327 695952
rect 173893 695947 173959 695950
rect 174261 695947 174327 695950
rect 509509 695874 509575 695877
rect 518065 695874 518131 695877
rect 509509 695872 518131 695874
rect 509509 695816 509514 695872
rect 509570 695816 518070 695872
rect 518126 695816 518131 695872
rect 509509 695814 518131 695816
rect 509509 695811 509575 695814
rect 518065 695811 518131 695814
rect 3417 695738 3483 695741
rect 545021 695738 545087 695741
rect 3417 695736 545087 695738
rect 3417 695680 3422 695736
rect 3478 695680 545026 695736
rect 545082 695680 545087 695736
rect 3417 695678 545087 695680
rect 3417 695675 3483 695678
rect 545021 695675 545087 695678
rect 19977 695602 20043 695605
rect 509509 695602 509575 695605
rect 19977 695600 509575 695602
rect 19977 695544 19982 695600
rect 20038 695544 509514 695600
rect 509570 695544 509575 695600
rect 19977 695542 509575 695544
rect 19977 695539 20043 695542
rect 509509 695539 509575 695542
rect 518065 695602 518131 695605
rect 576117 695602 576183 695605
rect 518065 695600 576183 695602
rect 518065 695544 518070 695600
rect 518126 695544 576122 695600
rect 576178 695544 576183 695600
rect 518065 695542 576183 695544
rect 518065 695539 518131 695542
rect 576117 695539 576183 695542
rect 15285 695332 15351 695333
rect 15285 695330 15332 695332
rect 15240 695328 15332 695330
rect 15240 695272 15290 695328
rect 15240 695270 15332 695272
rect 15285 695268 15332 695270
rect 15396 695268 15402 695332
rect 176193 695330 176259 695333
rect 521377 695332 521443 695333
rect 179638 695330 179644 695332
rect 176193 695328 179644 695330
rect 176193 695272 176198 695328
rect 176254 695272 179644 695328
rect 176193 695270 179644 695272
rect 15285 695267 15351 695268
rect 176193 695267 176259 695270
rect 179638 695268 179644 695270
rect 179708 695268 179714 695332
rect 521326 695330 521332 695332
rect 521286 695270 521332 695330
rect 521396 695328 521443 695332
rect 521438 695272 521443 695328
rect 521326 695268 521332 695270
rect 521396 695268 521443 695272
rect 521377 695267 521443 695268
rect 231894 694996 231900 695060
rect 231964 695058 231970 695060
rect 236862 695058 236868 695060
rect 231964 694998 236868 695058
rect 231964 694996 231970 694998
rect 236862 694996 236868 694998
rect 236932 694996 236938 695060
rect 251214 694996 251220 695060
rect 251284 695058 251290 695060
rect 256182 695058 256188 695060
rect 251284 694998 256188 695058
rect 251284 694996 251290 694998
rect 256182 694996 256188 694998
rect 256252 694996 256258 695060
rect 357382 694996 357388 695060
rect 357452 695058 357458 695060
rect 362166 695058 362172 695060
rect 357452 694998 362172 695058
rect 357452 694996 357458 694998
rect 362166 694996 362172 694998
rect 362236 694996 362242 695060
rect 434662 694996 434668 695060
rect 434732 695058 434738 695060
rect 439446 695058 439452 695060
rect 434732 694998 439452 695058
rect 434732 694996 434738 694998
rect 439446 694996 439452 694998
rect 439516 694996 439522 695060
rect 137318 694860 137324 694924
rect 137388 694922 137394 694924
rect 141918 694922 141924 694924
rect 137388 694862 141924 694922
rect 137388 694860 137394 694862
rect 141918 694860 141924 694862
rect 141988 694860 141994 694924
rect 196198 694860 196204 694924
rect 196268 694922 196274 694924
rect 202454 694922 202460 694924
rect 196268 694862 202460 694922
rect 196268 694860 196274 694862
rect 202454 694860 202460 694862
rect 202524 694860 202530 694924
rect 273110 694860 273116 694924
rect 273180 694922 273186 694924
rect 278814 694922 278820 694924
rect 273180 694862 278820 694922
rect 273180 694860 273186 694862
rect 278814 694860 278820 694862
rect 278884 694860 278890 694924
rect 280102 694860 280108 694924
rect 280172 694922 280178 694924
rect 283230 694922 283236 694924
rect 280172 694862 283236 694922
rect 280172 694860 280178 694862
rect 283230 694860 283236 694862
rect 283300 694860 283306 694924
rect 292798 694860 292804 694924
rect 292868 694922 292874 694924
rect 299054 694922 299060 694924
rect 292868 694862 299060 694922
rect 292868 694860 292874 694862
rect 299054 694860 299060 694862
rect 299124 694860 299130 694924
rect 346342 694860 346348 694924
rect 346412 694922 346418 694924
rect 351310 694922 351316 694924
rect 346412 694862 351316 694922
rect 346412 694860 346418 694862
rect 351310 694860 351316 694862
rect 351380 694860 351386 694924
rect 370078 694860 370084 694924
rect 370148 694922 370154 694924
rect 376334 694922 376340 694924
rect 370148 694862 376340 694922
rect 370148 694860 370154 694862
rect 376334 694860 376340 694862
rect 376404 694860 376410 694924
rect 389398 694860 389404 694924
rect 389468 694922 389474 694924
rect 395654 694922 395660 694924
rect 389468 694862 395660 694922
rect 389468 694860 389474 694862
rect 395654 694860 395660 694862
rect 395724 694860 395730 694924
rect 500902 694860 500908 694924
rect 500972 694922 500978 694924
rect 505686 694922 505692 694924
rect 500972 694862 505692 694922
rect 500972 694860 500978 694862
rect 505686 694860 505692 694862
rect 505756 694860 505762 694924
rect 134926 694724 134932 694788
rect 134996 694786 135002 694788
rect 138238 694786 138244 694788
rect 134996 694726 138244 694786
rect 134996 694724 135002 694726
rect 138238 694724 138244 694726
rect 138308 694724 138314 694788
rect 142102 694724 142108 694788
rect 142172 694786 142178 694788
rect 151670 694786 151676 694788
rect 142172 694726 151676 694786
rect 142172 694724 142178 694726
rect 151670 694724 151676 694726
rect 151740 694724 151746 694788
rect 152774 694724 152780 694788
rect 152844 694786 152850 694788
rect 159398 694786 159404 694788
rect 152844 694726 159404 694786
rect 152844 694724 152850 694726
rect 159398 694724 159404 694726
rect 159468 694724 159474 694788
rect 222142 694724 222148 694788
rect 222212 694786 222218 694788
rect 226926 694786 226932 694788
rect 222212 694726 226932 694786
rect 222212 694724 222218 694726
rect 226926 694724 226932 694726
rect 226996 694724 227002 694788
rect 236678 694786 236684 694788
rect 231902 694726 236684 694786
rect 106222 694588 106228 694652
rect 106292 694650 106298 694652
rect 115790 694650 115796 694652
rect 106292 694590 115796 694650
rect 106292 694588 106298 694590
rect 115790 694588 115796 694590
rect 115860 694588 115866 694652
rect 164182 694588 164188 694652
rect 164252 694650 164258 694652
rect 173566 694650 173572 694652
rect 164252 694590 173572 694650
rect 164252 694588 164258 694590
rect 173566 694588 173572 694590
rect 173636 694588 173642 694652
rect 176694 694588 176700 694652
rect 176764 694650 176770 694652
rect 176764 694590 177130 694650
rect 176764 694588 176770 694590
rect 15326 694452 15332 694516
rect 15396 694514 15402 694516
rect 15396 694454 24410 694514
rect 15396 694452 15402 694454
rect 24350 694378 24410 694454
rect 42006 694452 42012 694516
rect 42076 694514 42082 694516
rect 42076 694454 46858 694514
rect 42076 694452 42082 694454
rect 24350 694318 33794 694378
rect 9622 694180 9628 694244
rect 9692 694242 9698 694244
rect 33734 694242 33794 694318
rect 42006 694242 42012 694244
rect 9692 694182 19258 694242
rect 33734 694182 42012 694242
rect 9692 694180 9698 694182
rect 3509 693970 3575 693973
rect 9622 693970 9628 693972
rect 3509 693968 9628 693970
rect 3509 693912 3514 693968
rect 3570 693912 9628 693968
rect 3509 693910 9628 693912
rect 3509 693907 3575 693910
rect 9622 693908 9628 693910
rect 9692 693908 9698 693972
rect 19006 693908 19012 693972
rect 19076 693970 19082 693972
rect 19198 693970 19258 694182
rect 42006 694180 42012 694182
rect 42076 694180 42082 694244
rect 46798 694242 46858 694454
rect 85246 694452 85252 694516
rect 85316 694514 85322 694516
rect 85316 694454 98746 694514
rect 85316 694452 85322 694454
rect 79910 694378 79916 694380
rect 58022 694318 79916 694378
rect 58022 694242 58082 694318
rect 79910 694316 79916 694318
rect 79980 694316 79986 694380
rect 80094 694316 80100 694380
rect 80164 694378 80170 694380
rect 98310 694378 98316 694380
rect 80164 694318 98316 694378
rect 80164 694316 80170 694318
rect 98310 694316 98316 694318
rect 98380 694316 98386 694380
rect 46798 694182 58082 694242
rect 64822 694180 64828 694244
rect 64892 694242 64898 694244
rect 76966 694242 76972 694244
rect 64892 694182 76972 694242
rect 64892 694180 64898 694182
rect 76966 694180 76972 694182
rect 77036 694180 77042 694244
rect 86718 694180 86724 694244
rect 86788 694180 86794 694244
rect 37222 694044 37228 694108
rect 37292 694106 37298 694108
rect 41270 694106 41276 694108
rect 37292 694046 41276 694106
rect 37292 694044 37298 694046
rect 41270 694044 41276 694046
rect 41340 694044 41346 694108
rect 41454 694044 41460 694108
rect 41524 694106 41530 694108
rect 41524 694046 47042 694106
rect 41524 694044 41530 694046
rect 19076 693910 19258 693970
rect 19076 693908 19082 693910
rect 27286 693908 27292 693972
rect 27356 693970 27362 693972
rect 28942 693970 28948 693972
rect 27356 693910 28948 693970
rect 27356 693908 27362 693910
rect 28942 693908 28948 693910
rect 29012 693908 29018 693972
rect 46982 693970 47042 694046
rect 64822 693970 64828 693972
rect 46982 693910 64828 693970
rect 64822 693908 64828 693910
rect 64892 693908 64898 693972
rect 86726 693970 86786 694180
rect 98686 694106 98746 694454
rect 115974 694452 115980 694516
rect 116044 694514 116050 694516
rect 116044 694454 121010 694514
rect 116044 694452 116050 694454
rect 98862 694316 98868 694380
rect 98932 694378 98938 694380
rect 106222 694378 106228 694380
rect 98932 694318 106228 694378
rect 98932 694316 98938 694318
rect 106222 694316 106228 694318
rect 106292 694316 106298 694380
rect 106406 694316 106412 694380
rect 106476 694378 106482 694380
rect 120574 694378 120580 694380
rect 106476 694318 120580 694378
rect 106476 694316 106482 694318
rect 120574 694316 120580 694318
rect 120644 694316 120650 694380
rect 120950 694378 121010 694454
rect 130326 694452 130332 694516
rect 130396 694514 130402 694516
rect 134926 694514 134932 694516
rect 130396 694454 134932 694514
rect 130396 694452 130402 694454
rect 134926 694452 134932 694454
rect 134996 694452 135002 694516
rect 151670 694452 151676 694516
rect 151740 694514 151746 694516
rect 151854 694514 151860 694516
rect 151740 694454 151860 694514
rect 151740 694452 151746 694454
rect 151854 694452 151860 694454
rect 151924 694452 151930 694516
rect 166942 694452 166948 694516
rect 167012 694514 167018 694516
rect 176878 694514 176884 694516
rect 167012 694454 176884 694514
rect 167012 694452 167018 694454
rect 176878 694452 176884 694454
rect 176948 694452 176954 694516
rect 177070 694514 177130 694590
rect 186262 694588 186268 694652
rect 186332 694650 186338 694652
rect 215334 694650 215340 694652
rect 186332 694590 215340 694650
rect 186332 694588 186338 694590
rect 215334 694588 215340 694590
rect 215404 694588 215410 694652
rect 224350 694588 224356 694652
rect 224420 694650 224426 694652
rect 231902 694650 231962 694726
rect 236678 694724 236684 694726
rect 236748 694724 236754 694788
rect 241094 694724 241100 694788
rect 241164 694786 241170 694788
rect 246062 694786 246068 694788
rect 241164 694726 246068 694786
rect 241164 694724 241170 694726
rect 246062 694724 246068 694726
rect 246132 694724 246138 694788
rect 255998 694786 256004 694788
rect 251222 694726 256004 694786
rect 224420 694590 231962 694650
rect 224420 694588 224426 694590
rect 243854 694588 243860 694652
rect 243924 694650 243930 694652
rect 251222 694650 251282 694726
rect 255998 694724 256004 694726
rect 256068 694724 256074 694788
rect 264278 694724 264284 694788
rect 264348 694786 264354 694788
rect 270350 694786 270356 694788
rect 264348 694726 270356 694786
rect 264348 694724 264354 694726
rect 270350 694724 270356 694726
rect 270420 694724 270426 694788
rect 318742 694724 318748 694788
rect 318812 694786 318818 694788
rect 328310 694786 328316 694788
rect 318812 694726 328316 694786
rect 318812 694724 318818 694726
rect 328310 694724 328316 694726
rect 328380 694724 328386 694788
rect 350574 694724 350580 694788
rect 350644 694786 350650 694788
rect 357382 694786 357388 694788
rect 350644 694726 357388 694786
rect 350644 694724 350650 694726
rect 357382 694724 357388 694726
rect 357452 694724 357458 694788
rect 434662 694786 434668 694788
rect 424918 694726 434668 694786
rect 243924 694590 251282 694650
rect 243924 694588 243930 694590
rect 263174 694588 263180 694652
rect 263244 694650 263250 694652
rect 273110 694650 273116 694652
rect 263244 694590 273116 694650
rect 263244 694588 263250 694590
rect 273110 694588 273116 694590
rect 273180 694588 273186 694652
rect 282678 694588 282684 694652
rect 282748 694650 282754 694652
rect 311934 694650 311940 694652
rect 282748 694590 311940 694650
rect 282748 694588 282754 694590
rect 311934 694588 311940 694590
rect 312004 694588 312010 694652
rect 320950 694588 320956 694652
rect 321020 694650 321026 694652
rect 332910 694650 332916 694652
rect 321020 694590 332916 694650
rect 321020 694588 321026 694590
rect 332910 694588 332916 694590
rect 332980 694588 332986 694652
rect 338614 694650 338620 694652
rect 338070 694590 338620 694650
rect 177070 694454 186882 694514
rect 120950 694318 130578 694378
rect 106222 694106 106228 694108
rect 98686 694046 106228 694106
rect 106222 694044 106228 694046
rect 106292 694044 106298 694108
rect 120574 694044 120580 694108
rect 120644 694106 120650 694108
rect 130326 694106 130332 694108
rect 120644 694046 130332 694106
rect 120644 694044 120650 694046
rect 130326 694044 130332 694046
rect 130396 694044 130402 694108
rect 130518 694106 130578 694318
rect 141918 694316 141924 694380
rect 141988 694378 141994 694380
rect 142102 694378 142108 694380
rect 141988 694318 142108 694378
rect 141988 694316 141994 694318
rect 142102 694316 142108 694318
rect 142172 694316 142178 694380
rect 146886 694316 146892 694380
rect 146956 694378 146962 694380
rect 152774 694378 152780 694380
rect 146956 694318 152780 694378
rect 146956 694316 146962 694318
rect 152774 694316 152780 694318
rect 152844 694316 152850 694380
rect 164182 694378 164188 694380
rect 153150 694318 164188 694378
rect 137318 694106 137324 694108
rect 130518 694046 137324 694106
rect 137318 694044 137324 694046
rect 137388 694044 137394 694108
rect 138238 694044 138244 694108
rect 138308 694106 138314 694108
rect 146886 694106 146892 694108
rect 138308 694046 146892 694106
rect 138308 694044 138314 694046
rect 146886 694044 146892 694046
rect 146956 694044 146962 694108
rect 152038 694044 152044 694108
rect 152108 694106 152114 694108
rect 153150 694106 153210 694318
rect 164182 694316 164188 694318
rect 164252 694316 164258 694380
rect 179638 694316 179644 694380
rect 179708 694378 179714 694380
rect 186078 694378 186084 694380
rect 179708 694318 186084 694378
rect 179708 694316 179714 694318
rect 186078 694316 186084 694318
rect 186148 694316 186154 694380
rect 186822 694378 186882 694454
rect 202638 694452 202644 694516
rect 202708 694514 202714 694516
rect 202708 694454 212458 694514
rect 202708 694452 202714 694454
rect 196198 694378 196204 694380
rect 186822 694318 196204 694378
rect 196198 694316 196204 694318
rect 196268 694316 196274 694380
rect 212398 694378 212458 694454
rect 214966 694452 214972 694516
rect 215036 694514 215042 694516
rect 215518 694514 215524 694516
rect 215036 694454 215524 694514
rect 215036 694452 215042 694454
rect 215518 694452 215524 694454
rect 215588 694452 215594 694516
rect 265566 694514 265572 694516
rect 260422 694454 265572 694514
rect 222142 694378 222148 694380
rect 212398 694318 222148 694378
rect 222142 694316 222148 694318
rect 222212 694316 222218 694380
rect 226926 694316 226932 694380
rect 226996 694378 227002 694380
rect 226996 694318 231778 694378
rect 226996 694316 227002 694318
rect 173750 694180 173756 694244
rect 173820 694242 173826 694244
rect 176694 694242 176700 694244
rect 173820 694182 176700 694242
rect 173820 694180 173826 694182
rect 176694 694180 176700 694182
rect 176764 694180 176770 694244
rect 215702 694180 215708 694244
rect 215772 694242 215778 694244
rect 231718 694242 231778 694318
rect 231894 694316 231900 694380
rect 231964 694316 231970 694380
rect 232078 694316 232084 694380
rect 232148 694378 232154 694380
rect 235942 694378 235948 694380
rect 232148 694318 235948 694378
rect 232148 694316 232154 694318
rect 235942 694316 235948 694318
rect 236012 694316 236018 694380
rect 241094 694378 241100 694380
rect 236502 694318 241100 694378
rect 231902 694242 231962 694316
rect 215772 694182 224602 694242
rect 231718 694182 231962 694242
rect 215772 694180 215778 694182
rect 152108 694046 153210 694106
rect 152108 694044 152114 694046
rect 159398 694044 159404 694108
rect 159468 694106 159474 694108
rect 166942 694106 166948 694108
rect 159468 694046 166948 694106
rect 159468 694044 159474 694046
rect 166942 694044 166948 694046
rect 167012 694044 167018 694108
rect 176878 694044 176884 694108
rect 176948 694106 176954 694108
rect 185894 694106 185900 694108
rect 176948 694046 185900 694106
rect 176948 694044 176954 694046
rect 185894 694044 185900 694046
rect 185964 694044 185970 694108
rect 186078 694044 186084 694108
rect 186148 694106 186154 694108
rect 186262 694106 186268 694108
rect 186148 694046 186268 694106
rect 186148 694044 186154 694046
rect 186262 694044 186268 694046
rect 186332 694044 186338 694108
rect 186446 694044 186452 694108
rect 186516 694106 186522 694108
rect 205398 694106 205404 694108
rect 186516 694046 205404 694106
rect 186516 694044 186522 694046
rect 205398 694044 205404 694046
rect 205468 694044 205474 694108
rect 205950 694044 205956 694108
rect 206020 694106 206026 694108
rect 214966 694106 214972 694108
rect 206020 694046 214972 694106
rect 206020 694044 206026 694046
rect 214966 694044 214972 694046
rect 215036 694044 215042 694108
rect 215334 694044 215340 694108
rect 215404 694106 215410 694108
rect 224350 694106 224356 694108
rect 215404 694046 224356 694106
rect 215404 694044 215410 694046
rect 224350 694044 224356 694046
rect 224420 694044 224426 694108
rect 224542 694106 224602 694182
rect 236502 694106 236562 694318
rect 241094 694316 241100 694318
rect 241164 694316 241170 694380
rect 246062 694316 246068 694380
rect 246132 694316 246138 694380
rect 251214 694316 251220 694380
rect 251284 694316 251290 694380
rect 251398 694316 251404 694380
rect 251468 694378 251474 694380
rect 255262 694378 255268 694380
rect 251468 694318 255268 694378
rect 251468 694316 251474 694318
rect 255262 694316 255268 694318
rect 255332 694316 255338 694380
rect 260422 694378 260482 694454
rect 265566 694452 265572 694454
rect 265636 694452 265642 694516
rect 299238 694452 299244 694516
rect 299308 694514 299314 694516
rect 299308 694454 309058 694514
rect 299308 694452 299314 694454
rect 255822 694318 260482 694378
rect 236862 694180 236868 694244
rect 236932 694242 236938 694244
rect 245694 694242 245700 694244
rect 236932 694182 245700 694242
rect 236932 694180 236938 694182
rect 245694 694180 245700 694182
rect 245764 694180 245770 694244
rect 224542 694046 236562 694106
rect 236678 694044 236684 694108
rect 236748 694106 236754 694108
rect 243854 694106 243860 694108
rect 236748 694046 243860 694106
rect 236748 694044 236754 694046
rect 243854 694044 243860 694046
rect 243924 694044 243930 694108
rect 246070 694106 246130 694316
rect 246430 694180 246436 694244
rect 246500 694242 246506 694244
rect 251222 694242 251282 694316
rect 246500 694182 251282 694242
rect 246500 694180 246506 694182
rect 255822 694106 255882 694318
rect 270718 694316 270724 694380
rect 270788 694378 270794 694380
rect 283046 694378 283052 694380
rect 270788 694318 283052 694378
rect 270788 694316 270794 694318
rect 283046 694316 283052 694318
rect 283116 694316 283122 694380
rect 283230 694316 283236 694380
rect 283300 694378 283306 694380
rect 292798 694378 292804 694380
rect 283300 694318 292804 694378
rect 283300 694316 283306 694318
rect 292798 694316 292804 694318
rect 292868 694316 292874 694380
rect 308998 694378 309058 694454
rect 311566 694452 311572 694516
rect 311636 694514 311642 694516
rect 312118 694514 312124 694516
rect 311636 694454 312124 694514
rect 311636 694452 311642 694454
rect 312118 694452 312124 694454
rect 312188 694452 312194 694516
rect 333094 694514 333100 694516
rect 328502 694454 333100 694514
rect 318742 694378 318748 694380
rect 308998 694318 318748 694378
rect 318742 694316 318748 694318
rect 318812 694316 318818 694380
rect 328310 694316 328316 694380
rect 328380 694316 328386 694380
rect 256182 694180 256188 694244
rect 256252 694242 256258 694244
rect 264278 694242 264284 694244
rect 256252 694182 264284 694242
rect 256252 694180 256258 694182
rect 264278 694180 264284 694182
rect 264348 694180 264354 694244
rect 270350 694180 270356 694244
rect 270420 694242 270426 694244
rect 270420 694182 275386 694242
rect 270420 694180 270426 694182
rect 246070 694046 255882 694106
rect 255998 694044 256004 694108
rect 256068 694106 256074 694108
rect 263174 694106 263180 694108
rect 256068 694046 263180 694106
rect 256068 694044 256074 694046
rect 263174 694044 263180 694046
rect 263244 694044 263250 694108
rect 265566 694044 265572 694108
rect 265636 694106 265642 694108
rect 270534 694106 270540 694108
rect 265636 694046 270540 694106
rect 265636 694044 265642 694046
rect 270534 694044 270540 694046
rect 270604 694044 270610 694108
rect 275326 694106 275386 694182
rect 278814 694180 278820 694244
rect 278884 694242 278890 694244
rect 282678 694242 282684 694244
rect 278884 694182 282684 694242
rect 278884 694180 278890 694182
rect 282678 694180 282684 694182
rect 282748 694180 282754 694244
rect 312302 694180 312308 694244
rect 312372 694242 312378 694244
rect 328318 694242 328378 694316
rect 328502 694242 328562 694454
rect 333094 694452 333100 694454
rect 333164 694452 333170 694516
rect 338070 694378 338130 694590
rect 338614 694588 338620 694590
rect 338684 694588 338690 694652
rect 340454 694588 340460 694652
rect 340524 694650 340530 694652
rect 346342 694650 346348 694652
rect 340524 694590 346348 694650
rect 340524 694588 340530 694590
rect 346342 694588 346348 694590
rect 346412 694588 346418 694652
rect 359958 694588 359964 694652
rect 360028 694650 360034 694652
rect 424918 694650 424978 694726
rect 434662 694724 434668 694726
rect 434732 694724 434738 694788
rect 360028 694590 424978 694650
rect 360028 694588 360034 694590
rect 492806 694588 492812 694652
rect 492876 694650 492882 694652
rect 500902 694650 500908 694652
rect 492876 694590 500908 694650
rect 492876 694588 492882 694590
rect 500902 694588 500908 694590
rect 500972 694588 500978 694652
rect 531262 694588 531268 694652
rect 531332 694650 531338 694652
rect 531332 694590 540898 694650
rect 531332 694588 531338 694590
rect 341558 694514 341564 694516
rect 312372 694182 321202 694242
rect 328318 694182 328562 694242
rect 332734 694318 338130 694378
rect 338254 694454 341564 694514
rect 312372 694180 312378 694182
rect 279918 694106 279924 694108
rect 270726 694046 271338 694106
rect 275326 694046 279924 694106
rect 270726 693972 270786 694046
rect 86902 693970 86908 693972
rect 86726 693910 86908 693970
rect 86902 693908 86908 693910
rect 86972 693908 86978 693972
rect 87086 693908 87092 693972
rect 87156 693970 87162 693972
rect 270534 693970 270540 693972
rect 87156 693910 270540 693970
rect 87156 693908 87162 693910
rect 270534 693908 270540 693910
rect 270604 693908 270610 693972
rect 270718 693908 270724 693972
rect 270788 693908 270794 693972
rect 271278 693970 271338 694046
rect 279918 694044 279924 694046
rect 279988 694044 279994 694108
rect 283230 694044 283236 694108
rect 283300 694106 283306 694108
rect 301998 694106 302004 694108
rect 283300 694046 302004 694106
rect 283300 694044 283306 694046
rect 301998 694044 302004 694046
rect 302068 694044 302074 694108
rect 302550 694044 302556 694108
rect 302620 694106 302626 694108
rect 311566 694106 311572 694108
rect 302620 694046 311572 694106
rect 302620 694044 302626 694046
rect 311566 694044 311572 694046
rect 311636 694044 311642 694108
rect 311934 694044 311940 694108
rect 312004 694106 312010 694108
rect 320950 694106 320956 694108
rect 312004 694046 320956 694106
rect 312004 694044 312010 694046
rect 320950 694044 320956 694046
rect 321020 694044 321026 694108
rect 321142 694106 321202 694182
rect 332734 694106 332794 694318
rect 333094 694180 333100 694244
rect 333164 694242 333170 694244
rect 338254 694242 338314 694454
rect 341558 694452 341564 694454
rect 341628 694452 341634 694516
rect 376518 694452 376524 694516
rect 376588 694514 376594 694516
rect 376588 694454 380082 694514
rect 376588 694452 376594 694454
rect 338614 694316 338620 694380
rect 338684 694378 338690 694380
rect 338684 694318 340706 694378
rect 338684 694316 338690 694318
rect 333164 694182 338314 694242
rect 333164 694180 333170 694182
rect 321142 694046 332794 694106
rect 332910 694044 332916 694108
rect 332980 694106 332986 694108
rect 340454 694106 340460 694108
rect 332980 694046 340460 694106
rect 332980 694044 332986 694046
rect 340454 694044 340460 694046
rect 340524 694044 340530 694108
rect 340646 694106 340706 694318
rect 350390 694316 350396 694380
rect 350460 694378 350466 694380
rect 350758 694378 350764 694380
rect 350460 694318 350764 694378
rect 350460 694316 350466 694318
rect 350758 694316 350764 694318
rect 350828 694316 350834 694380
rect 351126 694316 351132 694380
rect 351196 694378 351202 694380
rect 351196 694318 361866 694378
rect 351196 694316 351202 694318
rect 341558 694180 341564 694244
rect 341628 694242 341634 694244
rect 350574 694242 350580 694244
rect 341628 694182 350580 694242
rect 341628 694180 341634 694182
rect 350574 694180 350580 694182
rect 350644 694180 350650 694244
rect 351310 694180 351316 694244
rect 351380 694242 351386 694244
rect 359958 694242 359964 694244
rect 351380 694182 359964 694242
rect 351380 694180 351386 694182
rect 359958 694180 359964 694182
rect 360028 694180 360034 694244
rect 350390 694106 350396 694108
rect 340646 694046 350396 694106
rect 350390 694044 350396 694046
rect 350460 694044 350466 694108
rect 361806 694106 361866 694318
rect 362166 694316 362172 694380
rect 362236 694378 362242 694380
rect 370078 694378 370084 694380
rect 362236 694318 370084 694378
rect 362236 694316 362242 694318
rect 370078 694316 370084 694318
rect 370148 694316 370154 694380
rect 380022 694378 380082 694454
rect 395838 694452 395844 694516
rect 395908 694514 395914 694516
rect 395908 694454 405658 694514
rect 395908 694452 395914 694454
rect 389398 694378 389404 694380
rect 380022 694318 389404 694378
rect 389398 694316 389404 694318
rect 389468 694316 389474 694380
rect 405598 694378 405658 694454
rect 427670 694452 427676 694516
rect 427740 694514 427746 694516
rect 427854 694514 427860 694516
rect 427740 694454 427860 694514
rect 427740 694452 427746 694454
rect 427854 694452 427860 694454
rect 427924 694452 427930 694516
rect 437238 694452 437244 694516
rect 437308 694514 437314 694516
rect 437422 694514 437428 694516
rect 437308 694454 437428 694514
rect 437308 694452 437314 694454
rect 437422 694452 437428 694454
rect 437492 694452 437498 694516
rect 446990 694452 446996 694516
rect 447060 694514 447066 694516
rect 447174 694514 447180 694516
rect 447060 694454 447180 694514
rect 447060 694452 447066 694454
rect 447174 694452 447180 694454
rect 447244 694452 447250 694516
rect 476062 694452 476068 694516
rect 476132 694514 476138 694516
rect 521694 694514 521700 694516
rect 476132 694454 490666 694514
rect 476132 694452 476138 694454
rect 417550 694378 417556 694380
rect 405598 694318 417556 694378
rect 417550 694316 417556 694318
rect 417620 694316 417626 694380
rect 417734 694316 417740 694380
rect 417804 694378 417810 694380
rect 417804 694318 418354 694378
rect 417804 694316 417810 694318
rect 410558 694180 410564 694244
rect 410628 694242 410634 694244
rect 414974 694242 414980 694244
rect 410628 694182 414980 694242
rect 410628 694180 410634 694182
rect 414974 694180 414980 694182
rect 415044 694180 415050 694244
rect 418294 694242 418354 694318
rect 418470 694316 418476 694380
rect 418540 694378 418546 694380
rect 418540 694318 432706 694378
rect 418540 694316 418546 694318
rect 432646 694242 432706 694318
rect 437430 694318 437858 694378
rect 437430 694242 437490 694318
rect 418294 694182 418538 694242
rect 432646 694182 437490 694242
rect 437798 694242 437858 694318
rect 439446 694316 439452 694380
rect 439516 694378 439522 694380
rect 451222 694378 451228 694380
rect 439516 694318 451228 694378
rect 439516 694316 439522 694318
rect 451222 694316 451228 694318
rect 451292 694316 451298 694380
rect 475878 694316 475884 694380
rect 475948 694378 475954 694380
rect 475948 694318 476498 694378
rect 475948 694316 475954 694318
rect 476062 694242 476068 694244
rect 437798 694182 476068 694242
rect 379278 694106 379284 694108
rect 361806 694046 379284 694106
rect 379278 694044 379284 694046
rect 379348 694044 379354 694108
rect 379830 694044 379836 694108
rect 379900 694106 379906 694108
rect 398598 694106 398604 694108
rect 379900 694046 398604 694106
rect 379900 694044 379906 694046
rect 398598 694044 398604 694046
rect 398668 694044 398674 694108
rect 399150 694044 399156 694108
rect 399220 694106 399226 694108
rect 417734 694106 417740 694108
rect 399220 694046 417740 694106
rect 399220 694044 399226 694046
rect 417734 694044 417740 694046
rect 417804 694044 417810 694108
rect 418478 694106 418538 694182
rect 476062 694180 476068 694182
rect 476132 694180 476138 694244
rect 427670 694106 427676 694108
rect 418478 694046 427676 694106
rect 427670 694044 427676 694046
rect 427740 694044 427746 694108
rect 427854 694044 427860 694108
rect 427924 694106 427930 694108
rect 437238 694106 437244 694108
rect 427924 694046 437244 694106
rect 427924 694044 427930 694046
rect 437238 694044 437244 694046
rect 437308 694044 437314 694108
rect 437422 694044 437428 694108
rect 437492 694106 437498 694108
rect 446990 694106 446996 694108
rect 437492 694046 446996 694106
rect 437492 694044 437498 694046
rect 446990 694044 446996 694046
rect 447060 694044 447066 694108
rect 451406 694044 451412 694108
rect 451476 694106 451482 694108
rect 475878 694106 475884 694108
rect 451476 694046 475884 694106
rect 451476 694044 451482 694046
rect 475878 694044 475884 694046
rect 475948 694044 475954 694108
rect 476438 694106 476498 694318
rect 490606 694242 490666 694454
rect 512134 694454 521700 694514
rect 505686 694316 505692 694380
rect 505756 694378 505762 694380
rect 512134 694378 512194 694454
rect 521694 694452 521700 694454
rect 521764 694452 521770 694516
rect 505756 694318 510538 694378
rect 505756 694316 505762 694318
rect 492622 694242 492628 694244
rect 490606 694182 492628 694242
rect 492622 694180 492628 694182
rect 492692 694180 492698 694244
rect 510478 694242 510538 694318
rect 511950 694318 512194 694378
rect 540838 694378 540898 694590
rect 543590 694378 543596 694380
rect 540838 694318 543596 694378
rect 511950 694242 512010 694318
rect 543590 694316 543596 694318
rect 543660 694316 543666 694380
rect 562910 694378 562916 694380
rect 555374 694318 562916 694378
rect 510478 694182 512010 694242
rect 521694 694180 521700 694244
rect 521764 694242 521770 694244
rect 531262 694242 531268 694244
rect 521764 694182 531268 694242
rect 521764 694180 521770 694182
rect 531262 694180 531268 694182
rect 531332 694180 531338 694244
rect 543774 694180 543780 694244
rect 543844 694242 543850 694244
rect 555374 694242 555434 694318
rect 562910 694316 562916 694318
rect 562980 694316 562986 694380
rect 568614 694316 568620 694380
rect 568684 694378 568690 694380
rect 568684 694344 572546 694378
rect 568684 694318 572730 694344
rect 568684 694316 568690 694318
rect 572486 694284 572730 694318
rect 543844 694182 555434 694242
rect 543844 694180 543850 694182
rect 563094 694180 563100 694244
rect 563164 694242 563170 694244
rect 568614 694242 568620 694244
rect 563164 694182 568620 694242
rect 563164 694180 563170 694182
rect 568614 694180 568620 694182
rect 568684 694180 568690 694244
rect 572670 694242 572730 694284
rect 574829 694242 574895 694245
rect 572670 694240 574895 694242
rect 572670 694184 574834 694240
rect 574890 694184 574895 694240
rect 572670 694182 574895 694184
rect 574829 694179 574895 694182
rect 529238 694106 529244 694108
rect 476438 694046 529244 694106
rect 529238 694044 529244 694046
rect 529308 694044 529314 694108
rect 538806 694044 538812 694108
rect 538876 694106 538882 694108
rect 548558 694106 548564 694108
rect 538876 694046 548564 694106
rect 538876 694044 538882 694046
rect 548558 694044 548564 694046
rect 548628 694044 548634 694108
rect 569861 694106 569927 694109
rect 579337 694106 579403 694109
rect 569861 694104 579403 694106
rect 569861 694048 569866 694104
rect 569922 694048 579342 694104
rect 579398 694048 579403 694104
rect 569861 694046 579403 694048
rect 569861 694043 569927 694046
rect 579337 694043 579403 694046
rect 410558 693970 410564 693972
rect 271278 693910 410564 693970
rect 410558 693908 410564 693910
rect 410628 693908 410634 693972
rect 410750 693910 415042 693970
rect 29126 693772 29132 693836
rect 29196 693834 29202 693836
rect 37222 693834 37228 693836
rect 29196 693774 37228 693834
rect 29196 693772 29202 693774
rect 37222 693772 37228 693774
rect 37292 693772 37298 693836
rect 71814 693772 71820 693836
rect 71884 693834 71890 693836
rect 231894 693834 231900 693836
rect 71884 693774 231900 693834
rect 71884 693772 71890 693774
rect 231894 693772 231900 693774
rect 231964 693772 231970 693836
rect 232630 693772 232636 693836
rect 232700 693834 232706 693836
rect 251214 693834 251220 693836
rect 232700 693774 251220 693834
rect 232700 693772 232706 693774
rect 251214 693772 251220 693774
rect 251284 693772 251290 693836
rect 251950 693772 251956 693836
rect 252020 693834 252026 693836
rect 410750 693834 410810 693910
rect 252020 693774 410810 693834
rect 414982 693834 415042 693910
rect 415158 693908 415164 693972
rect 415228 693970 415234 693972
rect 580533 693970 580599 693973
rect 415228 693968 580599 693970
rect 415228 693912 580538 693968
rect 580594 693912 580599 693968
rect 415228 693910 580599 693912
rect 415228 693908 415234 693910
rect 580533 693907 580599 693910
rect 580349 693834 580415 693837
rect 414982 693832 580415 693834
rect 414982 693776 580354 693832
rect 580410 693776 580415 693832
rect 414982 693774 580415 693776
rect 252020 693772 252026 693774
rect 580349 693771 580415 693774
rect 7649 693698 7715 693701
rect 102726 693698 102732 693700
rect 7649 693696 102732 693698
rect 7649 693640 7654 693696
rect 7710 693640 102732 693696
rect 7649 693638 102732 693640
rect 7649 693635 7715 693638
rect 102726 693636 102732 693638
rect 102796 693636 102802 693700
rect 103278 693636 103284 693700
rect 103348 693698 103354 693700
rect 232078 693698 232084 693700
rect 103348 693638 232084 693698
rect 103348 693636 103354 693638
rect 232078 693636 232084 693638
rect 232148 693636 232154 693700
rect 235942 693636 235948 693700
rect 236012 693698 236018 693700
rect 251398 693698 251404 693700
rect 236012 693638 251404 693698
rect 236012 693636 236018 693638
rect 251398 693636 251404 693638
rect 251468 693636 251474 693700
rect 255262 693636 255268 693700
rect 255332 693698 255338 693700
rect 270902 693698 270908 693700
rect 255332 693638 270908 693698
rect 255332 693636 255338 693638
rect 270902 693636 270908 693638
rect 270972 693636 270978 693700
rect 271270 693636 271276 693700
rect 271340 693698 271346 693700
rect 414422 693698 414428 693700
rect 271340 693638 414428 693698
rect 271340 693636 271346 693638
rect 414422 693636 414428 693638
rect 414492 693636 414498 693700
rect 415158 693636 415164 693700
rect 415228 693698 415234 693700
rect 521326 693698 521332 693700
rect 415228 693638 521332 693698
rect 415228 693636 415234 693638
rect 521326 693636 521332 693638
rect 521396 693636 521402 693700
rect 529238 693636 529244 693700
rect 529308 693698 529314 693700
rect 538806 693698 538812 693700
rect 529308 693638 538812 693698
rect 529308 693636 529314 693638
rect 538806 693636 538812 693638
rect 538876 693636 538882 693700
rect 548558 693636 548564 693700
rect 548628 693698 548634 693700
rect 569861 693698 569927 693701
rect 548628 693696 569927 693698
rect 548628 693640 569866 693696
rect 569922 693640 569927 693696
rect 548628 693638 569927 693640
rect 548628 693636 548634 693638
rect 569861 693635 569927 693638
rect 580901 686354 580967 686357
rect 583520 686354 584960 686444
rect 580901 686352 584960 686354
rect 580901 686296 580906 686352
rect 580962 686296 584960 686352
rect 580901 686294 584960 686296
rect 580901 686291 580967 686294
rect 583520 686204 584960 686294
rect -960 682274 480 682364
rect 2865 682274 2931 682277
rect -960 682272 2931 682274
rect -960 682216 2870 682272
rect 2926 682216 2931 682272
rect -960 682214 2931 682216
rect -960 682124 480 682214
rect 2865 682211 2931 682214
rect 574553 674930 574619 674933
rect 575473 674930 575539 674933
rect 574553 674928 575539 674930
rect 574553 674872 574558 674928
rect 574614 674872 575478 674928
rect 575534 674872 575539 674928
rect 574553 674870 575539 674872
rect 574553 674867 574619 674870
rect 575473 674867 575539 674870
rect 579797 674658 579863 674661
rect 583520 674658 584960 674748
rect 579797 674656 584960 674658
rect 579797 674600 579802 674656
rect 579858 674600 584960 674656
rect 579797 674598 584960 674600
rect 579797 674595 579863 674598
rect 583520 674508 584960 674598
rect -960 667994 480 668084
rect 2773 667994 2839 667997
rect -960 667992 2839 667994
rect -960 667936 2778 667992
rect 2834 667936 2839 667992
rect -960 667934 2839 667936
rect -960 667844 480 667934
rect 2773 667931 2839 667934
rect 583520 662676 584960 662916
rect -960 653578 480 653668
rect 3049 653578 3115 653581
rect -960 653576 3115 653578
rect -960 653520 3054 653576
rect 3110 653520 3115 653576
rect -960 653518 3115 653520
rect -960 653428 480 653518
rect 3049 653515 3115 653518
rect 579613 651130 579679 651133
rect 583520 651130 584960 651220
rect 579613 651128 584960 651130
rect 579613 651072 579618 651128
rect 579674 651072 584960 651128
rect 579613 651070 584960 651072
rect 579613 651067 579679 651070
rect 583520 650980 584960 651070
rect 579521 639434 579587 639437
rect 583520 639434 584960 639524
rect 579521 639432 584960 639434
rect 579521 639376 579526 639432
rect 579582 639376 584960 639432
rect 579521 639374 584960 639376
rect 579521 639371 579587 639374
rect 583520 639284 584960 639374
rect -960 639012 480 639252
rect 574645 628010 574711 628013
rect 575473 628010 575539 628013
rect 574645 628008 575539 628010
rect 574645 627952 574650 628008
rect 574706 627952 575478 628008
rect 575534 627952 575539 628008
rect 574645 627950 575539 627952
rect 574645 627947 574711 627950
rect 575473 627947 575539 627950
rect 579797 627738 579863 627741
rect 583520 627738 584960 627828
rect 579797 627736 584960 627738
rect 579797 627680 579802 627736
rect 579858 627680 584960 627736
rect 579797 627678 584960 627680
rect 579797 627675 579863 627678
rect 583520 627588 584960 627678
rect -960 624882 480 624972
rect 2957 624882 3023 624885
rect -960 624880 3023 624882
rect -960 624824 2962 624880
rect 3018 624824 3023 624880
rect -960 624822 3023 624824
rect -960 624732 480 624822
rect 2957 624819 3023 624822
rect 583520 615756 584960 615996
rect -960 610466 480 610556
rect 2773 610466 2839 610469
rect -960 610464 2839 610466
rect -960 610408 2778 610464
rect 2834 610408 2839 610464
rect -960 610406 2839 610408
rect -960 610316 480 610406
rect 2773 610403 2839 610406
rect 579613 604210 579679 604213
rect 583520 604210 584960 604300
rect 579613 604208 584960 604210
rect 579613 604152 579618 604208
rect 579674 604152 584960 604208
rect 579613 604150 584960 604152
rect 579613 604147 579679 604150
rect 583520 604060 584960 604150
rect -960 596050 480 596140
rect 3049 596050 3115 596053
rect -960 596048 3115 596050
rect -960 595992 3054 596048
rect 3110 595992 3115 596048
rect -960 595990 3115 595992
rect -960 595900 480 595990
rect 3049 595987 3115 595990
rect 579429 592514 579495 592517
rect 583520 592514 584960 592604
rect 579429 592512 584960 592514
rect 579429 592456 579434 592512
rect 579490 592456 584960 592512
rect 579429 592454 584960 592456
rect 579429 592451 579495 592454
rect 583520 592364 584960 592454
rect -960 581620 480 581860
rect 580165 580818 580231 580821
rect 583520 580818 584960 580908
rect 580165 580816 584960 580818
rect 580165 580760 580170 580816
rect 580226 580760 584960 580816
rect 580165 580758 584960 580760
rect 580165 580755 580231 580758
rect 583520 580668 584960 580758
rect 583520 568836 584960 569076
rect -960 567354 480 567444
rect 2957 567354 3023 567357
rect -960 567352 3023 567354
rect -960 567296 2962 567352
rect 3018 567296 3023 567352
rect -960 567294 3023 567296
rect -960 567204 480 567294
rect 2957 567291 3023 567294
rect 579613 557290 579679 557293
rect 583520 557290 584960 557380
rect 579613 557288 584960 557290
rect 579613 557232 579618 557288
rect 579674 557232 584960 557288
rect 579613 557230 584960 557232
rect 579613 557227 579679 557230
rect 583520 557140 584960 557230
rect -960 553074 480 553164
rect 3141 553074 3207 553077
rect -960 553072 3207 553074
rect -960 553016 3146 553072
rect 3202 553016 3207 553072
rect -960 553014 3207 553016
rect -960 552924 480 553014
rect 3141 553011 3207 553014
rect 579337 545594 579403 545597
rect 583520 545594 584960 545684
rect 579337 545592 584960 545594
rect 579337 545536 579342 545592
rect 579398 545536 584960 545592
rect 579337 545534 584960 545536
rect 579337 545531 579403 545534
rect 583520 545444 584960 545534
rect -960 538658 480 538748
rect 3233 538658 3299 538661
rect -960 538656 3299 538658
rect -960 538600 3238 538656
rect 3294 538600 3299 538656
rect -960 538598 3299 538600
rect -960 538508 480 538598
rect 3233 538595 3299 538598
rect 579705 533898 579771 533901
rect 583520 533898 584960 533988
rect 579705 533896 584960 533898
rect 579705 533840 579710 533896
rect 579766 533840 584960 533896
rect 579705 533838 584960 533840
rect 579705 533835 579771 533838
rect 583520 533748 584960 533838
rect -960 524092 480 524332
rect 583520 521916 584960 522156
rect 580165 510370 580231 510373
rect 583520 510370 584960 510460
rect 580165 510368 584960 510370
rect 580165 510312 580170 510368
rect 580226 510312 584960 510368
rect 580165 510310 584960 510312
rect 580165 510307 580231 510310
rect 583520 510220 584960 510310
rect -960 509962 480 510052
rect 3049 509962 3115 509965
rect -960 509960 3115 509962
rect -960 509904 3054 509960
rect 3110 509904 3115 509960
rect -960 509902 3115 509904
rect -960 509812 480 509902
rect 3049 509899 3115 509902
rect 580165 498674 580231 498677
rect 583520 498674 584960 498764
rect 580165 498672 584960 498674
rect 580165 498616 580170 498672
rect 580226 498616 584960 498672
rect 580165 498614 584960 498616
rect 580165 498611 580231 498614
rect 583520 498524 584960 498614
rect -960 495546 480 495636
rect 3969 495546 4035 495549
rect -960 495544 4035 495546
rect -960 495488 3974 495544
rect 4030 495488 4035 495544
rect -960 495486 4035 495488
rect -960 495396 480 495486
rect 3969 495483 4035 495486
rect 579981 486842 580047 486845
rect 583520 486842 584960 486932
rect 579981 486840 584960 486842
rect 579981 486784 579986 486840
rect 580042 486784 584960 486840
rect 579981 486782 584960 486784
rect 579981 486779 580047 486782
rect 583520 486692 584960 486782
rect -960 481130 480 481220
rect 3233 481130 3299 481133
rect -960 481128 3299 481130
rect -960 481072 3238 481128
rect 3294 481072 3299 481128
rect -960 481070 3299 481072
rect -960 480980 480 481070
rect 3233 481067 3299 481070
rect 583520 474996 584960 475236
rect -960 466700 480 466940
rect 579613 463450 579679 463453
rect 583520 463450 584960 463540
rect 579613 463448 584960 463450
rect 579613 463392 579618 463448
rect 579674 463392 584960 463448
rect 579613 463390 584960 463392
rect 579613 463387 579679 463390
rect 583520 463300 584960 463390
rect -960 452434 480 452524
rect 3049 452434 3115 452437
rect -960 452432 3115 452434
rect -960 452376 3054 452432
rect 3110 452376 3115 452432
rect -960 452374 3115 452376
rect -960 452284 480 452374
rect 3049 452371 3115 452374
rect 579245 451754 579311 451757
rect 583520 451754 584960 451844
rect 579245 451752 584960 451754
rect 579245 451696 579250 451752
rect 579306 451696 584960 451752
rect 579245 451694 584960 451696
rect 579245 451691 579311 451694
rect 583520 451604 584960 451694
rect 579981 439922 580047 439925
rect 583520 439922 584960 440012
rect 579981 439920 584960 439922
rect 579981 439864 579986 439920
rect 580042 439864 584960 439920
rect 579981 439862 584960 439864
rect 579981 439859 580047 439862
rect 583520 439772 584960 439862
rect -960 438018 480 438108
rect 3325 438018 3391 438021
rect -960 438016 3391 438018
rect -960 437960 3330 438016
rect 3386 437960 3391 438016
rect -960 437958 3391 437960
rect -960 437868 480 437958
rect 3325 437955 3391 437958
rect 583520 428076 584960 428316
rect -960 423738 480 423828
rect 3325 423738 3391 423741
rect -960 423736 3391 423738
rect -960 423680 3330 423736
rect 3386 423680 3391 423736
rect -960 423678 3391 423680
rect -960 423588 480 423678
rect 3325 423675 3391 423678
rect 580165 416530 580231 416533
rect 583520 416530 584960 416620
rect 580165 416528 584960 416530
rect 580165 416472 580170 416528
rect 580226 416472 584960 416528
rect 580165 416470 584960 416472
rect 580165 416467 580231 416470
rect 583520 416380 584960 416470
rect -960 409172 480 409412
rect 579153 404834 579219 404837
rect 583520 404834 584960 404924
rect 579153 404832 584960 404834
rect 579153 404776 579158 404832
rect 579214 404776 584960 404832
rect 579153 404774 584960 404776
rect 579153 404771 579219 404774
rect 583520 404684 584960 404774
rect -960 395042 480 395132
rect 3325 395042 3391 395045
rect -960 395040 3391 395042
rect -960 394984 3330 395040
rect 3386 394984 3391 395040
rect -960 394982 3391 394984
rect -960 394892 480 394982
rect 3325 394979 3391 394982
rect 579061 393002 579127 393005
rect 583520 393002 584960 393092
rect 579061 393000 584960 393002
rect 579061 392944 579066 393000
rect 579122 392944 584960 393000
rect 579061 392942 584960 392944
rect 579061 392939 579127 392942
rect 583520 392852 584960 392942
rect 583520 381156 584960 381396
rect -960 380626 480 380716
rect 4061 380626 4127 380629
rect -960 380624 4127 380626
rect -960 380568 4066 380624
rect 4122 380568 4127 380624
rect -960 380566 4127 380568
rect -960 380476 480 380566
rect 4061 380563 4127 380566
rect 580809 369610 580875 369613
rect 583520 369610 584960 369700
rect 580809 369608 584960 369610
rect 580809 369552 580814 369608
rect 580870 369552 584960 369608
rect 580809 369550 584960 369552
rect 580809 369547 580875 369550
rect 583520 369460 584960 369550
rect -960 366210 480 366300
rect 3325 366210 3391 366213
rect -960 366208 3391 366210
rect -960 366152 3330 366208
rect 3386 366152 3391 366208
rect -960 366150 3391 366152
rect -960 366060 480 366150
rect 3325 366147 3391 366150
rect 580809 357914 580875 357917
rect 583520 357914 584960 358004
rect 580809 357912 584960 357914
rect 580809 357856 580814 357912
rect 580870 357856 584960 357912
rect 580809 357854 584960 357856
rect 580809 357851 580875 357854
rect 583520 357764 584960 357854
rect -960 351780 480 352020
rect 579981 346082 580047 346085
rect 583520 346082 584960 346172
rect 579981 346080 584960 346082
rect 579981 346024 579986 346080
rect 580042 346024 584960 346080
rect 579981 346022 584960 346024
rect 579981 346019 580047 346022
rect 583520 345932 584960 346022
rect -960 337514 480 337604
rect 3325 337514 3391 337517
rect -960 337512 3391 337514
rect -960 337456 3330 337512
rect 3386 337456 3391 337512
rect -960 337454 3391 337456
rect -960 337364 480 337454
rect 3325 337451 3391 337454
rect 583520 334236 584960 334476
rect -960 323098 480 323188
rect 2773 323098 2839 323101
rect -960 323096 2839 323098
rect -960 323040 2778 323096
rect 2834 323040 2839 323096
rect -960 323038 2839 323040
rect -960 322948 480 323038
rect 2773 323035 2839 323038
rect 578969 322690 579035 322693
rect 583520 322690 584960 322780
rect 578969 322688 584960 322690
rect 578969 322632 578974 322688
rect 579030 322632 584960 322688
rect 578969 322630 584960 322632
rect 578969 322627 579035 322630
rect 583520 322540 584960 322630
rect 580809 310858 580875 310861
rect 583520 310858 584960 310948
rect 580809 310856 584960 310858
rect 580809 310800 580814 310856
rect 580870 310800 584960 310856
rect 580809 310798 584960 310800
rect 580809 310795 580875 310798
rect 583520 310708 584960 310798
rect -960 308818 480 308908
rect 3877 308818 3943 308821
rect -960 308816 3943 308818
rect -960 308760 3882 308816
rect 3938 308760 3943 308816
rect -960 308758 3943 308760
rect -960 308668 480 308758
rect 3877 308755 3943 308758
rect 579613 299162 579679 299165
rect 583520 299162 584960 299252
rect 579613 299160 584960 299162
rect 579613 299104 579618 299160
rect 579674 299104 584960 299160
rect 579613 299102 584960 299104
rect 579613 299099 579679 299102
rect 583520 299012 584960 299102
rect -960 294402 480 294492
rect 3325 294402 3391 294405
rect -960 294400 3391 294402
rect -960 294344 3330 294400
rect 3386 294344 3391 294400
rect -960 294342 3391 294344
rect -960 294252 480 294342
rect 3325 294339 3391 294342
rect 583520 287316 584960 287556
rect -960 280122 480 280212
rect 2773 280122 2839 280125
rect -960 280120 2839 280122
rect -960 280064 2778 280120
rect 2834 280064 2839 280120
rect -960 280062 2839 280064
rect -960 279972 480 280062
rect 2773 280059 2839 280062
rect 580717 275770 580783 275773
rect 583520 275770 584960 275860
rect 580717 275768 584960 275770
rect 580717 275712 580722 275768
rect 580778 275712 584960 275768
rect 580717 275710 584960 275712
rect 580717 275707 580783 275710
rect 583520 275620 584960 275710
rect -960 265706 480 265796
rect 3141 265706 3207 265709
rect -960 265704 3207 265706
rect -960 265648 3146 265704
rect 3202 265648 3207 265704
rect -960 265646 3207 265648
rect -960 265556 480 265646
rect 3141 265643 3207 265646
rect 580165 263938 580231 263941
rect 583520 263938 584960 264028
rect 580165 263936 584960 263938
rect 580165 263880 580170 263936
rect 580226 263880 584960 263936
rect 580165 263878 584960 263880
rect 580165 263875 580231 263878
rect 583520 263788 584960 263878
rect 580165 252242 580231 252245
rect 583520 252242 584960 252332
rect 580165 252240 584960 252242
rect 580165 252184 580170 252240
rect 580226 252184 584960 252240
rect 580165 252182 584960 252184
rect 580165 252179 580231 252182
rect 583520 252092 584960 252182
rect -960 251290 480 251380
rect 3233 251290 3299 251293
rect -960 251288 3299 251290
rect -960 251232 3238 251288
rect 3294 251232 3299 251288
rect -960 251230 3299 251232
rect -960 251140 480 251230
rect 3233 251227 3299 251230
rect 583520 240396 584960 240636
rect -960 237010 480 237100
rect 4061 237010 4127 237013
rect -960 237008 4127 237010
rect -960 236952 4066 237008
rect 4122 236952 4127 237008
rect -960 236950 4127 236952
rect -960 236860 480 236950
rect 4061 236947 4127 236950
rect 580625 228850 580691 228853
rect 583520 228850 584960 228940
rect 580625 228848 584960 228850
rect 580625 228792 580630 228848
rect 580686 228792 584960 228848
rect 580625 228790 584960 228792
rect 580625 228787 580691 228790
rect 583520 228700 584960 228790
rect -960 222594 480 222684
rect 3785 222594 3851 222597
rect -960 222592 3851 222594
rect -960 222536 3790 222592
rect 3846 222536 3851 222592
rect -960 222534 3851 222536
rect -960 222444 480 222534
rect 3785 222531 3851 222534
rect 578877 217018 578943 217021
rect 583520 217018 584960 217108
rect 578877 217016 584960 217018
rect 578877 216960 578882 217016
rect 578938 216960 584960 217016
rect 578877 216958 584960 216960
rect 578877 216955 578943 216958
rect 583520 216868 584960 216958
rect -960 208178 480 208268
rect 3141 208178 3207 208181
rect -960 208176 3207 208178
rect -960 208120 3146 208176
rect 3202 208120 3207 208176
rect -960 208118 3207 208120
rect -960 208028 480 208118
rect 3141 208115 3207 208118
rect 580165 205322 580231 205325
rect 583520 205322 584960 205412
rect 580165 205320 584960 205322
rect 580165 205264 580170 205320
rect 580226 205264 584960 205320
rect 580165 205262 584960 205264
rect 580165 205259 580231 205262
rect 583520 205172 584960 205262
rect -960 193898 480 193988
rect 2773 193898 2839 193901
rect -960 193896 2839 193898
rect -960 193840 2778 193896
rect 2834 193840 2839 193896
rect -960 193838 2839 193840
rect -960 193748 480 193838
rect 2773 193835 2839 193838
rect 583520 193476 584960 193716
rect 580165 181930 580231 181933
rect 583520 181930 584960 182020
rect 580165 181928 584960 181930
rect 580165 181872 580170 181928
rect 580226 181872 584960 181928
rect 580165 181870 584960 181872
rect 580165 181867 580231 181870
rect 583520 181780 584960 181870
rect -960 179482 480 179572
rect 3693 179482 3759 179485
rect -960 179480 3759 179482
rect -960 179424 3698 179480
rect 3754 179424 3759 179480
rect -960 179422 3759 179424
rect -960 179332 480 179422
rect 3693 179419 3759 179422
rect 579613 170098 579679 170101
rect 583520 170098 584960 170188
rect 579613 170096 584960 170098
rect 579613 170040 579618 170096
rect 579674 170040 584960 170096
rect 579613 170038 584960 170040
rect 579613 170035 579679 170038
rect 583520 169948 584960 170038
rect -960 165066 480 165156
rect 1117 165066 1183 165069
rect -960 165064 1183 165066
rect -960 165008 1122 165064
rect 1178 165008 1183 165064
rect -960 165006 1183 165008
rect -960 164916 480 165006
rect 1117 165003 1183 165006
rect 580625 158402 580691 158405
rect 583520 158402 584960 158492
rect 580625 158400 584960 158402
rect 580625 158344 580630 158400
rect 580686 158344 584960 158400
rect 580625 158342 584960 158344
rect 580625 158339 580691 158342
rect 583520 158252 584960 158342
rect -960 150786 480 150876
rect 2773 150786 2839 150789
rect -960 150784 2839 150786
rect -960 150728 2778 150784
rect 2834 150728 2839 150784
rect -960 150726 2839 150728
rect -960 150636 480 150726
rect 2773 150723 2839 150726
rect 583520 146556 584960 146796
rect -960 136370 480 136460
rect 3325 136370 3391 136373
rect -960 136368 3391 136370
rect -960 136312 3330 136368
rect 3386 136312 3391 136368
rect -960 136310 3391 136312
rect -960 136220 480 136310
rect 3325 136307 3391 136310
rect 580533 134874 580599 134877
rect 583520 134874 584960 134964
rect 580533 134872 584960 134874
rect 580533 134816 580538 134872
rect 580594 134816 584960 134872
rect 580533 134814 584960 134816
rect 580533 134811 580599 134814
rect 583520 134724 584960 134814
rect 580441 123178 580507 123181
rect 583520 123178 584960 123268
rect 580441 123176 584960 123178
rect 580441 123120 580446 123176
rect 580502 123120 584960 123176
rect 580441 123118 584960 123120
rect 580441 123115 580507 123118
rect 583520 123028 584960 123118
rect -960 122090 480 122180
rect 3325 122090 3391 122093
rect -960 122088 3391 122090
rect -960 122032 3330 122088
rect 3386 122032 3391 122088
rect -960 122030 3391 122032
rect -960 121940 480 122030
rect 3325 122027 3391 122030
rect 579613 111482 579679 111485
rect 583520 111482 584960 111572
rect 579613 111480 584960 111482
rect 579613 111424 579618 111480
rect 579674 111424 584960 111480
rect 579613 111422 584960 111424
rect 579613 111419 579679 111422
rect 583520 111332 584960 111422
rect -960 107674 480 107764
rect 3969 107674 4035 107677
rect -960 107672 4035 107674
rect -960 107616 3974 107672
rect 4030 107616 4035 107672
rect -960 107614 4035 107616
rect -960 107524 480 107614
rect 3969 107611 4035 107614
rect 583520 99636 584960 99876
rect -960 93258 480 93348
rect 3601 93258 3667 93261
rect -960 93256 3667 93258
rect -960 93200 3606 93256
rect 3662 93200 3667 93256
rect -960 93198 3667 93200
rect -960 93108 480 93198
rect 3601 93195 3667 93198
rect 580349 87954 580415 87957
rect 583520 87954 584960 88044
rect 580349 87952 584960 87954
rect 580349 87896 580354 87952
rect 580410 87896 584960 87952
rect 580349 87894 584960 87896
rect 580349 87891 580415 87894
rect 583520 87804 584960 87894
rect -960 78978 480 79068
rect 3049 78978 3115 78981
rect -960 78976 3115 78978
rect -960 78920 3054 78976
rect 3110 78920 3115 78976
rect -960 78918 3115 78920
rect -960 78828 480 78918
rect 3049 78915 3115 78918
rect 580257 76258 580323 76261
rect 583520 76258 584960 76348
rect 580257 76256 584960 76258
rect 580257 76200 580262 76256
rect 580318 76200 584960 76256
rect 580257 76198 584960 76200
rect 580257 76195 580323 76198
rect 583520 76108 584960 76198
rect -960 64562 480 64652
rect 2773 64562 2839 64565
rect -960 64560 2839 64562
rect -960 64504 2778 64560
rect 2834 64504 2839 64560
rect -960 64502 2839 64504
rect -960 64412 480 64502
rect 2773 64499 2839 64502
rect 579797 64562 579863 64565
rect 583520 64562 584960 64652
rect 579797 64560 584960 64562
rect 579797 64504 579802 64560
rect 579858 64504 584960 64560
rect 579797 64502 584960 64504
rect 579797 64499 579863 64502
rect 583520 64412 584960 64502
rect 583520 52716 584960 52956
rect -960 50146 480 50236
rect 3509 50146 3575 50149
rect -960 50144 3575 50146
rect -960 50088 3514 50144
rect 3570 50088 3575 50144
rect -960 50086 3575 50088
rect -960 49996 480 50086
rect 3509 50083 3575 50086
rect 580165 41034 580231 41037
rect 583520 41034 584960 41124
rect 580165 41032 584960 41034
rect 580165 40976 580170 41032
rect 580226 40976 584960 41032
rect 580165 40974 584960 40976
rect 580165 40971 580231 40974
rect 583520 40884 584960 40974
rect -960 35866 480 35956
rect 3509 35866 3575 35869
rect -960 35864 3575 35866
rect -960 35808 3514 35864
rect 3570 35808 3575 35864
rect -960 35806 3575 35808
rect -960 35716 480 35806
rect 3509 35803 3575 35806
rect 580165 29338 580231 29341
rect 583520 29338 584960 29428
rect 580165 29336 584960 29338
rect 580165 29280 580170 29336
rect 580226 29280 584960 29336
rect 580165 29278 584960 29280
rect 580165 29275 580231 29278
rect 583520 29188 584960 29278
rect -960 21450 480 21540
rect 3417 21450 3483 21453
rect -960 21448 3483 21450
rect -960 21392 3422 21448
rect 3478 21392 3483 21448
rect -960 21390 3483 21392
rect -960 21300 480 21390
rect 3417 21387 3483 21390
rect 580165 17642 580231 17645
rect 583520 17642 584960 17732
rect 580165 17640 584960 17642
rect 580165 17584 580170 17640
rect 580226 17584 584960 17640
rect 580165 17582 584960 17584
rect 580165 17579 580231 17582
rect 583520 17492 584960 17582
rect -960 7170 480 7260
rect 3141 7170 3207 7173
rect -960 7168 3207 7170
rect -960 7112 3146 7168
rect 3202 7112 3207 7168
rect -960 7110 3207 7112
rect -960 7020 480 7110
rect 3141 7107 3207 7110
rect 18804 6016 19404 6017
rect 18804 5952 18832 6016
rect 18896 5952 18912 6016
rect 18976 5952 18992 6016
rect 19056 5952 19072 6016
rect 19136 5952 19152 6016
rect 19216 5952 19232 6016
rect 19296 5952 19312 6016
rect 19376 5952 19404 6016
rect 18804 5951 19404 5952
rect 54804 6016 55404 6017
rect 54804 5952 54832 6016
rect 54896 5952 54912 6016
rect 54976 5952 54992 6016
rect 55056 5952 55072 6016
rect 55136 5952 55152 6016
rect 55216 5952 55232 6016
rect 55296 5952 55312 6016
rect 55376 5952 55404 6016
rect 54804 5951 55404 5952
rect 90804 6016 91404 6017
rect 90804 5952 90832 6016
rect 90896 5952 90912 6016
rect 90976 5952 90992 6016
rect 91056 5952 91072 6016
rect 91136 5952 91152 6016
rect 91216 5952 91232 6016
rect 91296 5952 91312 6016
rect 91376 5952 91404 6016
rect 90804 5951 91404 5952
rect 126804 6016 127404 6017
rect 126804 5952 126832 6016
rect 126896 5952 126912 6016
rect 126976 5952 126992 6016
rect 127056 5952 127072 6016
rect 127136 5952 127152 6016
rect 127216 5952 127232 6016
rect 127296 5952 127312 6016
rect 127376 5952 127404 6016
rect 126804 5951 127404 5952
rect 162804 6016 163404 6017
rect 162804 5952 162832 6016
rect 162896 5952 162912 6016
rect 162976 5952 162992 6016
rect 163056 5952 163072 6016
rect 163136 5952 163152 6016
rect 163216 5952 163232 6016
rect 163296 5952 163312 6016
rect 163376 5952 163404 6016
rect 162804 5951 163404 5952
rect 198804 6016 199404 6017
rect 198804 5952 198832 6016
rect 198896 5952 198912 6016
rect 198976 5952 198992 6016
rect 199056 5952 199072 6016
rect 199136 5952 199152 6016
rect 199216 5952 199232 6016
rect 199296 5952 199312 6016
rect 199376 5952 199404 6016
rect 198804 5951 199404 5952
rect 234804 6016 235404 6017
rect 234804 5952 234832 6016
rect 234896 5952 234912 6016
rect 234976 5952 234992 6016
rect 235056 5952 235072 6016
rect 235136 5952 235152 6016
rect 235216 5952 235232 6016
rect 235296 5952 235312 6016
rect 235376 5952 235404 6016
rect 234804 5951 235404 5952
rect 270804 6016 271404 6017
rect 270804 5952 270832 6016
rect 270896 5952 270912 6016
rect 270976 5952 270992 6016
rect 271056 5952 271072 6016
rect 271136 5952 271152 6016
rect 271216 5952 271232 6016
rect 271296 5952 271312 6016
rect 271376 5952 271404 6016
rect 270804 5951 271404 5952
rect 306804 6016 307404 6017
rect 306804 5952 306832 6016
rect 306896 5952 306912 6016
rect 306976 5952 306992 6016
rect 307056 5952 307072 6016
rect 307136 5952 307152 6016
rect 307216 5952 307232 6016
rect 307296 5952 307312 6016
rect 307376 5952 307404 6016
rect 306804 5951 307404 5952
rect 342804 6016 343404 6017
rect 342804 5952 342832 6016
rect 342896 5952 342912 6016
rect 342976 5952 342992 6016
rect 343056 5952 343072 6016
rect 343136 5952 343152 6016
rect 343216 5952 343232 6016
rect 343296 5952 343312 6016
rect 343376 5952 343404 6016
rect 342804 5951 343404 5952
rect 378804 6016 379404 6017
rect 378804 5952 378832 6016
rect 378896 5952 378912 6016
rect 378976 5952 378992 6016
rect 379056 5952 379072 6016
rect 379136 5952 379152 6016
rect 379216 5952 379232 6016
rect 379296 5952 379312 6016
rect 379376 5952 379404 6016
rect 378804 5951 379404 5952
rect 414804 6016 415404 6017
rect 414804 5952 414832 6016
rect 414896 5952 414912 6016
rect 414976 5952 414992 6016
rect 415056 5952 415072 6016
rect 415136 5952 415152 6016
rect 415216 5952 415232 6016
rect 415296 5952 415312 6016
rect 415376 5952 415404 6016
rect 414804 5951 415404 5952
rect 450804 6016 451404 6017
rect 450804 5952 450832 6016
rect 450896 5952 450912 6016
rect 450976 5952 450992 6016
rect 451056 5952 451072 6016
rect 451136 5952 451152 6016
rect 451216 5952 451232 6016
rect 451296 5952 451312 6016
rect 451376 5952 451404 6016
rect 450804 5951 451404 5952
rect 486804 6016 487404 6017
rect 486804 5952 486832 6016
rect 486896 5952 486912 6016
rect 486976 5952 486992 6016
rect 487056 5952 487072 6016
rect 487136 5952 487152 6016
rect 487216 5952 487232 6016
rect 487296 5952 487312 6016
rect 487376 5952 487404 6016
rect 486804 5951 487404 5952
rect 522804 6016 523404 6017
rect 522804 5952 522832 6016
rect 522896 5952 522912 6016
rect 522976 5952 522992 6016
rect 523056 5952 523072 6016
rect 523136 5952 523152 6016
rect 523216 5952 523232 6016
rect 523296 5952 523312 6016
rect 523376 5952 523404 6016
rect 522804 5951 523404 5952
rect 558804 6016 559404 6017
rect 558804 5952 558832 6016
rect 558896 5952 558912 6016
rect 558976 5952 558992 6016
rect 559056 5952 559072 6016
rect 559136 5952 559152 6016
rect 559216 5952 559232 6016
rect 559296 5952 559312 6016
rect 559376 5952 559404 6016
rect 558804 5951 559404 5952
rect 583520 5796 584960 6036
rect 36804 5472 37404 5473
rect 36804 5408 36832 5472
rect 36896 5408 36912 5472
rect 36976 5408 36992 5472
rect 37056 5408 37072 5472
rect 37136 5408 37152 5472
rect 37216 5408 37232 5472
rect 37296 5408 37312 5472
rect 37376 5408 37404 5472
rect 36804 5407 37404 5408
rect 72804 5472 73404 5473
rect 72804 5408 72832 5472
rect 72896 5408 72912 5472
rect 72976 5408 72992 5472
rect 73056 5408 73072 5472
rect 73136 5408 73152 5472
rect 73216 5408 73232 5472
rect 73296 5408 73312 5472
rect 73376 5408 73404 5472
rect 72804 5407 73404 5408
rect 108804 5472 109404 5473
rect 108804 5408 108832 5472
rect 108896 5408 108912 5472
rect 108976 5408 108992 5472
rect 109056 5408 109072 5472
rect 109136 5408 109152 5472
rect 109216 5408 109232 5472
rect 109296 5408 109312 5472
rect 109376 5408 109404 5472
rect 108804 5407 109404 5408
rect 144804 5472 145404 5473
rect 144804 5408 144832 5472
rect 144896 5408 144912 5472
rect 144976 5408 144992 5472
rect 145056 5408 145072 5472
rect 145136 5408 145152 5472
rect 145216 5408 145232 5472
rect 145296 5408 145312 5472
rect 145376 5408 145404 5472
rect 144804 5407 145404 5408
rect 180804 5472 181404 5473
rect 180804 5408 180832 5472
rect 180896 5408 180912 5472
rect 180976 5408 180992 5472
rect 181056 5408 181072 5472
rect 181136 5408 181152 5472
rect 181216 5408 181232 5472
rect 181296 5408 181312 5472
rect 181376 5408 181404 5472
rect 180804 5407 181404 5408
rect 216804 5472 217404 5473
rect 216804 5408 216832 5472
rect 216896 5408 216912 5472
rect 216976 5408 216992 5472
rect 217056 5408 217072 5472
rect 217136 5408 217152 5472
rect 217216 5408 217232 5472
rect 217296 5408 217312 5472
rect 217376 5408 217404 5472
rect 216804 5407 217404 5408
rect 252804 5472 253404 5473
rect 252804 5408 252832 5472
rect 252896 5408 252912 5472
rect 252976 5408 252992 5472
rect 253056 5408 253072 5472
rect 253136 5408 253152 5472
rect 253216 5408 253232 5472
rect 253296 5408 253312 5472
rect 253376 5408 253404 5472
rect 252804 5407 253404 5408
rect 288804 5472 289404 5473
rect 288804 5408 288832 5472
rect 288896 5408 288912 5472
rect 288976 5408 288992 5472
rect 289056 5408 289072 5472
rect 289136 5408 289152 5472
rect 289216 5408 289232 5472
rect 289296 5408 289312 5472
rect 289376 5408 289404 5472
rect 288804 5407 289404 5408
rect 324804 5472 325404 5473
rect 324804 5408 324832 5472
rect 324896 5408 324912 5472
rect 324976 5408 324992 5472
rect 325056 5408 325072 5472
rect 325136 5408 325152 5472
rect 325216 5408 325232 5472
rect 325296 5408 325312 5472
rect 325376 5408 325404 5472
rect 324804 5407 325404 5408
rect 360804 5472 361404 5473
rect 360804 5408 360832 5472
rect 360896 5408 360912 5472
rect 360976 5408 360992 5472
rect 361056 5408 361072 5472
rect 361136 5408 361152 5472
rect 361216 5408 361232 5472
rect 361296 5408 361312 5472
rect 361376 5408 361404 5472
rect 360804 5407 361404 5408
rect 396804 5472 397404 5473
rect 396804 5408 396832 5472
rect 396896 5408 396912 5472
rect 396976 5408 396992 5472
rect 397056 5408 397072 5472
rect 397136 5408 397152 5472
rect 397216 5408 397232 5472
rect 397296 5408 397312 5472
rect 397376 5408 397404 5472
rect 396804 5407 397404 5408
rect 432804 5472 433404 5473
rect 432804 5408 432832 5472
rect 432896 5408 432912 5472
rect 432976 5408 432992 5472
rect 433056 5408 433072 5472
rect 433136 5408 433152 5472
rect 433216 5408 433232 5472
rect 433296 5408 433312 5472
rect 433376 5408 433404 5472
rect 432804 5407 433404 5408
rect 468804 5472 469404 5473
rect 468804 5408 468832 5472
rect 468896 5408 468912 5472
rect 468976 5408 468992 5472
rect 469056 5408 469072 5472
rect 469136 5408 469152 5472
rect 469216 5408 469232 5472
rect 469296 5408 469312 5472
rect 469376 5408 469404 5472
rect 468804 5407 469404 5408
rect 504804 5472 505404 5473
rect 504804 5408 504832 5472
rect 504896 5408 504912 5472
rect 504976 5408 504992 5472
rect 505056 5408 505072 5472
rect 505136 5408 505152 5472
rect 505216 5408 505232 5472
rect 505296 5408 505312 5472
rect 505376 5408 505404 5472
rect 504804 5407 505404 5408
rect 540804 5472 541404 5473
rect 540804 5408 540832 5472
rect 540896 5408 540912 5472
rect 540976 5408 540992 5472
rect 541056 5408 541072 5472
rect 541136 5408 541152 5472
rect 541216 5408 541232 5472
rect 541296 5408 541312 5472
rect 541376 5408 541404 5472
rect 540804 5407 541404 5408
rect 576804 5472 577404 5473
rect 576804 5408 576832 5472
rect 576896 5408 576912 5472
rect 576976 5408 576992 5472
rect 577056 5408 577072 5472
rect 577136 5408 577152 5472
rect 577216 5408 577232 5472
rect 577296 5408 577312 5472
rect 577376 5408 577404 5472
rect 576804 5407 577404 5408
rect 18804 4928 19404 4929
rect 18804 4864 18832 4928
rect 18896 4864 18912 4928
rect 18976 4864 18992 4928
rect 19056 4864 19072 4928
rect 19136 4864 19152 4928
rect 19216 4864 19232 4928
rect 19296 4864 19312 4928
rect 19376 4864 19404 4928
rect 18804 4863 19404 4864
rect 54804 4928 55404 4929
rect 54804 4864 54832 4928
rect 54896 4864 54912 4928
rect 54976 4864 54992 4928
rect 55056 4864 55072 4928
rect 55136 4864 55152 4928
rect 55216 4864 55232 4928
rect 55296 4864 55312 4928
rect 55376 4864 55404 4928
rect 54804 4863 55404 4864
rect 90804 4928 91404 4929
rect 90804 4864 90832 4928
rect 90896 4864 90912 4928
rect 90976 4864 90992 4928
rect 91056 4864 91072 4928
rect 91136 4864 91152 4928
rect 91216 4864 91232 4928
rect 91296 4864 91312 4928
rect 91376 4864 91404 4928
rect 90804 4863 91404 4864
rect 126804 4928 127404 4929
rect 126804 4864 126832 4928
rect 126896 4864 126912 4928
rect 126976 4864 126992 4928
rect 127056 4864 127072 4928
rect 127136 4864 127152 4928
rect 127216 4864 127232 4928
rect 127296 4864 127312 4928
rect 127376 4864 127404 4928
rect 126804 4863 127404 4864
rect 162804 4928 163404 4929
rect 162804 4864 162832 4928
rect 162896 4864 162912 4928
rect 162976 4864 162992 4928
rect 163056 4864 163072 4928
rect 163136 4864 163152 4928
rect 163216 4864 163232 4928
rect 163296 4864 163312 4928
rect 163376 4864 163404 4928
rect 162804 4863 163404 4864
rect 198804 4928 199404 4929
rect 198804 4864 198832 4928
rect 198896 4864 198912 4928
rect 198976 4864 198992 4928
rect 199056 4864 199072 4928
rect 199136 4864 199152 4928
rect 199216 4864 199232 4928
rect 199296 4864 199312 4928
rect 199376 4864 199404 4928
rect 198804 4863 199404 4864
rect 234804 4928 235404 4929
rect 234804 4864 234832 4928
rect 234896 4864 234912 4928
rect 234976 4864 234992 4928
rect 235056 4864 235072 4928
rect 235136 4864 235152 4928
rect 235216 4864 235232 4928
rect 235296 4864 235312 4928
rect 235376 4864 235404 4928
rect 234804 4863 235404 4864
rect 270804 4928 271404 4929
rect 270804 4864 270832 4928
rect 270896 4864 270912 4928
rect 270976 4864 270992 4928
rect 271056 4864 271072 4928
rect 271136 4864 271152 4928
rect 271216 4864 271232 4928
rect 271296 4864 271312 4928
rect 271376 4864 271404 4928
rect 270804 4863 271404 4864
rect 306804 4928 307404 4929
rect 306804 4864 306832 4928
rect 306896 4864 306912 4928
rect 306976 4864 306992 4928
rect 307056 4864 307072 4928
rect 307136 4864 307152 4928
rect 307216 4864 307232 4928
rect 307296 4864 307312 4928
rect 307376 4864 307404 4928
rect 306804 4863 307404 4864
rect 342804 4928 343404 4929
rect 342804 4864 342832 4928
rect 342896 4864 342912 4928
rect 342976 4864 342992 4928
rect 343056 4864 343072 4928
rect 343136 4864 343152 4928
rect 343216 4864 343232 4928
rect 343296 4864 343312 4928
rect 343376 4864 343404 4928
rect 342804 4863 343404 4864
rect 378804 4928 379404 4929
rect 378804 4864 378832 4928
rect 378896 4864 378912 4928
rect 378976 4864 378992 4928
rect 379056 4864 379072 4928
rect 379136 4864 379152 4928
rect 379216 4864 379232 4928
rect 379296 4864 379312 4928
rect 379376 4864 379404 4928
rect 378804 4863 379404 4864
rect 414804 4928 415404 4929
rect 414804 4864 414832 4928
rect 414896 4864 414912 4928
rect 414976 4864 414992 4928
rect 415056 4864 415072 4928
rect 415136 4864 415152 4928
rect 415216 4864 415232 4928
rect 415296 4864 415312 4928
rect 415376 4864 415404 4928
rect 414804 4863 415404 4864
rect 450804 4928 451404 4929
rect 450804 4864 450832 4928
rect 450896 4864 450912 4928
rect 450976 4864 450992 4928
rect 451056 4864 451072 4928
rect 451136 4864 451152 4928
rect 451216 4864 451232 4928
rect 451296 4864 451312 4928
rect 451376 4864 451404 4928
rect 450804 4863 451404 4864
rect 486804 4928 487404 4929
rect 486804 4864 486832 4928
rect 486896 4864 486912 4928
rect 486976 4864 486992 4928
rect 487056 4864 487072 4928
rect 487136 4864 487152 4928
rect 487216 4864 487232 4928
rect 487296 4864 487312 4928
rect 487376 4864 487404 4928
rect 486804 4863 487404 4864
rect 522804 4928 523404 4929
rect 522804 4864 522832 4928
rect 522896 4864 522912 4928
rect 522976 4864 522992 4928
rect 523056 4864 523072 4928
rect 523136 4864 523152 4928
rect 523216 4864 523232 4928
rect 523296 4864 523312 4928
rect 523376 4864 523404 4928
rect 522804 4863 523404 4864
rect 558804 4928 559404 4929
rect 558804 4864 558832 4928
rect 558896 4864 558912 4928
rect 558976 4864 558992 4928
rect 559056 4864 559072 4928
rect 559136 4864 559152 4928
rect 559216 4864 559232 4928
rect 559296 4864 559312 4928
rect 559376 4864 559404 4928
rect 558804 4863 559404 4864
rect 36804 4384 37404 4385
rect 36804 4320 36832 4384
rect 36896 4320 36912 4384
rect 36976 4320 36992 4384
rect 37056 4320 37072 4384
rect 37136 4320 37152 4384
rect 37216 4320 37232 4384
rect 37296 4320 37312 4384
rect 37376 4320 37404 4384
rect 36804 4319 37404 4320
rect 72804 4384 73404 4385
rect 72804 4320 72832 4384
rect 72896 4320 72912 4384
rect 72976 4320 72992 4384
rect 73056 4320 73072 4384
rect 73136 4320 73152 4384
rect 73216 4320 73232 4384
rect 73296 4320 73312 4384
rect 73376 4320 73404 4384
rect 72804 4319 73404 4320
rect 108804 4384 109404 4385
rect 108804 4320 108832 4384
rect 108896 4320 108912 4384
rect 108976 4320 108992 4384
rect 109056 4320 109072 4384
rect 109136 4320 109152 4384
rect 109216 4320 109232 4384
rect 109296 4320 109312 4384
rect 109376 4320 109404 4384
rect 108804 4319 109404 4320
rect 144804 4384 145404 4385
rect 144804 4320 144832 4384
rect 144896 4320 144912 4384
rect 144976 4320 144992 4384
rect 145056 4320 145072 4384
rect 145136 4320 145152 4384
rect 145216 4320 145232 4384
rect 145296 4320 145312 4384
rect 145376 4320 145404 4384
rect 144804 4319 145404 4320
rect 180804 4384 181404 4385
rect 180804 4320 180832 4384
rect 180896 4320 180912 4384
rect 180976 4320 180992 4384
rect 181056 4320 181072 4384
rect 181136 4320 181152 4384
rect 181216 4320 181232 4384
rect 181296 4320 181312 4384
rect 181376 4320 181404 4384
rect 180804 4319 181404 4320
rect 216804 4384 217404 4385
rect 216804 4320 216832 4384
rect 216896 4320 216912 4384
rect 216976 4320 216992 4384
rect 217056 4320 217072 4384
rect 217136 4320 217152 4384
rect 217216 4320 217232 4384
rect 217296 4320 217312 4384
rect 217376 4320 217404 4384
rect 216804 4319 217404 4320
rect 252804 4384 253404 4385
rect 252804 4320 252832 4384
rect 252896 4320 252912 4384
rect 252976 4320 252992 4384
rect 253056 4320 253072 4384
rect 253136 4320 253152 4384
rect 253216 4320 253232 4384
rect 253296 4320 253312 4384
rect 253376 4320 253404 4384
rect 252804 4319 253404 4320
rect 288804 4384 289404 4385
rect 288804 4320 288832 4384
rect 288896 4320 288912 4384
rect 288976 4320 288992 4384
rect 289056 4320 289072 4384
rect 289136 4320 289152 4384
rect 289216 4320 289232 4384
rect 289296 4320 289312 4384
rect 289376 4320 289404 4384
rect 288804 4319 289404 4320
rect 324804 4384 325404 4385
rect 324804 4320 324832 4384
rect 324896 4320 324912 4384
rect 324976 4320 324992 4384
rect 325056 4320 325072 4384
rect 325136 4320 325152 4384
rect 325216 4320 325232 4384
rect 325296 4320 325312 4384
rect 325376 4320 325404 4384
rect 324804 4319 325404 4320
rect 360804 4384 361404 4385
rect 360804 4320 360832 4384
rect 360896 4320 360912 4384
rect 360976 4320 360992 4384
rect 361056 4320 361072 4384
rect 361136 4320 361152 4384
rect 361216 4320 361232 4384
rect 361296 4320 361312 4384
rect 361376 4320 361404 4384
rect 360804 4319 361404 4320
rect 396804 4384 397404 4385
rect 396804 4320 396832 4384
rect 396896 4320 396912 4384
rect 396976 4320 396992 4384
rect 397056 4320 397072 4384
rect 397136 4320 397152 4384
rect 397216 4320 397232 4384
rect 397296 4320 397312 4384
rect 397376 4320 397404 4384
rect 396804 4319 397404 4320
rect 432804 4384 433404 4385
rect 432804 4320 432832 4384
rect 432896 4320 432912 4384
rect 432976 4320 432992 4384
rect 433056 4320 433072 4384
rect 433136 4320 433152 4384
rect 433216 4320 433232 4384
rect 433296 4320 433312 4384
rect 433376 4320 433404 4384
rect 432804 4319 433404 4320
rect 468804 4384 469404 4385
rect 468804 4320 468832 4384
rect 468896 4320 468912 4384
rect 468976 4320 468992 4384
rect 469056 4320 469072 4384
rect 469136 4320 469152 4384
rect 469216 4320 469232 4384
rect 469296 4320 469312 4384
rect 469376 4320 469404 4384
rect 468804 4319 469404 4320
rect 504804 4384 505404 4385
rect 504804 4320 504832 4384
rect 504896 4320 504912 4384
rect 504976 4320 504992 4384
rect 505056 4320 505072 4384
rect 505136 4320 505152 4384
rect 505216 4320 505232 4384
rect 505296 4320 505312 4384
rect 505376 4320 505404 4384
rect 504804 4319 505404 4320
rect 540804 4384 541404 4385
rect 540804 4320 540832 4384
rect 540896 4320 540912 4384
rect 540976 4320 540992 4384
rect 541056 4320 541072 4384
rect 541136 4320 541152 4384
rect 541216 4320 541232 4384
rect 541296 4320 541312 4384
rect 541376 4320 541404 4384
rect 540804 4319 541404 4320
rect 576804 4384 577404 4385
rect 576804 4320 576832 4384
rect 576896 4320 576912 4384
rect 576976 4320 576992 4384
rect 577056 4320 577072 4384
rect 577136 4320 577152 4384
rect 577216 4320 577232 4384
rect 577296 4320 577312 4384
rect 577376 4320 577404 4384
rect 576804 4319 577404 4320
rect 18804 3840 19404 3841
rect 18804 3776 18832 3840
rect 18896 3776 18912 3840
rect 18976 3776 18992 3840
rect 19056 3776 19072 3840
rect 19136 3776 19152 3840
rect 19216 3776 19232 3840
rect 19296 3776 19312 3840
rect 19376 3776 19404 3840
rect 18804 3775 19404 3776
rect 54804 3840 55404 3841
rect 54804 3776 54832 3840
rect 54896 3776 54912 3840
rect 54976 3776 54992 3840
rect 55056 3776 55072 3840
rect 55136 3776 55152 3840
rect 55216 3776 55232 3840
rect 55296 3776 55312 3840
rect 55376 3776 55404 3840
rect 54804 3775 55404 3776
rect 90804 3840 91404 3841
rect 90804 3776 90832 3840
rect 90896 3776 90912 3840
rect 90976 3776 90992 3840
rect 91056 3776 91072 3840
rect 91136 3776 91152 3840
rect 91216 3776 91232 3840
rect 91296 3776 91312 3840
rect 91376 3776 91404 3840
rect 90804 3775 91404 3776
rect 126804 3840 127404 3841
rect 126804 3776 126832 3840
rect 126896 3776 126912 3840
rect 126976 3776 126992 3840
rect 127056 3776 127072 3840
rect 127136 3776 127152 3840
rect 127216 3776 127232 3840
rect 127296 3776 127312 3840
rect 127376 3776 127404 3840
rect 126804 3775 127404 3776
rect 162804 3840 163404 3841
rect 162804 3776 162832 3840
rect 162896 3776 162912 3840
rect 162976 3776 162992 3840
rect 163056 3776 163072 3840
rect 163136 3776 163152 3840
rect 163216 3776 163232 3840
rect 163296 3776 163312 3840
rect 163376 3776 163404 3840
rect 162804 3775 163404 3776
rect 198804 3840 199404 3841
rect 198804 3776 198832 3840
rect 198896 3776 198912 3840
rect 198976 3776 198992 3840
rect 199056 3776 199072 3840
rect 199136 3776 199152 3840
rect 199216 3776 199232 3840
rect 199296 3776 199312 3840
rect 199376 3776 199404 3840
rect 198804 3775 199404 3776
rect 234804 3840 235404 3841
rect 234804 3776 234832 3840
rect 234896 3776 234912 3840
rect 234976 3776 234992 3840
rect 235056 3776 235072 3840
rect 235136 3776 235152 3840
rect 235216 3776 235232 3840
rect 235296 3776 235312 3840
rect 235376 3776 235404 3840
rect 234804 3775 235404 3776
rect 270804 3840 271404 3841
rect 270804 3776 270832 3840
rect 270896 3776 270912 3840
rect 270976 3776 270992 3840
rect 271056 3776 271072 3840
rect 271136 3776 271152 3840
rect 271216 3776 271232 3840
rect 271296 3776 271312 3840
rect 271376 3776 271404 3840
rect 270804 3775 271404 3776
rect 306804 3840 307404 3841
rect 306804 3776 306832 3840
rect 306896 3776 306912 3840
rect 306976 3776 306992 3840
rect 307056 3776 307072 3840
rect 307136 3776 307152 3840
rect 307216 3776 307232 3840
rect 307296 3776 307312 3840
rect 307376 3776 307404 3840
rect 306804 3775 307404 3776
rect 342804 3840 343404 3841
rect 342804 3776 342832 3840
rect 342896 3776 342912 3840
rect 342976 3776 342992 3840
rect 343056 3776 343072 3840
rect 343136 3776 343152 3840
rect 343216 3776 343232 3840
rect 343296 3776 343312 3840
rect 343376 3776 343404 3840
rect 342804 3775 343404 3776
rect 378804 3840 379404 3841
rect 378804 3776 378832 3840
rect 378896 3776 378912 3840
rect 378976 3776 378992 3840
rect 379056 3776 379072 3840
rect 379136 3776 379152 3840
rect 379216 3776 379232 3840
rect 379296 3776 379312 3840
rect 379376 3776 379404 3840
rect 378804 3775 379404 3776
rect 414804 3840 415404 3841
rect 414804 3776 414832 3840
rect 414896 3776 414912 3840
rect 414976 3776 414992 3840
rect 415056 3776 415072 3840
rect 415136 3776 415152 3840
rect 415216 3776 415232 3840
rect 415296 3776 415312 3840
rect 415376 3776 415404 3840
rect 414804 3775 415404 3776
rect 450804 3840 451404 3841
rect 450804 3776 450832 3840
rect 450896 3776 450912 3840
rect 450976 3776 450992 3840
rect 451056 3776 451072 3840
rect 451136 3776 451152 3840
rect 451216 3776 451232 3840
rect 451296 3776 451312 3840
rect 451376 3776 451404 3840
rect 450804 3775 451404 3776
rect 486804 3840 487404 3841
rect 486804 3776 486832 3840
rect 486896 3776 486912 3840
rect 486976 3776 486992 3840
rect 487056 3776 487072 3840
rect 487136 3776 487152 3840
rect 487216 3776 487232 3840
rect 487296 3776 487312 3840
rect 487376 3776 487404 3840
rect 486804 3775 487404 3776
rect 522804 3840 523404 3841
rect 522804 3776 522832 3840
rect 522896 3776 522912 3840
rect 522976 3776 522992 3840
rect 523056 3776 523072 3840
rect 523136 3776 523152 3840
rect 523216 3776 523232 3840
rect 523296 3776 523312 3840
rect 523376 3776 523404 3840
rect 522804 3775 523404 3776
rect 558804 3840 559404 3841
rect 558804 3776 558832 3840
rect 558896 3776 558912 3840
rect 558976 3776 558992 3840
rect 559056 3776 559072 3840
rect 559136 3776 559152 3840
rect 559216 3776 559232 3840
rect 559296 3776 559312 3840
rect 559376 3776 559404 3840
rect 558804 3775 559404 3776
rect 36804 3296 37404 3297
rect 36804 3232 36832 3296
rect 36896 3232 36912 3296
rect 36976 3232 36992 3296
rect 37056 3232 37072 3296
rect 37136 3232 37152 3296
rect 37216 3232 37232 3296
rect 37296 3232 37312 3296
rect 37376 3232 37404 3296
rect 36804 3231 37404 3232
rect 72804 3296 73404 3297
rect 72804 3232 72832 3296
rect 72896 3232 72912 3296
rect 72976 3232 72992 3296
rect 73056 3232 73072 3296
rect 73136 3232 73152 3296
rect 73216 3232 73232 3296
rect 73296 3232 73312 3296
rect 73376 3232 73404 3296
rect 72804 3231 73404 3232
rect 108804 3296 109404 3297
rect 108804 3232 108832 3296
rect 108896 3232 108912 3296
rect 108976 3232 108992 3296
rect 109056 3232 109072 3296
rect 109136 3232 109152 3296
rect 109216 3232 109232 3296
rect 109296 3232 109312 3296
rect 109376 3232 109404 3296
rect 108804 3231 109404 3232
rect 144804 3296 145404 3297
rect 144804 3232 144832 3296
rect 144896 3232 144912 3296
rect 144976 3232 144992 3296
rect 145056 3232 145072 3296
rect 145136 3232 145152 3296
rect 145216 3232 145232 3296
rect 145296 3232 145312 3296
rect 145376 3232 145404 3296
rect 144804 3231 145404 3232
rect 180804 3296 181404 3297
rect 180804 3232 180832 3296
rect 180896 3232 180912 3296
rect 180976 3232 180992 3296
rect 181056 3232 181072 3296
rect 181136 3232 181152 3296
rect 181216 3232 181232 3296
rect 181296 3232 181312 3296
rect 181376 3232 181404 3296
rect 180804 3231 181404 3232
rect 216804 3296 217404 3297
rect 216804 3232 216832 3296
rect 216896 3232 216912 3296
rect 216976 3232 216992 3296
rect 217056 3232 217072 3296
rect 217136 3232 217152 3296
rect 217216 3232 217232 3296
rect 217296 3232 217312 3296
rect 217376 3232 217404 3296
rect 216804 3231 217404 3232
rect 252804 3296 253404 3297
rect 252804 3232 252832 3296
rect 252896 3232 252912 3296
rect 252976 3232 252992 3296
rect 253056 3232 253072 3296
rect 253136 3232 253152 3296
rect 253216 3232 253232 3296
rect 253296 3232 253312 3296
rect 253376 3232 253404 3296
rect 252804 3231 253404 3232
rect 288804 3296 289404 3297
rect 288804 3232 288832 3296
rect 288896 3232 288912 3296
rect 288976 3232 288992 3296
rect 289056 3232 289072 3296
rect 289136 3232 289152 3296
rect 289216 3232 289232 3296
rect 289296 3232 289312 3296
rect 289376 3232 289404 3296
rect 288804 3231 289404 3232
rect 324804 3296 325404 3297
rect 324804 3232 324832 3296
rect 324896 3232 324912 3296
rect 324976 3232 324992 3296
rect 325056 3232 325072 3296
rect 325136 3232 325152 3296
rect 325216 3232 325232 3296
rect 325296 3232 325312 3296
rect 325376 3232 325404 3296
rect 324804 3231 325404 3232
rect 360804 3296 361404 3297
rect 360804 3232 360832 3296
rect 360896 3232 360912 3296
rect 360976 3232 360992 3296
rect 361056 3232 361072 3296
rect 361136 3232 361152 3296
rect 361216 3232 361232 3296
rect 361296 3232 361312 3296
rect 361376 3232 361404 3296
rect 360804 3231 361404 3232
rect 396804 3296 397404 3297
rect 396804 3232 396832 3296
rect 396896 3232 396912 3296
rect 396976 3232 396992 3296
rect 397056 3232 397072 3296
rect 397136 3232 397152 3296
rect 397216 3232 397232 3296
rect 397296 3232 397312 3296
rect 397376 3232 397404 3296
rect 396804 3231 397404 3232
rect 432804 3296 433404 3297
rect 432804 3232 432832 3296
rect 432896 3232 432912 3296
rect 432976 3232 432992 3296
rect 433056 3232 433072 3296
rect 433136 3232 433152 3296
rect 433216 3232 433232 3296
rect 433296 3232 433312 3296
rect 433376 3232 433404 3296
rect 432804 3231 433404 3232
rect 468804 3296 469404 3297
rect 468804 3232 468832 3296
rect 468896 3232 468912 3296
rect 468976 3232 468992 3296
rect 469056 3232 469072 3296
rect 469136 3232 469152 3296
rect 469216 3232 469232 3296
rect 469296 3232 469312 3296
rect 469376 3232 469404 3296
rect 468804 3231 469404 3232
rect 504804 3296 505404 3297
rect 504804 3232 504832 3296
rect 504896 3232 504912 3296
rect 504976 3232 504992 3296
rect 505056 3232 505072 3296
rect 505136 3232 505152 3296
rect 505216 3232 505232 3296
rect 505296 3232 505312 3296
rect 505376 3232 505404 3296
rect 504804 3231 505404 3232
rect 540804 3296 541404 3297
rect 540804 3232 540832 3296
rect 540896 3232 540912 3296
rect 540976 3232 540992 3296
rect 541056 3232 541072 3296
rect 541136 3232 541152 3296
rect 541216 3232 541232 3296
rect 541296 3232 541312 3296
rect 541376 3232 541404 3296
rect 540804 3231 541404 3232
rect 576804 3296 577404 3297
rect 576804 3232 576832 3296
rect 576896 3232 576912 3296
rect 576976 3232 576992 3296
rect 577056 3232 577072 3296
rect 577136 3232 577152 3296
rect 577216 3232 577232 3296
rect 577296 3232 577312 3296
rect 577376 3232 577404 3296
rect 576804 3231 577404 3232
rect 18804 2752 19404 2753
rect 18804 2688 18832 2752
rect 18896 2688 18912 2752
rect 18976 2688 18992 2752
rect 19056 2688 19072 2752
rect 19136 2688 19152 2752
rect 19216 2688 19232 2752
rect 19296 2688 19312 2752
rect 19376 2688 19404 2752
rect 18804 2687 19404 2688
rect 54804 2752 55404 2753
rect 54804 2688 54832 2752
rect 54896 2688 54912 2752
rect 54976 2688 54992 2752
rect 55056 2688 55072 2752
rect 55136 2688 55152 2752
rect 55216 2688 55232 2752
rect 55296 2688 55312 2752
rect 55376 2688 55404 2752
rect 54804 2687 55404 2688
rect 90804 2752 91404 2753
rect 90804 2688 90832 2752
rect 90896 2688 90912 2752
rect 90976 2688 90992 2752
rect 91056 2688 91072 2752
rect 91136 2688 91152 2752
rect 91216 2688 91232 2752
rect 91296 2688 91312 2752
rect 91376 2688 91404 2752
rect 90804 2687 91404 2688
rect 126804 2752 127404 2753
rect 126804 2688 126832 2752
rect 126896 2688 126912 2752
rect 126976 2688 126992 2752
rect 127056 2688 127072 2752
rect 127136 2688 127152 2752
rect 127216 2688 127232 2752
rect 127296 2688 127312 2752
rect 127376 2688 127404 2752
rect 126804 2687 127404 2688
rect 162804 2752 163404 2753
rect 162804 2688 162832 2752
rect 162896 2688 162912 2752
rect 162976 2688 162992 2752
rect 163056 2688 163072 2752
rect 163136 2688 163152 2752
rect 163216 2688 163232 2752
rect 163296 2688 163312 2752
rect 163376 2688 163404 2752
rect 162804 2687 163404 2688
rect 198804 2752 199404 2753
rect 198804 2688 198832 2752
rect 198896 2688 198912 2752
rect 198976 2688 198992 2752
rect 199056 2688 199072 2752
rect 199136 2688 199152 2752
rect 199216 2688 199232 2752
rect 199296 2688 199312 2752
rect 199376 2688 199404 2752
rect 198804 2687 199404 2688
rect 234804 2752 235404 2753
rect 234804 2688 234832 2752
rect 234896 2688 234912 2752
rect 234976 2688 234992 2752
rect 235056 2688 235072 2752
rect 235136 2688 235152 2752
rect 235216 2688 235232 2752
rect 235296 2688 235312 2752
rect 235376 2688 235404 2752
rect 234804 2687 235404 2688
rect 270804 2752 271404 2753
rect 270804 2688 270832 2752
rect 270896 2688 270912 2752
rect 270976 2688 270992 2752
rect 271056 2688 271072 2752
rect 271136 2688 271152 2752
rect 271216 2688 271232 2752
rect 271296 2688 271312 2752
rect 271376 2688 271404 2752
rect 270804 2687 271404 2688
rect 306804 2752 307404 2753
rect 306804 2688 306832 2752
rect 306896 2688 306912 2752
rect 306976 2688 306992 2752
rect 307056 2688 307072 2752
rect 307136 2688 307152 2752
rect 307216 2688 307232 2752
rect 307296 2688 307312 2752
rect 307376 2688 307404 2752
rect 306804 2687 307404 2688
rect 342804 2752 343404 2753
rect 342804 2688 342832 2752
rect 342896 2688 342912 2752
rect 342976 2688 342992 2752
rect 343056 2688 343072 2752
rect 343136 2688 343152 2752
rect 343216 2688 343232 2752
rect 343296 2688 343312 2752
rect 343376 2688 343404 2752
rect 342804 2687 343404 2688
rect 378804 2752 379404 2753
rect 378804 2688 378832 2752
rect 378896 2688 378912 2752
rect 378976 2688 378992 2752
rect 379056 2688 379072 2752
rect 379136 2688 379152 2752
rect 379216 2688 379232 2752
rect 379296 2688 379312 2752
rect 379376 2688 379404 2752
rect 378804 2687 379404 2688
rect 414804 2752 415404 2753
rect 414804 2688 414832 2752
rect 414896 2688 414912 2752
rect 414976 2688 414992 2752
rect 415056 2688 415072 2752
rect 415136 2688 415152 2752
rect 415216 2688 415232 2752
rect 415296 2688 415312 2752
rect 415376 2688 415404 2752
rect 414804 2687 415404 2688
rect 450804 2752 451404 2753
rect 450804 2688 450832 2752
rect 450896 2688 450912 2752
rect 450976 2688 450992 2752
rect 451056 2688 451072 2752
rect 451136 2688 451152 2752
rect 451216 2688 451232 2752
rect 451296 2688 451312 2752
rect 451376 2688 451404 2752
rect 450804 2687 451404 2688
rect 486804 2752 487404 2753
rect 486804 2688 486832 2752
rect 486896 2688 486912 2752
rect 486976 2688 486992 2752
rect 487056 2688 487072 2752
rect 487136 2688 487152 2752
rect 487216 2688 487232 2752
rect 487296 2688 487312 2752
rect 487376 2688 487404 2752
rect 486804 2687 487404 2688
rect 522804 2752 523404 2753
rect 522804 2688 522832 2752
rect 522896 2688 522912 2752
rect 522976 2688 522992 2752
rect 523056 2688 523072 2752
rect 523136 2688 523152 2752
rect 523216 2688 523232 2752
rect 523296 2688 523312 2752
rect 523376 2688 523404 2752
rect 522804 2687 523404 2688
rect 558804 2752 559404 2753
rect 558804 2688 558832 2752
rect 558896 2688 558912 2752
rect 558976 2688 558992 2752
rect 559056 2688 559072 2752
rect 559136 2688 559152 2752
rect 559216 2688 559232 2752
rect 559296 2688 559312 2752
rect 559376 2688 559404 2752
rect 558804 2687 559404 2688
rect 36804 2208 37404 2209
rect 36804 2144 36832 2208
rect 36896 2144 36912 2208
rect 36976 2144 36992 2208
rect 37056 2144 37072 2208
rect 37136 2144 37152 2208
rect 37216 2144 37232 2208
rect 37296 2144 37312 2208
rect 37376 2144 37404 2208
rect 36804 2143 37404 2144
rect 72804 2208 73404 2209
rect 72804 2144 72832 2208
rect 72896 2144 72912 2208
rect 72976 2144 72992 2208
rect 73056 2144 73072 2208
rect 73136 2144 73152 2208
rect 73216 2144 73232 2208
rect 73296 2144 73312 2208
rect 73376 2144 73404 2208
rect 72804 2143 73404 2144
rect 108804 2208 109404 2209
rect 108804 2144 108832 2208
rect 108896 2144 108912 2208
rect 108976 2144 108992 2208
rect 109056 2144 109072 2208
rect 109136 2144 109152 2208
rect 109216 2144 109232 2208
rect 109296 2144 109312 2208
rect 109376 2144 109404 2208
rect 108804 2143 109404 2144
rect 144804 2208 145404 2209
rect 144804 2144 144832 2208
rect 144896 2144 144912 2208
rect 144976 2144 144992 2208
rect 145056 2144 145072 2208
rect 145136 2144 145152 2208
rect 145216 2144 145232 2208
rect 145296 2144 145312 2208
rect 145376 2144 145404 2208
rect 144804 2143 145404 2144
rect 180804 2208 181404 2209
rect 180804 2144 180832 2208
rect 180896 2144 180912 2208
rect 180976 2144 180992 2208
rect 181056 2144 181072 2208
rect 181136 2144 181152 2208
rect 181216 2144 181232 2208
rect 181296 2144 181312 2208
rect 181376 2144 181404 2208
rect 180804 2143 181404 2144
rect 216804 2208 217404 2209
rect 216804 2144 216832 2208
rect 216896 2144 216912 2208
rect 216976 2144 216992 2208
rect 217056 2144 217072 2208
rect 217136 2144 217152 2208
rect 217216 2144 217232 2208
rect 217296 2144 217312 2208
rect 217376 2144 217404 2208
rect 216804 2143 217404 2144
rect 252804 2208 253404 2209
rect 252804 2144 252832 2208
rect 252896 2144 252912 2208
rect 252976 2144 252992 2208
rect 253056 2144 253072 2208
rect 253136 2144 253152 2208
rect 253216 2144 253232 2208
rect 253296 2144 253312 2208
rect 253376 2144 253404 2208
rect 252804 2143 253404 2144
rect 288804 2208 289404 2209
rect 288804 2144 288832 2208
rect 288896 2144 288912 2208
rect 288976 2144 288992 2208
rect 289056 2144 289072 2208
rect 289136 2144 289152 2208
rect 289216 2144 289232 2208
rect 289296 2144 289312 2208
rect 289376 2144 289404 2208
rect 288804 2143 289404 2144
rect 324804 2208 325404 2209
rect 324804 2144 324832 2208
rect 324896 2144 324912 2208
rect 324976 2144 324992 2208
rect 325056 2144 325072 2208
rect 325136 2144 325152 2208
rect 325216 2144 325232 2208
rect 325296 2144 325312 2208
rect 325376 2144 325404 2208
rect 324804 2143 325404 2144
rect 360804 2208 361404 2209
rect 360804 2144 360832 2208
rect 360896 2144 360912 2208
rect 360976 2144 360992 2208
rect 361056 2144 361072 2208
rect 361136 2144 361152 2208
rect 361216 2144 361232 2208
rect 361296 2144 361312 2208
rect 361376 2144 361404 2208
rect 360804 2143 361404 2144
rect 396804 2208 397404 2209
rect 396804 2144 396832 2208
rect 396896 2144 396912 2208
rect 396976 2144 396992 2208
rect 397056 2144 397072 2208
rect 397136 2144 397152 2208
rect 397216 2144 397232 2208
rect 397296 2144 397312 2208
rect 397376 2144 397404 2208
rect 396804 2143 397404 2144
rect 432804 2208 433404 2209
rect 432804 2144 432832 2208
rect 432896 2144 432912 2208
rect 432976 2144 432992 2208
rect 433056 2144 433072 2208
rect 433136 2144 433152 2208
rect 433216 2144 433232 2208
rect 433296 2144 433312 2208
rect 433376 2144 433404 2208
rect 432804 2143 433404 2144
rect 468804 2208 469404 2209
rect 468804 2144 468832 2208
rect 468896 2144 468912 2208
rect 468976 2144 468992 2208
rect 469056 2144 469072 2208
rect 469136 2144 469152 2208
rect 469216 2144 469232 2208
rect 469296 2144 469312 2208
rect 469376 2144 469404 2208
rect 468804 2143 469404 2144
rect 504804 2208 505404 2209
rect 504804 2144 504832 2208
rect 504896 2144 504912 2208
rect 504976 2144 504992 2208
rect 505056 2144 505072 2208
rect 505136 2144 505152 2208
rect 505216 2144 505232 2208
rect 505296 2144 505312 2208
rect 505376 2144 505404 2208
rect 504804 2143 505404 2144
rect 540804 2208 541404 2209
rect 540804 2144 540832 2208
rect 540896 2144 540912 2208
rect 540976 2144 540992 2208
rect 541056 2144 541072 2208
rect 541136 2144 541152 2208
rect 541216 2144 541232 2208
rect 541296 2144 541312 2208
rect 541376 2144 541404 2208
rect 540804 2143 541404 2144
rect 576804 2208 577404 2209
rect 576804 2144 576832 2208
rect 576896 2144 576912 2208
rect 576976 2144 576992 2208
rect 577056 2144 577072 2208
rect 577136 2144 577152 2208
rect 577216 2144 577232 2208
rect 577296 2144 577312 2208
rect 577376 2144 577404 2208
rect 576804 2143 577404 2144
<< via3 >>
rect 36832 701788 36896 701792
rect 36832 701732 36836 701788
rect 36836 701732 36892 701788
rect 36892 701732 36896 701788
rect 36832 701728 36896 701732
rect 36912 701788 36976 701792
rect 36912 701732 36916 701788
rect 36916 701732 36972 701788
rect 36972 701732 36976 701788
rect 36912 701728 36976 701732
rect 36992 701788 37056 701792
rect 36992 701732 36996 701788
rect 36996 701732 37052 701788
rect 37052 701732 37056 701788
rect 36992 701728 37056 701732
rect 37072 701788 37136 701792
rect 37072 701732 37076 701788
rect 37076 701732 37132 701788
rect 37132 701732 37136 701788
rect 37072 701728 37136 701732
rect 37152 701788 37216 701792
rect 37152 701732 37156 701788
rect 37156 701732 37212 701788
rect 37212 701732 37216 701788
rect 37152 701728 37216 701732
rect 37232 701788 37296 701792
rect 37232 701732 37236 701788
rect 37236 701732 37292 701788
rect 37292 701732 37296 701788
rect 37232 701728 37296 701732
rect 37312 701788 37376 701792
rect 37312 701732 37316 701788
rect 37316 701732 37372 701788
rect 37372 701732 37376 701788
rect 37312 701728 37376 701732
rect 72832 701788 72896 701792
rect 72832 701732 72836 701788
rect 72836 701732 72892 701788
rect 72892 701732 72896 701788
rect 72832 701728 72896 701732
rect 72912 701788 72976 701792
rect 72912 701732 72916 701788
rect 72916 701732 72972 701788
rect 72972 701732 72976 701788
rect 72912 701728 72976 701732
rect 72992 701788 73056 701792
rect 72992 701732 72996 701788
rect 72996 701732 73052 701788
rect 73052 701732 73056 701788
rect 72992 701728 73056 701732
rect 73072 701788 73136 701792
rect 73072 701732 73076 701788
rect 73076 701732 73132 701788
rect 73132 701732 73136 701788
rect 73072 701728 73136 701732
rect 73152 701788 73216 701792
rect 73152 701732 73156 701788
rect 73156 701732 73212 701788
rect 73212 701732 73216 701788
rect 73152 701728 73216 701732
rect 73232 701788 73296 701792
rect 73232 701732 73236 701788
rect 73236 701732 73292 701788
rect 73292 701732 73296 701788
rect 73232 701728 73296 701732
rect 73312 701788 73376 701792
rect 73312 701732 73316 701788
rect 73316 701732 73372 701788
rect 73372 701732 73376 701788
rect 73312 701728 73376 701732
rect 108832 701788 108896 701792
rect 108832 701732 108836 701788
rect 108836 701732 108892 701788
rect 108892 701732 108896 701788
rect 108832 701728 108896 701732
rect 108912 701788 108976 701792
rect 108912 701732 108916 701788
rect 108916 701732 108972 701788
rect 108972 701732 108976 701788
rect 108912 701728 108976 701732
rect 108992 701788 109056 701792
rect 108992 701732 108996 701788
rect 108996 701732 109052 701788
rect 109052 701732 109056 701788
rect 108992 701728 109056 701732
rect 109072 701788 109136 701792
rect 109072 701732 109076 701788
rect 109076 701732 109132 701788
rect 109132 701732 109136 701788
rect 109072 701728 109136 701732
rect 109152 701788 109216 701792
rect 109152 701732 109156 701788
rect 109156 701732 109212 701788
rect 109212 701732 109216 701788
rect 109152 701728 109216 701732
rect 109232 701788 109296 701792
rect 109232 701732 109236 701788
rect 109236 701732 109292 701788
rect 109292 701732 109296 701788
rect 109232 701728 109296 701732
rect 109312 701788 109376 701792
rect 109312 701732 109316 701788
rect 109316 701732 109372 701788
rect 109372 701732 109376 701788
rect 109312 701728 109376 701732
rect 144832 701788 144896 701792
rect 144832 701732 144836 701788
rect 144836 701732 144892 701788
rect 144892 701732 144896 701788
rect 144832 701728 144896 701732
rect 144912 701788 144976 701792
rect 144912 701732 144916 701788
rect 144916 701732 144972 701788
rect 144972 701732 144976 701788
rect 144912 701728 144976 701732
rect 144992 701788 145056 701792
rect 144992 701732 144996 701788
rect 144996 701732 145052 701788
rect 145052 701732 145056 701788
rect 144992 701728 145056 701732
rect 145072 701788 145136 701792
rect 145072 701732 145076 701788
rect 145076 701732 145132 701788
rect 145132 701732 145136 701788
rect 145072 701728 145136 701732
rect 145152 701788 145216 701792
rect 145152 701732 145156 701788
rect 145156 701732 145212 701788
rect 145212 701732 145216 701788
rect 145152 701728 145216 701732
rect 145232 701788 145296 701792
rect 145232 701732 145236 701788
rect 145236 701732 145292 701788
rect 145292 701732 145296 701788
rect 145232 701728 145296 701732
rect 145312 701788 145376 701792
rect 145312 701732 145316 701788
rect 145316 701732 145372 701788
rect 145372 701732 145376 701788
rect 145312 701728 145376 701732
rect 180832 701788 180896 701792
rect 180832 701732 180836 701788
rect 180836 701732 180892 701788
rect 180892 701732 180896 701788
rect 180832 701728 180896 701732
rect 180912 701788 180976 701792
rect 180912 701732 180916 701788
rect 180916 701732 180972 701788
rect 180972 701732 180976 701788
rect 180912 701728 180976 701732
rect 180992 701788 181056 701792
rect 180992 701732 180996 701788
rect 180996 701732 181052 701788
rect 181052 701732 181056 701788
rect 180992 701728 181056 701732
rect 181072 701788 181136 701792
rect 181072 701732 181076 701788
rect 181076 701732 181132 701788
rect 181132 701732 181136 701788
rect 181072 701728 181136 701732
rect 181152 701788 181216 701792
rect 181152 701732 181156 701788
rect 181156 701732 181212 701788
rect 181212 701732 181216 701788
rect 181152 701728 181216 701732
rect 181232 701788 181296 701792
rect 181232 701732 181236 701788
rect 181236 701732 181292 701788
rect 181292 701732 181296 701788
rect 181232 701728 181296 701732
rect 181312 701788 181376 701792
rect 181312 701732 181316 701788
rect 181316 701732 181372 701788
rect 181372 701732 181376 701788
rect 181312 701728 181376 701732
rect 216832 701788 216896 701792
rect 216832 701732 216836 701788
rect 216836 701732 216892 701788
rect 216892 701732 216896 701788
rect 216832 701728 216896 701732
rect 216912 701788 216976 701792
rect 216912 701732 216916 701788
rect 216916 701732 216972 701788
rect 216972 701732 216976 701788
rect 216912 701728 216976 701732
rect 216992 701788 217056 701792
rect 216992 701732 216996 701788
rect 216996 701732 217052 701788
rect 217052 701732 217056 701788
rect 216992 701728 217056 701732
rect 217072 701788 217136 701792
rect 217072 701732 217076 701788
rect 217076 701732 217132 701788
rect 217132 701732 217136 701788
rect 217072 701728 217136 701732
rect 217152 701788 217216 701792
rect 217152 701732 217156 701788
rect 217156 701732 217212 701788
rect 217212 701732 217216 701788
rect 217152 701728 217216 701732
rect 217232 701788 217296 701792
rect 217232 701732 217236 701788
rect 217236 701732 217292 701788
rect 217292 701732 217296 701788
rect 217232 701728 217296 701732
rect 217312 701788 217376 701792
rect 217312 701732 217316 701788
rect 217316 701732 217372 701788
rect 217372 701732 217376 701788
rect 217312 701728 217376 701732
rect 252832 701788 252896 701792
rect 252832 701732 252836 701788
rect 252836 701732 252892 701788
rect 252892 701732 252896 701788
rect 252832 701728 252896 701732
rect 252912 701788 252976 701792
rect 252912 701732 252916 701788
rect 252916 701732 252972 701788
rect 252972 701732 252976 701788
rect 252912 701728 252976 701732
rect 252992 701788 253056 701792
rect 252992 701732 252996 701788
rect 252996 701732 253052 701788
rect 253052 701732 253056 701788
rect 252992 701728 253056 701732
rect 253072 701788 253136 701792
rect 253072 701732 253076 701788
rect 253076 701732 253132 701788
rect 253132 701732 253136 701788
rect 253072 701728 253136 701732
rect 253152 701788 253216 701792
rect 253152 701732 253156 701788
rect 253156 701732 253212 701788
rect 253212 701732 253216 701788
rect 253152 701728 253216 701732
rect 253232 701788 253296 701792
rect 253232 701732 253236 701788
rect 253236 701732 253292 701788
rect 253292 701732 253296 701788
rect 253232 701728 253296 701732
rect 253312 701788 253376 701792
rect 253312 701732 253316 701788
rect 253316 701732 253372 701788
rect 253372 701732 253376 701788
rect 253312 701728 253376 701732
rect 288832 701788 288896 701792
rect 288832 701732 288836 701788
rect 288836 701732 288892 701788
rect 288892 701732 288896 701788
rect 288832 701728 288896 701732
rect 288912 701788 288976 701792
rect 288912 701732 288916 701788
rect 288916 701732 288972 701788
rect 288972 701732 288976 701788
rect 288912 701728 288976 701732
rect 288992 701788 289056 701792
rect 288992 701732 288996 701788
rect 288996 701732 289052 701788
rect 289052 701732 289056 701788
rect 288992 701728 289056 701732
rect 289072 701788 289136 701792
rect 289072 701732 289076 701788
rect 289076 701732 289132 701788
rect 289132 701732 289136 701788
rect 289072 701728 289136 701732
rect 289152 701788 289216 701792
rect 289152 701732 289156 701788
rect 289156 701732 289212 701788
rect 289212 701732 289216 701788
rect 289152 701728 289216 701732
rect 289232 701788 289296 701792
rect 289232 701732 289236 701788
rect 289236 701732 289292 701788
rect 289292 701732 289296 701788
rect 289232 701728 289296 701732
rect 289312 701788 289376 701792
rect 289312 701732 289316 701788
rect 289316 701732 289372 701788
rect 289372 701732 289376 701788
rect 289312 701728 289376 701732
rect 324832 701788 324896 701792
rect 324832 701732 324836 701788
rect 324836 701732 324892 701788
rect 324892 701732 324896 701788
rect 324832 701728 324896 701732
rect 324912 701788 324976 701792
rect 324912 701732 324916 701788
rect 324916 701732 324972 701788
rect 324972 701732 324976 701788
rect 324912 701728 324976 701732
rect 324992 701788 325056 701792
rect 324992 701732 324996 701788
rect 324996 701732 325052 701788
rect 325052 701732 325056 701788
rect 324992 701728 325056 701732
rect 325072 701788 325136 701792
rect 325072 701732 325076 701788
rect 325076 701732 325132 701788
rect 325132 701732 325136 701788
rect 325072 701728 325136 701732
rect 325152 701788 325216 701792
rect 325152 701732 325156 701788
rect 325156 701732 325212 701788
rect 325212 701732 325216 701788
rect 325152 701728 325216 701732
rect 325232 701788 325296 701792
rect 325232 701732 325236 701788
rect 325236 701732 325292 701788
rect 325292 701732 325296 701788
rect 325232 701728 325296 701732
rect 325312 701788 325376 701792
rect 325312 701732 325316 701788
rect 325316 701732 325372 701788
rect 325372 701732 325376 701788
rect 325312 701728 325376 701732
rect 360832 701788 360896 701792
rect 360832 701732 360836 701788
rect 360836 701732 360892 701788
rect 360892 701732 360896 701788
rect 360832 701728 360896 701732
rect 360912 701788 360976 701792
rect 360912 701732 360916 701788
rect 360916 701732 360972 701788
rect 360972 701732 360976 701788
rect 360912 701728 360976 701732
rect 360992 701788 361056 701792
rect 360992 701732 360996 701788
rect 360996 701732 361052 701788
rect 361052 701732 361056 701788
rect 360992 701728 361056 701732
rect 361072 701788 361136 701792
rect 361072 701732 361076 701788
rect 361076 701732 361132 701788
rect 361132 701732 361136 701788
rect 361072 701728 361136 701732
rect 361152 701788 361216 701792
rect 361152 701732 361156 701788
rect 361156 701732 361212 701788
rect 361212 701732 361216 701788
rect 361152 701728 361216 701732
rect 361232 701788 361296 701792
rect 361232 701732 361236 701788
rect 361236 701732 361292 701788
rect 361292 701732 361296 701788
rect 361232 701728 361296 701732
rect 361312 701788 361376 701792
rect 361312 701732 361316 701788
rect 361316 701732 361372 701788
rect 361372 701732 361376 701788
rect 361312 701728 361376 701732
rect 396832 701788 396896 701792
rect 396832 701732 396836 701788
rect 396836 701732 396892 701788
rect 396892 701732 396896 701788
rect 396832 701728 396896 701732
rect 396912 701788 396976 701792
rect 396912 701732 396916 701788
rect 396916 701732 396972 701788
rect 396972 701732 396976 701788
rect 396912 701728 396976 701732
rect 396992 701788 397056 701792
rect 396992 701732 396996 701788
rect 396996 701732 397052 701788
rect 397052 701732 397056 701788
rect 396992 701728 397056 701732
rect 397072 701788 397136 701792
rect 397072 701732 397076 701788
rect 397076 701732 397132 701788
rect 397132 701732 397136 701788
rect 397072 701728 397136 701732
rect 397152 701788 397216 701792
rect 397152 701732 397156 701788
rect 397156 701732 397212 701788
rect 397212 701732 397216 701788
rect 397152 701728 397216 701732
rect 397232 701788 397296 701792
rect 397232 701732 397236 701788
rect 397236 701732 397292 701788
rect 397292 701732 397296 701788
rect 397232 701728 397296 701732
rect 397312 701788 397376 701792
rect 397312 701732 397316 701788
rect 397316 701732 397372 701788
rect 397372 701732 397376 701788
rect 397312 701728 397376 701732
rect 432832 701788 432896 701792
rect 432832 701732 432836 701788
rect 432836 701732 432892 701788
rect 432892 701732 432896 701788
rect 432832 701728 432896 701732
rect 432912 701788 432976 701792
rect 432912 701732 432916 701788
rect 432916 701732 432972 701788
rect 432972 701732 432976 701788
rect 432912 701728 432976 701732
rect 432992 701788 433056 701792
rect 432992 701732 432996 701788
rect 432996 701732 433052 701788
rect 433052 701732 433056 701788
rect 432992 701728 433056 701732
rect 433072 701788 433136 701792
rect 433072 701732 433076 701788
rect 433076 701732 433132 701788
rect 433132 701732 433136 701788
rect 433072 701728 433136 701732
rect 433152 701788 433216 701792
rect 433152 701732 433156 701788
rect 433156 701732 433212 701788
rect 433212 701732 433216 701788
rect 433152 701728 433216 701732
rect 433232 701788 433296 701792
rect 433232 701732 433236 701788
rect 433236 701732 433292 701788
rect 433292 701732 433296 701788
rect 433232 701728 433296 701732
rect 433312 701788 433376 701792
rect 433312 701732 433316 701788
rect 433316 701732 433372 701788
rect 433372 701732 433376 701788
rect 433312 701728 433376 701732
rect 468832 701788 468896 701792
rect 468832 701732 468836 701788
rect 468836 701732 468892 701788
rect 468892 701732 468896 701788
rect 468832 701728 468896 701732
rect 468912 701788 468976 701792
rect 468912 701732 468916 701788
rect 468916 701732 468972 701788
rect 468972 701732 468976 701788
rect 468912 701728 468976 701732
rect 468992 701788 469056 701792
rect 468992 701732 468996 701788
rect 468996 701732 469052 701788
rect 469052 701732 469056 701788
rect 468992 701728 469056 701732
rect 469072 701788 469136 701792
rect 469072 701732 469076 701788
rect 469076 701732 469132 701788
rect 469132 701732 469136 701788
rect 469072 701728 469136 701732
rect 469152 701788 469216 701792
rect 469152 701732 469156 701788
rect 469156 701732 469212 701788
rect 469212 701732 469216 701788
rect 469152 701728 469216 701732
rect 469232 701788 469296 701792
rect 469232 701732 469236 701788
rect 469236 701732 469292 701788
rect 469292 701732 469296 701788
rect 469232 701728 469296 701732
rect 469312 701788 469376 701792
rect 469312 701732 469316 701788
rect 469316 701732 469372 701788
rect 469372 701732 469376 701788
rect 469312 701728 469376 701732
rect 504832 701788 504896 701792
rect 504832 701732 504836 701788
rect 504836 701732 504892 701788
rect 504892 701732 504896 701788
rect 504832 701728 504896 701732
rect 504912 701788 504976 701792
rect 504912 701732 504916 701788
rect 504916 701732 504972 701788
rect 504972 701732 504976 701788
rect 504912 701728 504976 701732
rect 504992 701788 505056 701792
rect 504992 701732 504996 701788
rect 504996 701732 505052 701788
rect 505052 701732 505056 701788
rect 504992 701728 505056 701732
rect 505072 701788 505136 701792
rect 505072 701732 505076 701788
rect 505076 701732 505132 701788
rect 505132 701732 505136 701788
rect 505072 701728 505136 701732
rect 505152 701788 505216 701792
rect 505152 701732 505156 701788
rect 505156 701732 505212 701788
rect 505212 701732 505216 701788
rect 505152 701728 505216 701732
rect 505232 701788 505296 701792
rect 505232 701732 505236 701788
rect 505236 701732 505292 701788
rect 505292 701732 505296 701788
rect 505232 701728 505296 701732
rect 505312 701788 505376 701792
rect 505312 701732 505316 701788
rect 505316 701732 505372 701788
rect 505372 701732 505376 701788
rect 505312 701728 505376 701732
rect 540832 701788 540896 701792
rect 540832 701732 540836 701788
rect 540836 701732 540892 701788
rect 540892 701732 540896 701788
rect 540832 701728 540896 701732
rect 540912 701788 540976 701792
rect 540912 701732 540916 701788
rect 540916 701732 540972 701788
rect 540972 701732 540976 701788
rect 540912 701728 540976 701732
rect 540992 701788 541056 701792
rect 540992 701732 540996 701788
rect 540996 701732 541052 701788
rect 541052 701732 541056 701788
rect 540992 701728 541056 701732
rect 541072 701788 541136 701792
rect 541072 701732 541076 701788
rect 541076 701732 541132 701788
rect 541132 701732 541136 701788
rect 541072 701728 541136 701732
rect 541152 701788 541216 701792
rect 541152 701732 541156 701788
rect 541156 701732 541212 701788
rect 541212 701732 541216 701788
rect 541152 701728 541216 701732
rect 541232 701788 541296 701792
rect 541232 701732 541236 701788
rect 541236 701732 541292 701788
rect 541292 701732 541296 701788
rect 541232 701728 541296 701732
rect 541312 701788 541376 701792
rect 541312 701732 541316 701788
rect 541316 701732 541372 701788
rect 541372 701732 541376 701788
rect 541312 701728 541376 701732
rect 576832 701788 576896 701792
rect 576832 701732 576836 701788
rect 576836 701732 576892 701788
rect 576892 701732 576896 701788
rect 576832 701728 576896 701732
rect 576912 701788 576976 701792
rect 576912 701732 576916 701788
rect 576916 701732 576972 701788
rect 576972 701732 576976 701788
rect 576912 701728 576976 701732
rect 576992 701788 577056 701792
rect 576992 701732 576996 701788
rect 576996 701732 577052 701788
rect 577052 701732 577056 701788
rect 576992 701728 577056 701732
rect 577072 701788 577136 701792
rect 577072 701732 577076 701788
rect 577076 701732 577132 701788
rect 577132 701732 577136 701788
rect 577072 701728 577136 701732
rect 577152 701788 577216 701792
rect 577152 701732 577156 701788
rect 577156 701732 577212 701788
rect 577212 701732 577216 701788
rect 577152 701728 577216 701732
rect 577232 701788 577296 701792
rect 577232 701732 577236 701788
rect 577236 701732 577292 701788
rect 577292 701732 577296 701788
rect 577232 701728 577296 701732
rect 577312 701788 577376 701792
rect 577312 701732 577316 701788
rect 577316 701732 577372 701788
rect 577372 701732 577376 701788
rect 577312 701728 577376 701732
rect 18832 701244 18896 701248
rect 18832 701188 18836 701244
rect 18836 701188 18892 701244
rect 18892 701188 18896 701244
rect 18832 701184 18896 701188
rect 18912 701244 18976 701248
rect 18912 701188 18916 701244
rect 18916 701188 18972 701244
rect 18972 701188 18976 701244
rect 18912 701184 18976 701188
rect 18992 701244 19056 701248
rect 18992 701188 18996 701244
rect 18996 701188 19052 701244
rect 19052 701188 19056 701244
rect 18992 701184 19056 701188
rect 19072 701244 19136 701248
rect 19072 701188 19076 701244
rect 19076 701188 19132 701244
rect 19132 701188 19136 701244
rect 19072 701184 19136 701188
rect 19152 701244 19216 701248
rect 19152 701188 19156 701244
rect 19156 701188 19212 701244
rect 19212 701188 19216 701244
rect 19152 701184 19216 701188
rect 19232 701244 19296 701248
rect 19232 701188 19236 701244
rect 19236 701188 19292 701244
rect 19292 701188 19296 701244
rect 19232 701184 19296 701188
rect 19312 701244 19376 701248
rect 19312 701188 19316 701244
rect 19316 701188 19372 701244
rect 19372 701188 19376 701244
rect 19312 701184 19376 701188
rect 54832 701244 54896 701248
rect 54832 701188 54836 701244
rect 54836 701188 54892 701244
rect 54892 701188 54896 701244
rect 54832 701184 54896 701188
rect 54912 701244 54976 701248
rect 54912 701188 54916 701244
rect 54916 701188 54972 701244
rect 54972 701188 54976 701244
rect 54912 701184 54976 701188
rect 54992 701244 55056 701248
rect 54992 701188 54996 701244
rect 54996 701188 55052 701244
rect 55052 701188 55056 701244
rect 54992 701184 55056 701188
rect 55072 701244 55136 701248
rect 55072 701188 55076 701244
rect 55076 701188 55132 701244
rect 55132 701188 55136 701244
rect 55072 701184 55136 701188
rect 55152 701244 55216 701248
rect 55152 701188 55156 701244
rect 55156 701188 55212 701244
rect 55212 701188 55216 701244
rect 55152 701184 55216 701188
rect 55232 701244 55296 701248
rect 55232 701188 55236 701244
rect 55236 701188 55292 701244
rect 55292 701188 55296 701244
rect 55232 701184 55296 701188
rect 55312 701244 55376 701248
rect 55312 701188 55316 701244
rect 55316 701188 55372 701244
rect 55372 701188 55376 701244
rect 55312 701184 55376 701188
rect 90832 701244 90896 701248
rect 90832 701188 90836 701244
rect 90836 701188 90892 701244
rect 90892 701188 90896 701244
rect 90832 701184 90896 701188
rect 90912 701244 90976 701248
rect 90912 701188 90916 701244
rect 90916 701188 90972 701244
rect 90972 701188 90976 701244
rect 90912 701184 90976 701188
rect 90992 701244 91056 701248
rect 90992 701188 90996 701244
rect 90996 701188 91052 701244
rect 91052 701188 91056 701244
rect 90992 701184 91056 701188
rect 91072 701244 91136 701248
rect 91072 701188 91076 701244
rect 91076 701188 91132 701244
rect 91132 701188 91136 701244
rect 91072 701184 91136 701188
rect 91152 701244 91216 701248
rect 91152 701188 91156 701244
rect 91156 701188 91212 701244
rect 91212 701188 91216 701244
rect 91152 701184 91216 701188
rect 91232 701244 91296 701248
rect 91232 701188 91236 701244
rect 91236 701188 91292 701244
rect 91292 701188 91296 701244
rect 91232 701184 91296 701188
rect 91312 701244 91376 701248
rect 91312 701188 91316 701244
rect 91316 701188 91372 701244
rect 91372 701188 91376 701244
rect 91312 701184 91376 701188
rect 126832 701244 126896 701248
rect 126832 701188 126836 701244
rect 126836 701188 126892 701244
rect 126892 701188 126896 701244
rect 126832 701184 126896 701188
rect 126912 701244 126976 701248
rect 126912 701188 126916 701244
rect 126916 701188 126972 701244
rect 126972 701188 126976 701244
rect 126912 701184 126976 701188
rect 126992 701244 127056 701248
rect 126992 701188 126996 701244
rect 126996 701188 127052 701244
rect 127052 701188 127056 701244
rect 126992 701184 127056 701188
rect 127072 701244 127136 701248
rect 127072 701188 127076 701244
rect 127076 701188 127132 701244
rect 127132 701188 127136 701244
rect 127072 701184 127136 701188
rect 127152 701244 127216 701248
rect 127152 701188 127156 701244
rect 127156 701188 127212 701244
rect 127212 701188 127216 701244
rect 127152 701184 127216 701188
rect 127232 701244 127296 701248
rect 127232 701188 127236 701244
rect 127236 701188 127292 701244
rect 127292 701188 127296 701244
rect 127232 701184 127296 701188
rect 127312 701244 127376 701248
rect 127312 701188 127316 701244
rect 127316 701188 127372 701244
rect 127372 701188 127376 701244
rect 127312 701184 127376 701188
rect 162832 701244 162896 701248
rect 162832 701188 162836 701244
rect 162836 701188 162892 701244
rect 162892 701188 162896 701244
rect 162832 701184 162896 701188
rect 162912 701244 162976 701248
rect 162912 701188 162916 701244
rect 162916 701188 162972 701244
rect 162972 701188 162976 701244
rect 162912 701184 162976 701188
rect 162992 701244 163056 701248
rect 162992 701188 162996 701244
rect 162996 701188 163052 701244
rect 163052 701188 163056 701244
rect 162992 701184 163056 701188
rect 163072 701244 163136 701248
rect 163072 701188 163076 701244
rect 163076 701188 163132 701244
rect 163132 701188 163136 701244
rect 163072 701184 163136 701188
rect 163152 701244 163216 701248
rect 163152 701188 163156 701244
rect 163156 701188 163212 701244
rect 163212 701188 163216 701244
rect 163152 701184 163216 701188
rect 163232 701244 163296 701248
rect 163232 701188 163236 701244
rect 163236 701188 163292 701244
rect 163292 701188 163296 701244
rect 163232 701184 163296 701188
rect 163312 701244 163376 701248
rect 163312 701188 163316 701244
rect 163316 701188 163372 701244
rect 163372 701188 163376 701244
rect 163312 701184 163376 701188
rect 198832 701244 198896 701248
rect 198832 701188 198836 701244
rect 198836 701188 198892 701244
rect 198892 701188 198896 701244
rect 198832 701184 198896 701188
rect 198912 701244 198976 701248
rect 198912 701188 198916 701244
rect 198916 701188 198972 701244
rect 198972 701188 198976 701244
rect 198912 701184 198976 701188
rect 198992 701244 199056 701248
rect 198992 701188 198996 701244
rect 198996 701188 199052 701244
rect 199052 701188 199056 701244
rect 198992 701184 199056 701188
rect 199072 701244 199136 701248
rect 199072 701188 199076 701244
rect 199076 701188 199132 701244
rect 199132 701188 199136 701244
rect 199072 701184 199136 701188
rect 199152 701244 199216 701248
rect 199152 701188 199156 701244
rect 199156 701188 199212 701244
rect 199212 701188 199216 701244
rect 199152 701184 199216 701188
rect 199232 701244 199296 701248
rect 199232 701188 199236 701244
rect 199236 701188 199292 701244
rect 199292 701188 199296 701244
rect 199232 701184 199296 701188
rect 199312 701244 199376 701248
rect 199312 701188 199316 701244
rect 199316 701188 199372 701244
rect 199372 701188 199376 701244
rect 199312 701184 199376 701188
rect 234832 701244 234896 701248
rect 234832 701188 234836 701244
rect 234836 701188 234892 701244
rect 234892 701188 234896 701244
rect 234832 701184 234896 701188
rect 234912 701244 234976 701248
rect 234912 701188 234916 701244
rect 234916 701188 234972 701244
rect 234972 701188 234976 701244
rect 234912 701184 234976 701188
rect 234992 701244 235056 701248
rect 234992 701188 234996 701244
rect 234996 701188 235052 701244
rect 235052 701188 235056 701244
rect 234992 701184 235056 701188
rect 235072 701244 235136 701248
rect 235072 701188 235076 701244
rect 235076 701188 235132 701244
rect 235132 701188 235136 701244
rect 235072 701184 235136 701188
rect 235152 701244 235216 701248
rect 235152 701188 235156 701244
rect 235156 701188 235212 701244
rect 235212 701188 235216 701244
rect 235152 701184 235216 701188
rect 235232 701244 235296 701248
rect 235232 701188 235236 701244
rect 235236 701188 235292 701244
rect 235292 701188 235296 701244
rect 235232 701184 235296 701188
rect 235312 701244 235376 701248
rect 235312 701188 235316 701244
rect 235316 701188 235372 701244
rect 235372 701188 235376 701244
rect 235312 701184 235376 701188
rect 270832 701244 270896 701248
rect 270832 701188 270836 701244
rect 270836 701188 270892 701244
rect 270892 701188 270896 701244
rect 270832 701184 270896 701188
rect 270912 701244 270976 701248
rect 270912 701188 270916 701244
rect 270916 701188 270972 701244
rect 270972 701188 270976 701244
rect 270912 701184 270976 701188
rect 270992 701244 271056 701248
rect 270992 701188 270996 701244
rect 270996 701188 271052 701244
rect 271052 701188 271056 701244
rect 270992 701184 271056 701188
rect 271072 701244 271136 701248
rect 271072 701188 271076 701244
rect 271076 701188 271132 701244
rect 271132 701188 271136 701244
rect 271072 701184 271136 701188
rect 271152 701244 271216 701248
rect 271152 701188 271156 701244
rect 271156 701188 271212 701244
rect 271212 701188 271216 701244
rect 271152 701184 271216 701188
rect 271232 701244 271296 701248
rect 271232 701188 271236 701244
rect 271236 701188 271292 701244
rect 271292 701188 271296 701244
rect 271232 701184 271296 701188
rect 271312 701244 271376 701248
rect 271312 701188 271316 701244
rect 271316 701188 271372 701244
rect 271372 701188 271376 701244
rect 271312 701184 271376 701188
rect 306832 701244 306896 701248
rect 306832 701188 306836 701244
rect 306836 701188 306892 701244
rect 306892 701188 306896 701244
rect 306832 701184 306896 701188
rect 306912 701244 306976 701248
rect 306912 701188 306916 701244
rect 306916 701188 306972 701244
rect 306972 701188 306976 701244
rect 306912 701184 306976 701188
rect 306992 701244 307056 701248
rect 306992 701188 306996 701244
rect 306996 701188 307052 701244
rect 307052 701188 307056 701244
rect 306992 701184 307056 701188
rect 307072 701244 307136 701248
rect 307072 701188 307076 701244
rect 307076 701188 307132 701244
rect 307132 701188 307136 701244
rect 307072 701184 307136 701188
rect 307152 701244 307216 701248
rect 307152 701188 307156 701244
rect 307156 701188 307212 701244
rect 307212 701188 307216 701244
rect 307152 701184 307216 701188
rect 307232 701244 307296 701248
rect 307232 701188 307236 701244
rect 307236 701188 307292 701244
rect 307292 701188 307296 701244
rect 307232 701184 307296 701188
rect 307312 701244 307376 701248
rect 307312 701188 307316 701244
rect 307316 701188 307372 701244
rect 307372 701188 307376 701244
rect 307312 701184 307376 701188
rect 342832 701244 342896 701248
rect 342832 701188 342836 701244
rect 342836 701188 342892 701244
rect 342892 701188 342896 701244
rect 342832 701184 342896 701188
rect 342912 701244 342976 701248
rect 342912 701188 342916 701244
rect 342916 701188 342972 701244
rect 342972 701188 342976 701244
rect 342912 701184 342976 701188
rect 342992 701244 343056 701248
rect 342992 701188 342996 701244
rect 342996 701188 343052 701244
rect 343052 701188 343056 701244
rect 342992 701184 343056 701188
rect 343072 701244 343136 701248
rect 343072 701188 343076 701244
rect 343076 701188 343132 701244
rect 343132 701188 343136 701244
rect 343072 701184 343136 701188
rect 343152 701244 343216 701248
rect 343152 701188 343156 701244
rect 343156 701188 343212 701244
rect 343212 701188 343216 701244
rect 343152 701184 343216 701188
rect 343232 701244 343296 701248
rect 343232 701188 343236 701244
rect 343236 701188 343292 701244
rect 343292 701188 343296 701244
rect 343232 701184 343296 701188
rect 343312 701244 343376 701248
rect 343312 701188 343316 701244
rect 343316 701188 343372 701244
rect 343372 701188 343376 701244
rect 343312 701184 343376 701188
rect 378832 701244 378896 701248
rect 378832 701188 378836 701244
rect 378836 701188 378892 701244
rect 378892 701188 378896 701244
rect 378832 701184 378896 701188
rect 378912 701244 378976 701248
rect 378912 701188 378916 701244
rect 378916 701188 378972 701244
rect 378972 701188 378976 701244
rect 378912 701184 378976 701188
rect 378992 701244 379056 701248
rect 378992 701188 378996 701244
rect 378996 701188 379052 701244
rect 379052 701188 379056 701244
rect 378992 701184 379056 701188
rect 379072 701244 379136 701248
rect 379072 701188 379076 701244
rect 379076 701188 379132 701244
rect 379132 701188 379136 701244
rect 379072 701184 379136 701188
rect 379152 701244 379216 701248
rect 379152 701188 379156 701244
rect 379156 701188 379212 701244
rect 379212 701188 379216 701244
rect 379152 701184 379216 701188
rect 379232 701244 379296 701248
rect 379232 701188 379236 701244
rect 379236 701188 379292 701244
rect 379292 701188 379296 701244
rect 379232 701184 379296 701188
rect 379312 701244 379376 701248
rect 379312 701188 379316 701244
rect 379316 701188 379372 701244
rect 379372 701188 379376 701244
rect 379312 701184 379376 701188
rect 414832 701244 414896 701248
rect 414832 701188 414836 701244
rect 414836 701188 414892 701244
rect 414892 701188 414896 701244
rect 414832 701184 414896 701188
rect 414912 701244 414976 701248
rect 414912 701188 414916 701244
rect 414916 701188 414972 701244
rect 414972 701188 414976 701244
rect 414912 701184 414976 701188
rect 414992 701244 415056 701248
rect 414992 701188 414996 701244
rect 414996 701188 415052 701244
rect 415052 701188 415056 701244
rect 414992 701184 415056 701188
rect 415072 701244 415136 701248
rect 415072 701188 415076 701244
rect 415076 701188 415132 701244
rect 415132 701188 415136 701244
rect 415072 701184 415136 701188
rect 415152 701244 415216 701248
rect 415152 701188 415156 701244
rect 415156 701188 415212 701244
rect 415212 701188 415216 701244
rect 415152 701184 415216 701188
rect 415232 701244 415296 701248
rect 415232 701188 415236 701244
rect 415236 701188 415292 701244
rect 415292 701188 415296 701244
rect 415232 701184 415296 701188
rect 415312 701244 415376 701248
rect 415312 701188 415316 701244
rect 415316 701188 415372 701244
rect 415372 701188 415376 701244
rect 415312 701184 415376 701188
rect 450832 701244 450896 701248
rect 450832 701188 450836 701244
rect 450836 701188 450892 701244
rect 450892 701188 450896 701244
rect 450832 701184 450896 701188
rect 450912 701244 450976 701248
rect 450912 701188 450916 701244
rect 450916 701188 450972 701244
rect 450972 701188 450976 701244
rect 450912 701184 450976 701188
rect 450992 701244 451056 701248
rect 450992 701188 450996 701244
rect 450996 701188 451052 701244
rect 451052 701188 451056 701244
rect 450992 701184 451056 701188
rect 451072 701244 451136 701248
rect 451072 701188 451076 701244
rect 451076 701188 451132 701244
rect 451132 701188 451136 701244
rect 451072 701184 451136 701188
rect 451152 701244 451216 701248
rect 451152 701188 451156 701244
rect 451156 701188 451212 701244
rect 451212 701188 451216 701244
rect 451152 701184 451216 701188
rect 451232 701244 451296 701248
rect 451232 701188 451236 701244
rect 451236 701188 451292 701244
rect 451292 701188 451296 701244
rect 451232 701184 451296 701188
rect 451312 701244 451376 701248
rect 451312 701188 451316 701244
rect 451316 701188 451372 701244
rect 451372 701188 451376 701244
rect 451312 701184 451376 701188
rect 486832 701244 486896 701248
rect 486832 701188 486836 701244
rect 486836 701188 486892 701244
rect 486892 701188 486896 701244
rect 486832 701184 486896 701188
rect 486912 701244 486976 701248
rect 486912 701188 486916 701244
rect 486916 701188 486972 701244
rect 486972 701188 486976 701244
rect 486912 701184 486976 701188
rect 486992 701244 487056 701248
rect 486992 701188 486996 701244
rect 486996 701188 487052 701244
rect 487052 701188 487056 701244
rect 486992 701184 487056 701188
rect 487072 701244 487136 701248
rect 487072 701188 487076 701244
rect 487076 701188 487132 701244
rect 487132 701188 487136 701244
rect 487072 701184 487136 701188
rect 487152 701244 487216 701248
rect 487152 701188 487156 701244
rect 487156 701188 487212 701244
rect 487212 701188 487216 701244
rect 487152 701184 487216 701188
rect 487232 701244 487296 701248
rect 487232 701188 487236 701244
rect 487236 701188 487292 701244
rect 487292 701188 487296 701244
rect 487232 701184 487296 701188
rect 487312 701244 487376 701248
rect 487312 701188 487316 701244
rect 487316 701188 487372 701244
rect 487372 701188 487376 701244
rect 487312 701184 487376 701188
rect 522832 701244 522896 701248
rect 522832 701188 522836 701244
rect 522836 701188 522892 701244
rect 522892 701188 522896 701244
rect 522832 701184 522896 701188
rect 522912 701244 522976 701248
rect 522912 701188 522916 701244
rect 522916 701188 522972 701244
rect 522972 701188 522976 701244
rect 522912 701184 522976 701188
rect 522992 701244 523056 701248
rect 522992 701188 522996 701244
rect 522996 701188 523052 701244
rect 523052 701188 523056 701244
rect 522992 701184 523056 701188
rect 523072 701244 523136 701248
rect 523072 701188 523076 701244
rect 523076 701188 523132 701244
rect 523132 701188 523136 701244
rect 523072 701184 523136 701188
rect 523152 701244 523216 701248
rect 523152 701188 523156 701244
rect 523156 701188 523212 701244
rect 523212 701188 523216 701244
rect 523152 701184 523216 701188
rect 523232 701244 523296 701248
rect 523232 701188 523236 701244
rect 523236 701188 523292 701244
rect 523292 701188 523296 701244
rect 523232 701184 523296 701188
rect 523312 701244 523376 701248
rect 523312 701188 523316 701244
rect 523316 701188 523372 701244
rect 523372 701188 523376 701244
rect 523312 701184 523376 701188
rect 558832 701244 558896 701248
rect 558832 701188 558836 701244
rect 558836 701188 558892 701244
rect 558892 701188 558896 701244
rect 558832 701184 558896 701188
rect 558912 701244 558976 701248
rect 558912 701188 558916 701244
rect 558916 701188 558972 701244
rect 558972 701188 558976 701244
rect 558912 701184 558976 701188
rect 558992 701244 559056 701248
rect 558992 701188 558996 701244
rect 558996 701188 559052 701244
rect 559052 701188 559056 701244
rect 558992 701184 559056 701188
rect 559072 701244 559136 701248
rect 559072 701188 559076 701244
rect 559076 701188 559132 701244
rect 559132 701188 559136 701244
rect 559072 701184 559136 701188
rect 559152 701244 559216 701248
rect 559152 701188 559156 701244
rect 559156 701188 559212 701244
rect 559212 701188 559216 701244
rect 559152 701184 559216 701188
rect 559232 701244 559296 701248
rect 559232 701188 559236 701244
rect 559236 701188 559292 701244
rect 559292 701188 559296 701244
rect 559232 701184 559296 701188
rect 559312 701244 559376 701248
rect 559312 701188 559316 701244
rect 559316 701188 559372 701244
rect 559372 701188 559376 701244
rect 559312 701184 559376 701188
rect 36832 700700 36896 700704
rect 36832 700644 36836 700700
rect 36836 700644 36892 700700
rect 36892 700644 36896 700700
rect 36832 700640 36896 700644
rect 36912 700700 36976 700704
rect 36912 700644 36916 700700
rect 36916 700644 36972 700700
rect 36972 700644 36976 700700
rect 36912 700640 36976 700644
rect 36992 700700 37056 700704
rect 36992 700644 36996 700700
rect 36996 700644 37052 700700
rect 37052 700644 37056 700700
rect 36992 700640 37056 700644
rect 37072 700700 37136 700704
rect 37072 700644 37076 700700
rect 37076 700644 37132 700700
rect 37132 700644 37136 700700
rect 37072 700640 37136 700644
rect 37152 700700 37216 700704
rect 37152 700644 37156 700700
rect 37156 700644 37212 700700
rect 37212 700644 37216 700700
rect 37152 700640 37216 700644
rect 37232 700700 37296 700704
rect 37232 700644 37236 700700
rect 37236 700644 37292 700700
rect 37292 700644 37296 700700
rect 37232 700640 37296 700644
rect 37312 700700 37376 700704
rect 37312 700644 37316 700700
rect 37316 700644 37372 700700
rect 37372 700644 37376 700700
rect 37312 700640 37376 700644
rect 72832 700700 72896 700704
rect 72832 700644 72836 700700
rect 72836 700644 72892 700700
rect 72892 700644 72896 700700
rect 72832 700640 72896 700644
rect 72912 700700 72976 700704
rect 72912 700644 72916 700700
rect 72916 700644 72972 700700
rect 72972 700644 72976 700700
rect 72912 700640 72976 700644
rect 72992 700700 73056 700704
rect 72992 700644 72996 700700
rect 72996 700644 73052 700700
rect 73052 700644 73056 700700
rect 72992 700640 73056 700644
rect 73072 700700 73136 700704
rect 73072 700644 73076 700700
rect 73076 700644 73132 700700
rect 73132 700644 73136 700700
rect 73072 700640 73136 700644
rect 73152 700700 73216 700704
rect 73152 700644 73156 700700
rect 73156 700644 73212 700700
rect 73212 700644 73216 700700
rect 73152 700640 73216 700644
rect 73232 700700 73296 700704
rect 73232 700644 73236 700700
rect 73236 700644 73292 700700
rect 73292 700644 73296 700700
rect 73232 700640 73296 700644
rect 73312 700700 73376 700704
rect 73312 700644 73316 700700
rect 73316 700644 73372 700700
rect 73372 700644 73376 700700
rect 73312 700640 73376 700644
rect 108832 700700 108896 700704
rect 108832 700644 108836 700700
rect 108836 700644 108892 700700
rect 108892 700644 108896 700700
rect 108832 700640 108896 700644
rect 108912 700700 108976 700704
rect 108912 700644 108916 700700
rect 108916 700644 108972 700700
rect 108972 700644 108976 700700
rect 108912 700640 108976 700644
rect 108992 700700 109056 700704
rect 108992 700644 108996 700700
rect 108996 700644 109052 700700
rect 109052 700644 109056 700700
rect 108992 700640 109056 700644
rect 109072 700700 109136 700704
rect 109072 700644 109076 700700
rect 109076 700644 109132 700700
rect 109132 700644 109136 700700
rect 109072 700640 109136 700644
rect 109152 700700 109216 700704
rect 109152 700644 109156 700700
rect 109156 700644 109212 700700
rect 109212 700644 109216 700700
rect 109152 700640 109216 700644
rect 109232 700700 109296 700704
rect 109232 700644 109236 700700
rect 109236 700644 109292 700700
rect 109292 700644 109296 700700
rect 109232 700640 109296 700644
rect 109312 700700 109376 700704
rect 109312 700644 109316 700700
rect 109316 700644 109372 700700
rect 109372 700644 109376 700700
rect 109312 700640 109376 700644
rect 144832 700700 144896 700704
rect 144832 700644 144836 700700
rect 144836 700644 144892 700700
rect 144892 700644 144896 700700
rect 144832 700640 144896 700644
rect 144912 700700 144976 700704
rect 144912 700644 144916 700700
rect 144916 700644 144972 700700
rect 144972 700644 144976 700700
rect 144912 700640 144976 700644
rect 144992 700700 145056 700704
rect 144992 700644 144996 700700
rect 144996 700644 145052 700700
rect 145052 700644 145056 700700
rect 144992 700640 145056 700644
rect 145072 700700 145136 700704
rect 145072 700644 145076 700700
rect 145076 700644 145132 700700
rect 145132 700644 145136 700700
rect 145072 700640 145136 700644
rect 145152 700700 145216 700704
rect 145152 700644 145156 700700
rect 145156 700644 145212 700700
rect 145212 700644 145216 700700
rect 145152 700640 145216 700644
rect 145232 700700 145296 700704
rect 145232 700644 145236 700700
rect 145236 700644 145292 700700
rect 145292 700644 145296 700700
rect 145232 700640 145296 700644
rect 145312 700700 145376 700704
rect 145312 700644 145316 700700
rect 145316 700644 145372 700700
rect 145372 700644 145376 700700
rect 145312 700640 145376 700644
rect 180832 700700 180896 700704
rect 180832 700644 180836 700700
rect 180836 700644 180892 700700
rect 180892 700644 180896 700700
rect 180832 700640 180896 700644
rect 180912 700700 180976 700704
rect 180912 700644 180916 700700
rect 180916 700644 180972 700700
rect 180972 700644 180976 700700
rect 180912 700640 180976 700644
rect 180992 700700 181056 700704
rect 180992 700644 180996 700700
rect 180996 700644 181052 700700
rect 181052 700644 181056 700700
rect 180992 700640 181056 700644
rect 181072 700700 181136 700704
rect 181072 700644 181076 700700
rect 181076 700644 181132 700700
rect 181132 700644 181136 700700
rect 181072 700640 181136 700644
rect 181152 700700 181216 700704
rect 181152 700644 181156 700700
rect 181156 700644 181212 700700
rect 181212 700644 181216 700700
rect 181152 700640 181216 700644
rect 181232 700700 181296 700704
rect 181232 700644 181236 700700
rect 181236 700644 181292 700700
rect 181292 700644 181296 700700
rect 181232 700640 181296 700644
rect 181312 700700 181376 700704
rect 181312 700644 181316 700700
rect 181316 700644 181372 700700
rect 181372 700644 181376 700700
rect 181312 700640 181376 700644
rect 216832 700700 216896 700704
rect 216832 700644 216836 700700
rect 216836 700644 216892 700700
rect 216892 700644 216896 700700
rect 216832 700640 216896 700644
rect 216912 700700 216976 700704
rect 216912 700644 216916 700700
rect 216916 700644 216972 700700
rect 216972 700644 216976 700700
rect 216912 700640 216976 700644
rect 216992 700700 217056 700704
rect 216992 700644 216996 700700
rect 216996 700644 217052 700700
rect 217052 700644 217056 700700
rect 216992 700640 217056 700644
rect 217072 700700 217136 700704
rect 217072 700644 217076 700700
rect 217076 700644 217132 700700
rect 217132 700644 217136 700700
rect 217072 700640 217136 700644
rect 217152 700700 217216 700704
rect 217152 700644 217156 700700
rect 217156 700644 217212 700700
rect 217212 700644 217216 700700
rect 217152 700640 217216 700644
rect 217232 700700 217296 700704
rect 217232 700644 217236 700700
rect 217236 700644 217292 700700
rect 217292 700644 217296 700700
rect 217232 700640 217296 700644
rect 217312 700700 217376 700704
rect 217312 700644 217316 700700
rect 217316 700644 217372 700700
rect 217372 700644 217376 700700
rect 217312 700640 217376 700644
rect 252832 700700 252896 700704
rect 252832 700644 252836 700700
rect 252836 700644 252892 700700
rect 252892 700644 252896 700700
rect 252832 700640 252896 700644
rect 252912 700700 252976 700704
rect 252912 700644 252916 700700
rect 252916 700644 252972 700700
rect 252972 700644 252976 700700
rect 252912 700640 252976 700644
rect 252992 700700 253056 700704
rect 252992 700644 252996 700700
rect 252996 700644 253052 700700
rect 253052 700644 253056 700700
rect 252992 700640 253056 700644
rect 253072 700700 253136 700704
rect 253072 700644 253076 700700
rect 253076 700644 253132 700700
rect 253132 700644 253136 700700
rect 253072 700640 253136 700644
rect 253152 700700 253216 700704
rect 253152 700644 253156 700700
rect 253156 700644 253212 700700
rect 253212 700644 253216 700700
rect 253152 700640 253216 700644
rect 253232 700700 253296 700704
rect 253232 700644 253236 700700
rect 253236 700644 253292 700700
rect 253292 700644 253296 700700
rect 253232 700640 253296 700644
rect 253312 700700 253376 700704
rect 253312 700644 253316 700700
rect 253316 700644 253372 700700
rect 253372 700644 253376 700700
rect 253312 700640 253376 700644
rect 288832 700700 288896 700704
rect 288832 700644 288836 700700
rect 288836 700644 288892 700700
rect 288892 700644 288896 700700
rect 288832 700640 288896 700644
rect 288912 700700 288976 700704
rect 288912 700644 288916 700700
rect 288916 700644 288972 700700
rect 288972 700644 288976 700700
rect 288912 700640 288976 700644
rect 288992 700700 289056 700704
rect 288992 700644 288996 700700
rect 288996 700644 289052 700700
rect 289052 700644 289056 700700
rect 288992 700640 289056 700644
rect 289072 700700 289136 700704
rect 289072 700644 289076 700700
rect 289076 700644 289132 700700
rect 289132 700644 289136 700700
rect 289072 700640 289136 700644
rect 289152 700700 289216 700704
rect 289152 700644 289156 700700
rect 289156 700644 289212 700700
rect 289212 700644 289216 700700
rect 289152 700640 289216 700644
rect 289232 700700 289296 700704
rect 289232 700644 289236 700700
rect 289236 700644 289292 700700
rect 289292 700644 289296 700700
rect 289232 700640 289296 700644
rect 289312 700700 289376 700704
rect 289312 700644 289316 700700
rect 289316 700644 289372 700700
rect 289372 700644 289376 700700
rect 289312 700640 289376 700644
rect 324832 700700 324896 700704
rect 324832 700644 324836 700700
rect 324836 700644 324892 700700
rect 324892 700644 324896 700700
rect 324832 700640 324896 700644
rect 324912 700700 324976 700704
rect 324912 700644 324916 700700
rect 324916 700644 324972 700700
rect 324972 700644 324976 700700
rect 324912 700640 324976 700644
rect 324992 700700 325056 700704
rect 324992 700644 324996 700700
rect 324996 700644 325052 700700
rect 325052 700644 325056 700700
rect 324992 700640 325056 700644
rect 325072 700700 325136 700704
rect 325072 700644 325076 700700
rect 325076 700644 325132 700700
rect 325132 700644 325136 700700
rect 325072 700640 325136 700644
rect 325152 700700 325216 700704
rect 325152 700644 325156 700700
rect 325156 700644 325212 700700
rect 325212 700644 325216 700700
rect 325152 700640 325216 700644
rect 325232 700700 325296 700704
rect 325232 700644 325236 700700
rect 325236 700644 325292 700700
rect 325292 700644 325296 700700
rect 325232 700640 325296 700644
rect 325312 700700 325376 700704
rect 325312 700644 325316 700700
rect 325316 700644 325372 700700
rect 325372 700644 325376 700700
rect 325312 700640 325376 700644
rect 360832 700700 360896 700704
rect 360832 700644 360836 700700
rect 360836 700644 360892 700700
rect 360892 700644 360896 700700
rect 360832 700640 360896 700644
rect 360912 700700 360976 700704
rect 360912 700644 360916 700700
rect 360916 700644 360972 700700
rect 360972 700644 360976 700700
rect 360912 700640 360976 700644
rect 360992 700700 361056 700704
rect 360992 700644 360996 700700
rect 360996 700644 361052 700700
rect 361052 700644 361056 700700
rect 360992 700640 361056 700644
rect 361072 700700 361136 700704
rect 361072 700644 361076 700700
rect 361076 700644 361132 700700
rect 361132 700644 361136 700700
rect 361072 700640 361136 700644
rect 361152 700700 361216 700704
rect 361152 700644 361156 700700
rect 361156 700644 361212 700700
rect 361212 700644 361216 700700
rect 361152 700640 361216 700644
rect 361232 700700 361296 700704
rect 361232 700644 361236 700700
rect 361236 700644 361292 700700
rect 361292 700644 361296 700700
rect 361232 700640 361296 700644
rect 361312 700700 361376 700704
rect 361312 700644 361316 700700
rect 361316 700644 361372 700700
rect 361372 700644 361376 700700
rect 361312 700640 361376 700644
rect 396832 700700 396896 700704
rect 396832 700644 396836 700700
rect 396836 700644 396892 700700
rect 396892 700644 396896 700700
rect 396832 700640 396896 700644
rect 396912 700700 396976 700704
rect 396912 700644 396916 700700
rect 396916 700644 396972 700700
rect 396972 700644 396976 700700
rect 396912 700640 396976 700644
rect 396992 700700 397056 700704
rect 396992 700644 396996 700700
rect 396996 700644 397052 700700
rect 397052 700644 397056 700700
rect 396992 700640 397056 700644
rect 397072 700700 397136 700704
rect 397072 700644 397076 700700
rect 397076 700644 397132 700700
rect 397132 700644 397136 700700
rect 397072 700640 397136 700644
rect 397152 700700 397216 700704
rect 397152 700644 397156 700700
rect 397156 700644 397212 700700
rect 397212 700644 397216 700700
rect 397152 700640 397216 700644
rect 397232 700700 397296 700704
rect 397232 700644 397236 700700
rect 397236 700644 397292 700700
rect 397292 700644 397296 700700
rect 397232 700640 397296 700644
rect 397312 700700 397376 700704
rect 397312 700644 397316 700700
rect 397316 700644 397372 700700
rect 397372 700644 397376 700700
rect 397312 700640 397376 700644
rect 432832 700700 432896 700704
rect 432832 700644 432836 700700
rect 432836 700644 432892 700700
rect 432892 700644 432896 700700
rect 432832 700640 432896 700644
rect 432912 700700 432976 700704
rect 432912 700644 432916 700700
rect 432916 700644 432972 700700
rect 432972 700644 432976 700700
rect 432912 700640 432976 700644
rect 432992 700700 433056 700704
rect 432992 700644 432996 700700
rect 432996 700644 433052 700700
rect 433052 700644 433056 700700
rect 432992 700640 433056 700644
rect 433072 700700 433136 700704
rect 433072 700644 433076 700700
rect 433076 700644 433132 700700
rect 433132 700644 433136 700700
rect 433072 700640 433136 700644
rect 433152 700700 433216 700704
rect 433152 700644 433156 700700
rect 433156 700644 433212 700700
rect 433212 700644 433216 700700
rect 433152 700640 433216 700644
rect 433232 700700 433296 700704
rect 433232 700644 433236 700700
rect 433236 700644 433292 700700
rect 433292 700644 433296 700700
rect 433232 700640 433296 700644
rect 433312 700700 433376 700704
rect 433312 700644 433316 700700
rect 433316 700644 433372 700700
rect 433372 700644 433376 700700
rect 433312 700640 433376 700644
rect 468832 700700 468896 700704
rect 468832 700644 468836 700700
rect 468836 700644 468892 700700
rect 468892 700644 468896 700700
rect 468832 700640 468896 700644
rect 468912 700700 468976 700704
rect 468912 700644 468916 700700
rect 468916 700644 468972 700700
rect 468972 700644 468976 700700
rect 468912 700640 468976 700644
rect 468992 700700 469056 700704
rect 468992 700644 468996 700700
rect 468996 700644 469052 700700
rect 469052 700644 469056 700700
rect 468992 700640 469056 700644
rect 469072 700700 469136 700704
rect 469072 700644 469076 700700
rect 469076 700644 469132 700700
rect 469132 700644 469136 700700
rect 469072 700640 469136 700644
rect 469152 700700 469216 700704
rect 469152 700644 469156 700700
rect 469156 700644 469212 700700
rect 469212 700644 469216 700700
rect 469152 700640 469216 700644
rect 469232 700700 469296 700704
rect 469232 700644 469236 700700
rect 469236 700644 469292 700700
rect 469292 700644 469296 700700
rect 469232 700640 469296 700644
rect 469312 700700 469376 700704
rect 469312 700644 469316 700700
rect 469316 700644 469372 700700
rect 469372 700644 469376 700700
rect 469312 700640 469376 700644
rect 504832 700700 504896 700704
rect 504832 700644 504836 700700
rect 504836 700644 504892 700700
rect 504892 700644 504896 700700
rect 504832 700640 504896 700644
rect 504912 700700 504976 700704
rect 504912 700644 504916 700700
rect 504916 700644 504972 700700
rect 504972 700644 504976 700700
rect 504912 700640 504976 700644
rect 504992 700700 505056 700704
rect 504992 700644 504996 700700
rect 504996 700644 505052 700700
rect 505052 700644 505056 700700
rect 504992 700640 505056 700644
rect 505072 700700 505136 700704
rect 505072 700644 505076 700700
rect 505076 700644 505132 700700
rect 505132 700644 505136 700700
rect 505072 700640 505136 700644
rect 505152 700700 505216 700704
rect 505152 700644 505156 700700
rect 505156 700644 505212 700700
rect 505212 700644 505216 700700
rect 505152 700640 505216 700644
rect 505232 700700 505296 700704
rect 505232 700644 505236 700700
rect 505236 700644 505292 700700
rect 505292 700644 505296 700700
rect 505232 700640 505296 700644
rect 505312 700700 505376 700704
rect 505312 700644 505316 700700
rect 505316 700644 505372 700700
rect 505372 700644 505376 700700
rect 505312 700640 505376 700644
rect 540832 700700 540896 700704
rect 540832 700644 540836 700700
rect 540836 700644 540892 700700
rect 540892 700644 540896 700700
rect 540832 700640 540896 700644
rect 540912 700700 540976 700704
rect 540912 700644 540916 700700
rect 540916 700644 540972 700700
rect 540972 700644 540976 700700
rect 540912 700640 540976 700644
rect 540992 700700 541056 700704
rect 540992 700644 540996 700700
rect 540996 700644 541052 700700
rect 541052 700644 541056 700700
rect 540992 700640 541056 700644
rect 541072 700700 541136 700704
rect 541072 700644 541076 700700
rect 541076 700644 541132 700700
rect 541132 700644 541136 700700
rect 541072 700640 541136 700644
rect 541152 700700 541216 700704
rect 541152 700644 541156 700700
rect 541156 700644 541212 700700
rect 541212 700644 541216 700700
rect 541152 700640 541216 700644
rect 541232 700700 541296 700704
rect 541232 700644 541236 700700
rect 541236 700644 541292 700700
rect 541292 700644 541296 700700
rect 541232 700640 541296 700644
rect 541312 700700 541376 700704
rect 541312 700644 541316 700700
rect 541316 700644 541372 700700
rect 541372 700644 541376 700700
rect 541312 700640 541376 700644
rect 576832 700700 576896 700704
rect 576832 700644 576836 700700
rect 576836 700644 576892 700700
rect 576892 700644 576896 700700
rect 576832 700640 576896 700644
rect 576912 700700 576976 700704
rect 576912 700644 576916 700700
rect 576916 700644 576972 700700
rect 576972 700644 576976 700700
rect 576912 700640 576976 700644
rect 576992 700700 577056 700704
rect 576992 700644 576996 700700
rect 576996 700644 577052 700700
rect 577052 700644 577056 700700
rect 576992 700640 577056 700644
rect 577072 700700 577136 700704
rect 577072 700644 577076 700700
rect 577076 700644 577132 700700
rect 577132 700644 577136 700700
rect 577072 700640 577136 700644
rect 577152 700700 577216 700704
rect 577152 700644 577156 700700
rect 577156 700644 577212 700700
rect 577212 700644 577216 700700
rect 577152 700640 577216 700644
rect 577232 700700 577296 700704
rect 577232 700644 577236 700700
rect 577236 700644 577292 700700
rect 577292 700644 577296 700700
rect 577232 700640 577296 700644
rect 577312 700700 577376 700704
rect 577312 700644 577316 700700
rect 577316 700644 577372 700700
rect 577372 700644 577376 700700
rect 577312 700640 577376 700644
rect 18832 700156 18896 700160
rect 18832 700100 18836 700156
rect 18836 700100 18892 700156
rect 18892 700100 18896 700156
rect 18832 700096 18896 700100
rect 18912 700156 18976 700160
rect 18912 700100 18916 700156
rect 18916 700100 18972 700156
rect 18972 700100 18976 700156
rect 18912 700096 18976 700100
rect 18992 700156 19056 700160
rect 18992 700100 18996 700156
rect 18996 700100 19052 700156
rect 19052 700100 19056 700156
rect 18992 700096 19056 700100
rect 19072 700156 19136 700160
rect 19072 700100 19076 700156
rect 19076 700100 19132 700156
rect 19132 700100 19136 700156
rect 19072 700096 19136 700100
rect 19152 700156 19216 700160
rect 19152 700100 19156 700156
rect 19156 700100 19212 700156
rect 19212 700100 19216 700156
rect 19152 700096 19216 700100
rect 19232 700156 19296 700160
rect 19232 700100 19236 700156
rect 19236 700100 19292 700156
rect 19292 700100 19296 700156
rect 19232 700096 19296 700100
rect 19312 700156 19376 700160
rect 19312 700100 19316 700156
rect 19316 700100 19372 700156
rect 19372 700100 19376 700156
rect 19312 700096 19376 700100
rect 54832 700156 54896 700160
rect 54832 700100 54836 700156
rect 54836 700100 54892 700156
rect 54892 700100 54896 700156
rect 54832 700096 54896 700100
rect 54912 700156 54976 700160
rect 54912 700100 54916 700156
rect 54916 700100 54972 700156
rect 54972 700100 54976 700156
rect 54912 700096 54976 700100
rect 54992 700156 55056 700160
rect 54992 700100 54996 700156
rect 54996 700100 55052 700156
rect 55052 700100 55056 700156
rect 54992 700096 55056 700100
rect 55072 700156 55136 700160
rect 55072 700100 55076 700156
rect 55076 700100 55132 700156
rect 55132 700100 55136 700156
rect 55072 700096 55136 700100
rect 55152 700156 55216 700160
rect 55152 700100 55156 700156
rect 55156 700100 55212 700156
rect 55212 700100 55216 700156
rect 55152 700096 55216 700100
rect 55232 700156 55296 700160
rect 55232 700100 55236 700156
rect 55236 700100 55292 700156
rect 55292 700100 55296 700156
rect 55232 700096 55296 700100
rect 55312 700156 55376 700160
rect 55312 700100 55316 700156
rect 55316 700100 55372 700156
rect 55372 700100 55376 700156
rect 55312 700096 55376 700100
rect 90832 700156 90896 700160
rect 90832 700100 90836 700156
rect 90836 700100 90892 700156
rect 90892 700100 90896 700156
rect 90832 700096 90896 700100
rect 90912 700156 90976 700160
rect 90912 700100 90916 700156
rect 90916 700100 90972 700156
rect 90972 700100 90976 700156
rect 90912 700096 90976 700100
rect 90992 700156 91056 700160
rect 90992 700100 90996 700156
rect 90996 700100 91052 700156
rect 91052 700100 91056 700156
rect 90992 700096 91056 700100
rect 91072 700156 91136 700160
rect 91072 700100 91076 700156
rect 91076 700100 91132 700156
rect 91132 700100 91136 700156
rect 91072 700096 91136 700100
rect 91152 700156 91216 700160
rect 91152 700100 91156 700156
rect 91156 700100 91212 700156
rect 91212 700100 91216 700156
rect 91152 700096 91216 700100
rect 91232 700156 91296 700160
rect 91232 700100 91236 700156
rect 91236 700100 91292 700156
rect 91292 700100 91296 700156
rect 91232 700096 91296 700100
rect 91312 700156 91376 700160
rect 91312 700100 91316 700156
rect 91316 700100 91372 700156
rect 91372 700100 91376 700156
rect 91312 700096 91376 700100
rect 126832 700156 126896 700160
rect 126832 700100 126836 700156
rect 126836 700100 126892 700156
rect 126892 700100 126896 700156
rect 126832 700096 126896 700100
rect 126912 700156 126976 700160
rect 126912 700100 126916 700156
rect 126916 700100 126972 700156
rect 126972 700100 126976 700156
rect 126912 700096 126976 700100
rect 126992 700156 127056 700160
rect 126992 700100 126996 700156
rect 126996 700100 127052 700156
rect 127052 700100 127056 700156
rect 126992 700096 127056 700100
rect 127072 700156 127136 700160
rect 127072 700100 127076 700156
rect 127076 700100 127132 700156
rect 127132 700100 127136 700156
rect 127072 700096 127136 700100
rect 127152 700156 127216 700160
rect 127152 700100 127156 700156
rect 127156 700100 127212 700156
rect 127212 700100 127216 700156
rect 127152 700096 127216 700100
rect 127232 700156 127296 700160
rect 127232 700100 127236 700156
rect 127236 700100 127292 700156
rect 127292 700100 127296 700156
rect 127232 700096 127296 700100
rect 127312 700156 127376 700160
rect 127312 700100 127316 700156
rect 127316 700100 127372 700156
rect 127372 700100 127376 700156
rect 127312 700096 127376 700100
rect 162832 700156 162896 700160
rect 162832 700100 162836 700156
rect 162836 700100 162892 700156
rect 162892 700100 162896 700156
rect 162832 700096 162896 700100
rect 162912 700156 162976 700160
rect 162912 700100 162916 700156
rect 162916 700100 162972 700156
rect 162972 700100 162976 700156
rect 162912 700096 162976 700100
rect 162992 700156 163056 700160
rect 162992 700100 162996 700156
rect 162996 700100 163052 700156
rect 163052 700100 163056 700156
rect 162992 700096 163056 700100
rect 163072 700156 163136 700160
rect 163072 700100 163076 700156
rect 163076 700100 163132 700156
rect 163132 700100 163136 700156
rect 163072 700096 163136 700100
rect 163152 700156 163216 700160
rect 163152 700100 163156 700156
rect 163156 700100 163212 700156
rect 163212 700100 163216 700156
rect 163152 700096 163216 700100
rect 163232 700156 163296 700160
rect 163232 700100 163236 700156
rect 163236 700100 163292 700156
rect 163292 700100 163296 700156
rect 163232 700096 163296 700100
rect 163312 700156 163376 700160
rect 163312 700100 163316 700156
rect 163316 700100 163372 700156
rect 163372 700100 163376 700156
rect 163312 700096 163376 700100
rect 198832 700156 198896 700160
rect 198832 700100 198836 700156
rect 198836 700100 198892 700156
rect 198892 700100 198896 700156
rect 198832 700096 198896 700100
rect 198912 700156 198976 700160
rect 198912 700100 198916 700156
rect 198916 700100 198972 700156
rect 198972 700100 198976 700156
rect 198912 700096 198976 700100
rect 198992 700156 199056 700160
rect 198992 700100 198996 700156
rect 198996 700100 199052 700156
rect 199052 700100 199056 700156
rect 198992 700096 199056 700100
rect 199072 700156 199136 700160
rect 199072 700100 199076 700156
rect 199076 700100 199132 700156
rect 199132 700100 199136 700156
rect 199072 700096 199136 700100
rect 199152 700156 199216 700160
rect 199152 700100 199156 700156
rect 199156 700100 199212 700156
rect 199212 700100 199216 700156
rect 199152 700096 199216 700100
rect 199232 700156 199296 700160
rect 199232 700100 199236 700156
rect 199236 700100 199292 700156
rect 199292 700100 199296 700156
rect 199232 700096 199296 700100
rect 199312 700156 199376 700160
rect 199312 700100 199316 700156
rect 199316 700100 199372 700156
rect 199372 700100 199376 700156
rect 199312 700096 199376 700100
rect 234832 700156 234896 700160
rect 234832 700100 234836 700156
rect 234836 700100 234892 700156
rect 234892 700100 234896 700156
rect 234832 700096 234896 700100
rect 234912 700156 234976 700160
rect 234912 700100 234916 700156
rect 234916 700100 234972 700156
rect 234972 700100 234976 700156
rect 234912 700096 234976 700100
rect 234992 700156 235056 700160
rect 234992 700100 234996 700156
rect 234996 700100 235052 700156
rect 235052 700100 235056 700156
rect 234992 700096 235056 700100
rect 235072 700156 235136 700160
rect 235072 700100 235076 700156
rect 235076 700100 235132 700156
rect 235132 700100 235136 700156
rect 235072 700096 235136 700100
rect 235152 700156 235216 700160
rect 235152 700100 235156 700156
rect 235156 700100 235212 700156
rect 235212 700100 235216 700156
rect 235152 700096 235216 700100
rect 235232 700156 235296 700160
rect 235232 700100 235236 700156
rect 235236 700100 235292 700156
rect 235292 700100 235296 700156
rect 235232 700096 235296 700100
rect 235312 700156 235376 700160
rect 235312 700100 235316 700156
rect 235316 700100 235372 700156
rect 235372 700100 235376 700156
rect 235312 700096 235376 700100
rect 270832 700156 270896 700160
rect 270832 700100 270836 700156
rect 270836 700100 270892 700156
rect 270892 700100 270896 700156
rect 270832 700096 270896 700100
rect 270912 700156 270976 700160
rect 270912 700100 270916 700156
rect 270916 700100 270972 700156
rect 270972 700100 270976 700156
rect 270912 700096 270976 700100
rect 270992 700156 271056 700160
rect 270992 700100 270996 700156
rect 270996 700100 271052 700156
rect 271052 700100 271056 700156
rect 270992 700096 271056 700100
rect 271072 700156 271136 700160
rect 271072 700100 271076 700156
rect 271076 700100 271132 700156
rect 271132 700100 271136 700156
rect 271072 700096 271136 700100
rect 271152 700156 271216 700160
rect 271152 700100 271156 700156
rect 271156 700100 271212 700156
rect 271212 700100 271216 700156
rect 271152 700096 271216 700100
rect 271232 700156 271296 700160
rect 271232 700100 271236 700156
rect 271236 700100 271292 700156
rect 271292 700100 271296 700156
rect 271232 700096 271296 700100
rect 271312 700156 271376 700160
rect 271312 700100 271316 700156
rect 271316 700100 271372 700156
rect 271372 700100 271376 700156
rect 271312 700096 271376 700100
rect 306832 700156 306896 700160
rect 306832 700100 306836 700156
rect 306836 700100 306892 700156
rect 306892 700100 306896 700156
rect 306832 700096 306896 700100
rect 306912 700156 306976 700160
rect 306912 700100 306916 700156
rect 306916 700100 306972 700156
rect 306972 700100 306976 700156
rect 306912 700096 306976 700100
rect 306992 700156 307056 700160
rect 306992 700100 306996 700156
rect 306996 700100 307052 700156
rect 307052 700100 307056 700156
rect 306992 700096 307056 700100
rect 307072 700156 307136 700160
rect 307072 700100 307076 700156
rect 307076 700100 307132 700156
rect 307132 700100 307136 700156
rect 307072 700096 307136 700100
rect 307152 700156 307216 700160
rect 307152 700100 307156 700156
rect 307156 700100 307212 700156
rect 307212 700100 307216 700156
rect 307152 700096 307216 700100
rect 307232 700156 307296 700160
rect 307232 700100 307236 700156
rect 307236 700100 307292 700156
rect 307292 700100 307296 700156
rect 307232 700096 307296 700100
rect 307312 700156 307376 700160
rect 307312 700100 307316 700156
rect 307316 700100 307372 700156
rect 307372 700100 307376 700156
rect 307312 700096 307376 700100
rect 342832 700156 342896 700160
rect 342832 700100 342836 700156
rect 342836 700100 342892 700156
rect 342892 700100 342896 700156
rect 342832 700096 342896 700100
rect 342912 700156 342976 700160
rect 342912 700100 342916 700156
rect 342916 700100 342972 700156
rect 342972 700100 342976 700156
rect 342912 700096 342976 700100
rect 342992 700156 343056 700160
rect 342992 700100 342996 700156
rect 342996 700100 343052 700156
rect 343052 700100 343056 700156
rect 342992 700096 343056 700100
rect 343072 700156 343136 700160
rect 343072 700100 343076 700156
rect 343076 700100 343132 700156
rect 343132 700100 343136 700156
rect 343072 700096 343136 700100
rect 343152 700156 343216 700160
rect 343152 700100 343156 700156
rect 343156 700100 343212 700156
rect 343212 700100 343216 700156
rect 343152 700096 343216 700100
rect 343232 700156 343296 700160
rect 343232 700100 343236 700156
rect 343236 700100 343292 700156
rect 343292 700100 343296 700156
rect 343232 700096 343296 700100
rect 343312 700156 343376 700160
rect 343312 700100 343316 700156
rect 343316 700100 343372 700156
rect 343372 700100 343376 700156
rect 343312 700096 343376 700100
rect 378832 700156 378896 700160
rect 378832 700100 378836 700156
rect 378836 700100 378892 700156
rect 378892 700100 378896 700156
rect 378832 700096 378896 700100
rect 378912 700156 378976 700160
rect 378912 700100 378916 700156
rect 378916 700100 378972 700156
rect 378972 700100 378976 700156
rect 378912 700096 378976 700100
rect 378992 700156 379056 700160
rect 378992 700100 378996 700156
rect 378996 700100 379052 700156
rect 379052 700100 379056 700156
rect 378992 700096 379056 700100
rect 379072 700156 379136 700160
rect 379072 700100 379076 700156
rect 379076 700100 379132 700156
rect 379132 700100 379136 700156
rect 379072 700096 379136 700100
rect 379152 700156 379216 700160
rect 379152 700100 379156 700156
rect 379156 700100 379212 700156
rect 379212 700100 379216 700156
rect 379152 700096 379216 700100
rect 379232 700156 379296 700160
rect 379232 700100 379236 700156
rect 379236 700100 379292 700156
rect 379292 700100 379296 700156
rect 379232 700096 379296 700100
rect 379312 700156 379376 700160
rect 379312 700100 379316 700156
rect 379316 700100 379372 700156
rect 379372 700100 379376 700156
rect 379312 700096 379376 700100
rect 414832 700156 414896 700160
rect 414832 700100 414836 700156
rect 414836 700100 414892 700156
rect 414892 700100 414896 700156
rect 414832 700096 414896 700100
rect 414912 700156 414976 700160
rect 414912 700100 414916 700156
rect 414916 700100 414972 700156
rect 414972 700100 414976 700156
rect 414912 700096 414976 700100
rect 414992 700156 415056 700160
rect 414992 700100 414996 700156
rect 414996 700100 415052 700156
rect 415052 700100 415056 700156
rect 414992 700096 415056 700100
rect 415072 700156 415136 700160
rect 415072 700100 415076 700156
rect 415076 700100 415132 700156
rect 415132 700100 415136 700156
rect 415072 700096 415136 700100
rect 415152 700156 415216 700160
rect 415152 700100 415156 700156
rect 415156 700100 415212 700156
rect 415212 700100 415216 700156
rect 415152 700096 415216 700100
rect 415232 700156 415296 700160
rect 415232 700100 415236 700156
rect 415236 700100 415292 700156
rect 415292 700100 415296 700156
rect 415232 700096 415296 700100
rect 415312 700156 415376 700160
rect 415312 700100 415316 700156
rect 415316 700100 415372 700156
rect 415372 700100 415376 700156
rect 415312 700096 415376 700100
rect 450832 700156 450896 700160
rect 450832 700100 450836 700156
rect 450836 700100 450892 700156
rect 450892 700100 450896 700156
rect 450832 700096 450896 700100
rect 450912 700156 450976 700160
rect 450912 700100 450916 700156
rect 450916 700100 450972 700156
rect 450972 700100 450976 700156
rect 450912 700096 450976 700100
rect 450992 700156 451056 700160
rect 450992 700100 450996 700156
rect 450996 700100 451052 700156
rect 451052 700100 451056 700156
rect 450992 700096 451056 700100
rect 451072 700156 451136 700160
rect 451072 700100 451076 700156
rect 451076 700100 451132 700156
rect 451132 700100 451136 700156
rect 451072 700096 451136 700100
rect 451152 700156 451216 700160
rect 451152 700100 451156 700156
rect 451156 700100 451212 700156
rect 451212 700100 451216 700156
rect 451152 700096 451216 700100
rect 451232 700156 451296 700160
rect 451232 700100 451236 700156
rect 451236 700100 451292 700156
rect 451292 700100 451296 700156
rect 451232 700096 451296 700100
rect 451312 700156 451376 700160
rect 451312 700100 451316 700156
rect 451316 700100 451372 700156
rect 451372 700100 451376 700156
rect 451312 700096 451376 700100
rect 486832 700156 486896 700160
rect 486832 700100 486836 700156
rect 486836 700100 486892 700156
rect 486892 700100 486896 700156
rect 486832 700096 486896 700100
rect 486912 700156 486976 700160
rect 486912 700100 486916 700156
rect 486916 700100 486972 700156
rect 486972 700100 486976 700156
rect 486912 700096 486976 700100
rect 486992 700156 487056 700160
rect 486992 700100 486996 700156
rect 486996 700100 487052 700156
rect 487052 700100 487056 700156
rect 486992 700096 487056 700100
rect 487072 700156 487136 700160
rect 487072 700100 487076 700156
rect 487076 700100 487132 700156
rect 487132 700100 487136 700156
rect 487072 700096 487136 700100
rect 487152 700156 487216 700160
rect 487152 700100 487156 700156
rect 487156 700100 487212 700156
rect 487212 700100 487216 700156
rect 487152 700096 487216 700100
rect 487232 700156 487296 700160
rect 487232 700100 487236 700156
rect 487236 700100 487292 700156
rect 487292 700100 487296 700156
rect 487232 700096 487296 700100
rect 487312 700156 487376 700160
rect 487312 700100 487316 700156
rect 487316 700100 487372 700156
rect 487372 700100 487376 700156
rect 487312 700096 487376 700100
rect 522832 700156 522896 700160
rect 522832 700100 522836 700156
rect 522836 700100 522892 700156
rect 522892 700100 522896 700156
rect 522832 700096 522896 700100
rect 522912 700156 522976 700160
rect 522912 700100 522916 700156
rect 522916 700100 522972 700156
rect 522972 700100 522976 700156
rect 522912 700096 522976 700100
rect 522992 700156 523056 700160
rect 522992 700100 522996 700156
rect 522996 700100 523052 700156
rect 523052 700100 523056 700156
rect 522992 700096 523056 700100
rect 523072 700156 523136 700160
rect 523072 700100 523076 700156
rect 523076 700100 523132 700156
rect 523132 700100 523136 700156
rect 523072 700096 523136 700100
rect 523152 700156 523216 700160
rect 523152 700100 523156 700156
rect 523156 700100 523212 700156
rect 523212 700100 523216 700156
rect 523152 700096 523216 700100
rect 523232 700156 523296 700160
rect 523232 700100 523236 700156
rect 523236 700100 523292 700156
rect 523292 700100 523296 700156
rect 523232 700096 523296 700100
rect 523312 700156 523376 700160
rect 523312 700100 523316 700156
rect 523316 700100 523372 700156
rect 523372 700100 523376 700156
rect 523312 700096 523376 700100
rect 558832 700156 558896 700160
rect 558832 700100 558836 700156
rect 558836 700100 558892 700156
rect 558892 700100 558896 700156
rect 558832 700096 558896 700100
rect 558912 700156 558976 700160
rect 558912 700100 558916 700156
rect 558916 700100 558972 700156
rect 558972 700100 558976 700156
rect 558912 700096 558976 700100
rect 558992 700156 559056 700160
rect 558992 700100 558996 700156
rect 558996 700100 559052 700156
rect 559052 700100 559056 700156
rect 558992 700096 559056 700100
rect 559072 700156 559136 700160
rect 559072 700100 559076 700156
rect 559076 700100 559132 700156
rect 559132 700100 559136 700156
rect 559072 700096 559136 700100
rect 559152 700156 559216 700160
rect 559152 700100 559156 700156
rect 559156 700100 559212 700156
rect 559212 700100 559216 700156
rect 559152 700096 559216 700100
rect 559232 700156 559296 700160
rect 559232 700100 559236 700156
rect 559236 700100 559292 700156
rect 559292 700100 559296 700156
rect 559232 700096 559296 700100
rect 559312 700156 559376 700160
rect 559312 700100 559316 700156
rect 559316 700100 559372 700156
rect 559372 700100 559376 700156
rect 559312 700096 559376 700100
rect 36832 699612 36896 699616
rect 36832 699556 36836 699612
rect 36836 699556 36892 699612
rect 36892 699556 36896 699612
rect 36832 699552 36896 699556
rect 36912 699612 36976 699616
rect 36912 699556 36916 699612
rect 36916 699556 36972 699612
rect 36972 699556 36976 699612
rect 36912 699552 36976 699556
rect 36992 699612 37056 699616
rect 36992 699556 36996 699612
rect 36996 699556 37052 699612
rect 37052 699556 37056 699612
rect 36992 699552 37056 699556
rect 37072 699612 37136 699616
rect 37072 699556 37076 699612
rect 37076 699556 37132 699612
rect 37132 699556 37136 699612
rect 37072 699552 37136 699556
rect 37152 699612 37216 699616
rect 37152 699556 37156 699612
rect 37156 699556 37212 699612
rect 37212 699556 37216 699612
rect 37152 699552 37216 699556
rect 37232 699612 37296 699616
rect 37232 699556 37236 699612
rect 37236 699556 37292 699612
rect 37292 699556 37296 699612
rect 37232 699552 37296 699556
rect 37312 699612 37376 699616
rect 37312 699556 37316 699612
rect 37316 699556 37372 699612
rect 37372 699556 37376 699612
rect 37312 699552 37376 699556
rect 72832 699612 72896 699616
rect 72832 699556 72836 699612
rect 72836 699556 72892 699612
rect 72892 699556 72896 699612
rect 72832 699552 72896 699556
rect 72912 699612 72976 699616
rect 72912 699556 72916 699612
rect 72916 699556 72972 699612
rect 72972 699556 72976 699612
rect 72912 699552 72976 699556
rect 72992 699612 73056 699616
rect 72992 699556 72996 699612
rect 72996 699556 73052 699612
rect 73052 699556 73056 699612
rect 72992 699552 73056 699556
rect 73072 699612 73136 699616
rect 73072 699556 73076 699612
rect 73076 699556 73132 699612
rect 73132 699556 73136 699612
rect 73072 699552 73136 699556
rect 73152 699612 73216 699616
rect 73152 699556 73156 699612
rect 73156 699556 73212 699612
rect 73212 699556 73216 699612
rect 73152 699552 73216 699556
rect 73232 699612 73296 699616
rect 73232 699556 73236 699612
rect 73236 699556 73292 699612
rect 73292 699556 73296 699612
rect 73232 699552 73296 699556
rect 73312 699612 73376 699616
rect 73312 699556 73316 699612
rect 73316 699556 73372 699612
rect 73372 699556 73376 699612
rect 73312 699552 73376 699556
rect 108832 699612 108896 699616
rect 108832 699556 108836 699612
rect 108836 699556 108892 699612
rect 108892 699556 108896 699612
rect 108832 699552 108896 699556
rect 108912 699612 108976 699616
rect 108912 699556 108916 699612
rect 108916 699556 108972 699612
rect 108972 699556 108976 699612
rect 108912 699552 108976 699556
rect 108992 699612 109056 699616
rect 108992 699556 108996 699612
rect 108996 699556 109052 699612
rect 109052 699556 109056 699612
rect 108992 699552 109056 699556
rect 109072 699612 109136 699616
rect 109072 699556 109076 699612
rect 109076 699556 109132 699612
rect 109132 699556 109136 699612
rect 109072 699552 109136 699556
rect 109152 699612 109216 699616
rect 109152 699556 109156 699612
rect 109156 699556 109212 699612
rect 109212 699556 109216 699612
rect 109152 699552 109216 699556
rect 109232 699612 109296 699616
rect 109232 699556 109236 699612
rect 109236 699556 109292 699612
rect 109292 699556 109296 699612
rect 109232 699552 109296 699556
rect 109312 699612 109376 699616
rect 109312 699556 109316 699612
rect 109316 699556 109372 699612
rect 109372 699556 109376 699612
rect 109312 699552 109376 699556
rect 144832 699612 144896 699616
rect 144832 699556 144836 699612
rect 144836 699556 144892 699612
rect 144892 699556 144896 699612
rect 144832 699552 144896 699556
rect 144912 699612 144976 699616
rect 144912 699556 144916 699612
rect 144916 699556 144972 699612
rect 144972 699556 144976 699612
rect 144912 699552 144976 699556
rect 144992 699612 145056 699616
rect 144992 699556 144996 699612
rect 144996 699556 145052 699612
rect 145052 699556 145056 699612
rect 144992 699552 145056 699556
rect 145072 699612 145136 699616
rect 145072 699556 145076 699612
rect 145076 699556 145132 699612
rect 145132 699556 145136 699612
rect 145072 699552 145136 699556
rect 145152 699612 145216 699616
rect 145152 699556 145156 699612
rect 145156 699556 145212 699612
rect 145212 699556 145216 699612
rect 145152 699552 145216 699556
rect 145232 699612 145296 699616
rect 145232 699556 145236 699612
rect 145236 699556 145292 699612
rect 145292 699556 145296 699612
rect 145232 699552 145296 699556
rect 145312 699612 145376 699616
rect 145312 699556 145316 699612
rect 145316 699556 145372 699612
rect 145372 699556 145376 699612
rect 145312 699552 145376 699556
rect 180832 699612 180896 699616
rect 180832 699556 180836 699612
rect 180836 699556 180892 699612
rect 180892 699556 180896 699612
rect 180832 699552 180896 699556
rect 180912 699612 180976 699616
rect 180912 699556 180916 699612
rect 180916 699556 180972 699612
rect 180972 699556 180976 699612
rect 180912 699552 180976 699556
rect 180992 699612 181056 699616
rect 180992 699556 180996 699612
rect 180996 699556 181052 699612
rect 181052 699556 181056 699612
rect 180992 699552 181056 699556
rect 181072 699612 181136 699616
rect 181072 699556 181076 699612
rect 181076 699556 181132 699612
rect 181132 699556 181136 699612
rect 181072 699552 181136 699556
rect 181152 699612 181216 699616
rect 181152 699556 181156 699612
rect 181156 699556 181212 699612
rect 181212 699556 181216 699612
rect 181152 699552 181216 699556
rect 181232 699612 181296 699616
rect 181232 699556 181236 699612
rect 181236 699556 181292 699612
rect 181292 699556 181296 699612
rect 181232 699552 181296 699556
rect 181312 699612 181376 699616
rect 181312 699556 181316 699612
rect 181316 699556 181372 699612
rect 181372 699556 181376 699612
rect 181312 699552 181376 699556
rect 216832 699612 216896 699616
rect 216832 699556 216836 699612
rect 216836 699556 216892 699612
rect 216892 699556 216896 699612
rect 216832 699552 216896 699556
rect 216912 699612 216976 699616
rect 216912 699556 216916 699612
rect 216916 699556 216972 699612
rect 216972 699556 216976 699612
rect 216912 699552 216976 699556
rect 216992 699612 217056 699616
rect 216992 699556 216996 699612
rect 216996 699556 217052 699612
rect 217052 699556 217056 699612
rect 216992 699552 217056 699556
rect 217072 699612 217136 699616
rect 217072 699556 217076 699612
rect 217076 699556 217132 699612
rect 217132 699556 217136 699612
rect 217072 699552 217136 699556
rect 217152 699612 217216 699616
rect 217152 699556 217156 699612
rect 217156 699556 217212 699612
rect 217212 699556 217216 699612
rect 217152 699552 217216 699556
rect 217232 699612 217296 699616
rect 217232 699556 217236 699612
rect 217236 699556 217292 699612
rect 217292 699556 217296 699612
rect 217232 699552 217296 699556
rect 217312 699612 217376 699616
rect 217312 699556 217316 699612
rect 217316 699556 217372 699612
rect 217372 699556 217376 699612
rect 217312 699552 217376 699556
rect 252832 699612 252896 699616
rect 252832 699556 252836 699612
rect 252836 699556 252892 699612
rect 252892 699556 252896 699612
rect 252832 699552 252896 699556
rect 252912 699612 252976 699616
rect 252912 699556 252916 699612
rect 252916 699556 252972 699612
rect 252972 699556 252976 699612
rect 252912 699552 252976 699556
rect 252992 699612 253056 699616
rect 252992 699556 252996 699612
rect 252996 699556 253052 699612
rect 253052 699556 253056 699612
rect 252992 699552 253056 699556
rect 253072 699612 253136 699616
rect 253072 699556 253076 699612
rect 253076 699556 253132 699612
rect 253132 699556 253136 699612
rect 253072 699552 253136 699556
rect 253152 699612 253216 699616
rect 253152 699556 253156 699612
rect 253156 699556 253212 699612
rect 253212 699556 253216 699612
rect 253152 699552 253216 699556
rect 253232 699612 253296 699616
rect 253232 699556 253236 699612
rect 253236 699556 253292 699612
rect 253292 699556 253296 699612
rect 253232 699552 253296 699556
rect 253312 699612 253376 699616
rect 253312 699556 253316 699612
rect 253316 699556 253372 699612
rect 253372 699556 253376 699612
rect 253312 699552 253376 699556
rect 288832 699612 288896 699616
rect 288832 699556 288836 699612
rect 288836 699556 288892 699612
rect 288892 699556 288896 699612
rect 288832 699552 288896 699556
rect 288912 699612 288976 699616
rect 288912 699556 288916 699612
rect 288916 699556 288972 699612
rect 288972 699556 288976 699612
rect 288912 699552 288976 699556
rect 288992 699612 289056 699616
rect 288992 699556 288996 699612
rect 288996 699556 289052 699612
rect 289052 699556 289056 699612
rect 288992 699552 289056 699556
rect 289072 699612 289136 699616
rect 289072 699556 289076 699612
rect 289076 699556 289132 699612
rect 289132 699556 289136 699612
rect 289072 699552 289136 699556
rect 289152 699612 289216 699616
rect 289152 699556 289156 699612
rect 289156 699556 289212 699612
rect 289212 699556 289216 699612
rect 289152 699552 289216 699556
rect 289232 699612 289296 699616
rect 289232 699556 289236 699612
rect 289236 699556 289292 699612
rect 289292 699556 289296 699612
rect 289232 699552 289296 699556
rect 289312 699612 289376 699616
rect 289312 699556 289316 699612
rect 289316 699556 289372 699612
rect 289372 699556 289376 699612
rect 289312 699552 289376 699556
rect 324832 699612 324896 699616
rect 324832 699556 324836 699612
rect 324836 699556 324892 699612
rect 324892 699556 324896 699612
rect 324832 699552 324896 699556
rect 324912 699612 324976 699616
rect 324912 699556 324916 699612
rect 324916 699556 324972 699612
rect 324972 699556 324976 699612
rect 324912 699552 324976 699556
rect 324992 699612 325056 699616
rect 324992 699556 324996 699612
rect 324996 699556 325052 699612
rect 325052 699556 325056 699612
rect 324992 699552 325056 699556
rect 325072 699612 325136 699616
rect 325072 699556 325076 699612
rect 325076 699556 325132 699612
rect 325132 699556 325136 699612
rect 325072 699552 325136 699556
rect 325152 699612 325216 699616
rect 325152 699556 325156 699612
rect 325156 699556 325212 699612
rect 325212 699556 325216 699612
rect 325152 699552 325216 699556
rect 325232 699612 325296 699616
rect 325232 699556 325236 699612
rect 325236 699556 325292 699612
rect 325292 699556 325296 699612
rect 325232 699552 325296 699556
rect 325312 699612 325376 699616
rect 325312 699556 325316 699612
rect 325316 699556 325372 699612
rect 325372 699556 325376 699612
rect 325312 699552 325376 699556
rect 360832 699612 360896 699616
rect 360832 699556 360836 699612
rect 360836 699556 360892 699612
rect 360892 699556 360896 699612
rect 360832 699552 360896 699556
rect 360912 699612 360976 699616
rect 360912 699556 360916 699612
rect 360916 699556 360972 699612
rect 360972 699556 360976 699612
rect 360912 699552 360976 699556
rect 360992 699612 361056 699616
rect 360992 699556 360996 699612
rect 360996 699556 361052 699612
rect 361052 699556 361056 699612
rect 360992 699552 361056 699556
rect 361072 699612 361136 699616
rect 361072 699556 361076 699612
rect 361076 699556 361132 699612
rect 361132 699556 361136 699612
rect 361072 699552 361136 699556
rect 361152 699612 361216 699616
rect 361152 699556 361156 699612
rect 361156 699556 361212 699612
rect 361212 699556 361216 699612
rect 361152 699552 361216 699556
rect 361232 699612 361296 699616
rect 361232 699556 361236 699612
rect 361236 699556 361292 699612
rect 361292 699556 361296 699612
rect 361232 699552 361296 699556
rect 361312 699612 361376 699616
rect 361312 699556 361316 699612
rect 361316 699556 361372 699612
rect 361372 699556 361376 699612
rect 361312 699552 361376 699556
rect 396832 699612 396896 699616
rect 396832 699556 396836 699612
rect 396836 699556 396892 699612
rect 396892 699556 396896 699612
rect 396832 699552 396896 699556
rect 396912 699612 396976 699616
rect 396912 699556 396916 699612
rect 396916 699556 396972 699612
rect 396972 699556 396976 699612
rect 396912 699552 396976 699556
rect 396992 699612 397056 699616
rect 396992 699556 396996 699612
rect 396996 699556 397052 699612
rect 397052 699556 397056 699612
rect 396992 699552 397056 699556
rect 397072 699612 397136 699616
rect 397072 699556 397076 699612
rect 397076 699556 397132 699612
rect 397132 699556 397136 699612
rect 397072 699552 397136 699556
rect 397152 699612 397216 699616
rect 397152 699556 397156 699612
rect 397156 699556 397212 699612
rect 397212 699556 397216 699612
rect 397152 699552 397216 699556
rect 397232 699612 397296 699616
rect 397232 699556 397236 699612
rect 397236 699556 397292 699612
rect 397292 699556 397296 699612
rect 397232 699552 397296 699556
rect 397312 699612 397376 699616
rect 397312 699556 397316 699612
rect 397316 699556 397372 699612
rect 397372 699556 397376 699612
rect 397312 699552 397376 699556
rect 432832 699612 432896 699616
rect 432832 699556 432836 699612
rect 432836 699556 432892 699612
rect 432892 699556 432896 699612
rect 432832 699552 432896 699556
rect 432912 699612 432976 699616
rect 432912 699556 432916 699612
rect 432916 699556 432972 699612
rect 432972 699556 432976 699612
rect 432912 699552 432976 699556
rect 432992 699612 433056 699616
rect 432992 699556 432996 699612
rect 432996 699556 433052 699612
rect 433052 699556 433056 699612
rect 432992 699552 433056 699556
rect 433072 699612 433136 699616
rect 433072 699556 433076 699612
rect 433076 699556 433132 699612
rect 433132 699556 433136 699612
rect 433072 699552 433136 699556
rect 433152 699612 433216 699616
rect 433152 699556 433156 699612
rect 433156 699556 433212 699612
rect 433212 699556 433216 699612
rect 433152 699552 433216 699556
rect 433232 699612 433296 699616
rect 433232 699556 433236 699612
rect 433236 699556 433292 699612
rect 433292 699556 433296 699612
rect 433232 699552 433296 699556
rect 433312 699612 433376 699616
rect 433312 699556 433316 699612
rect 433316 699556 433372 699612
rect 433372 699556 433376 699612
rect 433312 699552 433376 699556
rect 468832 699612 468896 699616
rect 468832 699556 468836 699612
rect 468836 699556 468892 699612
rect 468892 699556 468896 699612
rect 468832 699552 468896 699556
rect 468912 699612 468976 699616
rect 468912 699556 468916 699612
rect 468916 699556 468972 699612
rect 468972 699556 468976 699612
rect 468912 699552 468976 699556
rect 468992 699612 469056 699616
rect 468992 699556 468996 699612
rect 468996 699556 469052 699612
rect 469052 699556 469056 699612
rect 468992 699552 469056 699556
rect 469072 699612 469136 699616
rect 469072 699556 469076 699612
rect 469076 699556 469132 699612
rect 469132 699556 469136 699612
rect 469072 699552 469136 699556
rect 469152 699612 469216 699616
rect 469152 699556 469156 699612
rect 469156 699556 469212 699612
rect 469212 699556 469216 699612
rect 469152 699552 469216 699556
rect 469232 699612 469296 699616
rect 469232 699556 469236 699612
rect 469236 699556 469292 699612
rect 469292 699556 469296 699612
rect 469232 699552 469296 699556
rect 469312 699612 469376 699616
rect 469312 699556 469316 699612
rect 469316 699556 469372 699612
rect 469372 699556 469376 699612
rect 469312 699552 469376 699556
rect 504832 699612 504896 699616
rect 504832 699556 504836 699612
rect 504836 699556 504892 699612
rect 504892 699556 504896 699612
rect 504832 699552 504896 699556
rect 504912 699612 504976 699616
rect 504912 699556 504916 699612
rect 504916 699556 504972 699612
rect 504972 699556 504976 699612
rect 504912 699552 504976 699556
rect 504992 699612 505056 699616
rect 504992 699556 504996 699612
rect 504996 699556 505052 699612
rect 505052 699556 505056 699612
rect 504992 699552 505056 699556
rect 505072 699612 505136 699616
rect 505072 699556 505076 699612
rect 505076 699556 505132 699612
rect 505132 699556 505136 699612
rect 505072 699552 505136 699556
rect 505152 699612 505216 699616
rect 505152 699556 505156 699612
rect 505156 699556 505212 699612
rect 505212 699556 505216 699612
rect 505152 699552 505216 699556
rect 505232 699612 505296 699616
rect 505232 699556 505236 699612
rect 505236 699556 505292 699612
rect 505292 699556 505296 699612
rect 505232 699552 505296 699556
rect 505312 699612 505376 699616
rect 505312 699556 505316 699612
rect 505316 699556 505372 699612
rect 505372 699556 505376 699612
rect 505312 699552 505376 699556
rect 540832 699612 540896 699616
rect 540832 699556 540836 699612
rect 540836 699556 540892 699612
rect 540892 699556 540896 699612
rect 540832 699552 540896 699556
rect 540912 699612 540976 699616
rect 540912 699556 540916 699612
rect 540916 699556 540972 699612
rect 540972 699556 540976 699612
rect 540912 699552 540976 699556
rect 540992 699612 541056 699616
rect 540992 699556 540996 699612
rect 540996 699556 541052 699612
rect 541052 699556 541056 699612
rect 540992 699552 541056 699556
rect 541072 699612 541136 699616
rect 541072 699556 541076 699612
rect 541076 699556 541132 699612
rect 541132 699556 541136 699612
rect 541072 699552 541136 699556
rect 541152 699612 541216 699616
rect 541152 699556 541156 699612
rect 541156 699556 541212 699612
rect 541212 699556 541216 699612
rect 541152 699552 541216 699556
rect 541232 699612 541296 699616
rect 541232 699556 541236 699612
rect 541236 699556 541292 699612
rect 541292 699556 541296 699612
rect 541232 699552 541296 699556
rect 541312 699612 541376 699616
rect 541312 699556 541316 699612
rect 541316 699556 541372 699612
rect 541372 699556 541376 699612
rect 541312 699552 541376 699556
rect 576832 699612 576896 699616
rect 576832 699556 576836 699612
rect 576836 699556 576892 699612
rect 576892 699556 576896 699612
rect 576832 699552 576896 699556
rect 576912 699612 576976 699616
rect 576912 699556 576916 699612
rect 576916 699556 576972 699612
rect 576972 699556 576976 699612
rect 576912 699552 576976 699556
rect 576992 699612 577056 699616
rect 576992 699556 576996 699612
rect 576996 699556 577052 699612
rect 577052 699556 577056 699612
rect 576992 699552 577056 699556
rect 577072 699612 577136 699616
rect 577072 699556 577076 699612
rect 577076 699556 577132 699612
rect 577132 699556 577136 699612
rect 577072 699552 577136 699556
rect 577152 699612 577216 699616
rect 577152 699556 577156 699612
rect 577156 699556 577212 699612
rect 577212 699556 577216 699612
rect 577152 699552 577216 699556
rect 577232 699612 577296 699616
rect 577232 699556 577236 699612
rect 577236 699556 577292 699612
rect 577292 699556 577296 699612
rect 577232 699552 577296 699556
rect 577312 699612 577376 699616
rect 577312 699556 577316 699612
rect 577316 699556 577372 699612
rect 577372 699556 577376 699612
rect 577312 699552 577376 699556
rect 282868 699076 282932 699140
rect 18832 699068 18896 699072
rect 18832 699012 18836 699068
rect 18836 699012 18892 699068
rect 18892 699012 18896 699068
rect 18832 699008 18896 699012
rect 18912 699068 18976 699072
rect 18912 699012 18916 699068
rect 18916 699012 18972 699068
rect 18972 699012 18976 699068
rect 18912 699008 18976 699012
rect 18992 699068 19056 699072
rect 18992 699012 18996 699068
rect 18996 699012 19052 699068
rect 19052 699012 19056 699068
rect 18992 699008 19056 699012
rect 19072 699068 19136 699072
rect 19072 699012 19076 699068
rect 19076 699012 19132 699068
rect 19132 699012 19136 699068
rect 19072 699008 19136 699012
rect 19152 699068 19216 699072
rect 19152 699012 19156 699068
rect 19156 699012 19212 699068
rect 19212 699012 19216 699068
rect 19152 699008 19216 699012
rect 19232 699068 19296 699072
rect 19232 699012 19236 699068
rect 19236 699012 19292 699068
rect 19292 699012 19296 699068
rect 19232 699008 19296 699012
rect 19312 699068 19376 699072
rect 19312 699012 19316 699068
rect 19316 699012 19372 699068
rect 19372 699012 19376 699068
rect 19312 699008 19376 699012
rect 54832 699068 54896 699072
rect 54832 699012 54836 699068
rect 54836 699012 54892 699068
rect 54892 699012 54896 699068
rect 54832 699008 54896 699012
rect 54912 699068 54976 699072
rect 54912 699012 54916 699068
rect 54916 699012 54972 699068
rect 54972 699012 54976 699068
rect 54912 699008 54976 699012
rect 54992 699068 55056 699072
rect 54992 699012 54996 699068
rect 54996 699012 55052 699068
rect 55052 699012 55056 699068
rect 54992 699008 55056 699012
rect 55072 699068 55136 699072
rect 55072 699012 55076 699068
rect 55076 699012 55132 699068
rect 55132 699012 55136 699068
rect 55072 699008 55136 699012
rect 55152 699068 55216 699072
rect 55152 699012 55156 699068
rect 55156 699012 55212 699068
rect 55212 699012 55216 699068
rect 55152 699008 55216 699012
rect 55232 699068 55296 699072
rect 55232 699012 55236 699068
rect 55236 699012 55292 699068
rect 55292 699012 55296 699068
rect 55232 699008 55296 699012
rect 55312 699068 55376 699072
rect 55312 699012 55316 699068
rect 55316 699012 55372 699068
rect 55372 699012 55376 699068
rect 55312 699008 55376 699012
rect 90832 699068 90896 699072
rect 90832 699012 90836 699068
rect 90836 699012 90892 699068
rect 90892 699012 90896 699068
rect 90832 699008 90896 699012
rect 90912 699068 90976 699072
rect 90912 699012 90916 699068
rect 90916 699012 90972 699068
rect 90972 699012 90976 699068
rect 90912 699008 90976 699012
rect 90992 699068 91056 699072
rect 90992 699012 90996 699068
rect 90996 699012 91052 699068
rect 91052 699012 91056 699068
rect 90992 699008 91056 699012
rect 91072 699068 91136 699072
rect 91072 699012 91076 699068
rect 91076 699012 91132 699068
rect 91132 699012 91136 699068
rect 91072 699008 91136 699012
rect 91152 699068 91216 699072
rect 91152 699012 91156 699068
rect 91156 699012 91212 699068
rect 91212 699012 91216 699068
rect 91152 699008 91216 699012
rect 91232 699068 91296 699072
rect 91232 699012 91236 699068
rect 91236 699012 91292 699068
rect 91292 699012 91296 699068
rect 91232 699008 91296 699012
rect 91312 699068 91376 699072
rect 91312 699012 91316 699068
rect 91316 699012 91372 699068
rect 91372 699012 91376 699068
rect 91312 699008 91376 699012
rect 126832 699068 126896 699072
rect 126832 699012 126836 699068
rect 126836 699012 126892 699068
rect 126892 699012 126896 699068
rect 126832 699008 126896 699012
rect 126912 699068 126976 699072
rect 126912 699012 126916 699068
rect 126916 699012 126972 699068
rect 126972 699012 126976 699068
rect 126912 699008 126976 699012
rect 126992 699068 127056 699072
rect 126992 699012 126996 699068
rect 126996 699012 127052 699068
rect 127052 699012 127056 699068
rect 126992 699008 127056 699012
rect 127072 699068 127136 699072
rect 127072 699012 127076 699068
rect 127076 699012 127132 699068
rect 127132 699012 127136 699068
rect 127072 699008 127136 699012
rect 127152 699068 127216 699072
rect 127152 699012 127156 699068
rect 127156 699012 127212 699068
rect 127212 699012 127216 699068
rect 127152 699008 127216 699012
rect 127232 699068 127296 699072
rect 127232 699012 127236 699068
rect 127236 699012 127292 699068
rect 127292 699012 127296 699068
rect 127232 699008 127296 699012
rect 127312 699068 127376 699072
rect 127312 699012 127316 699068
rect 127316 699012 127372 699068
rect 127372 699012 127376 699068
rect 127312 699008 127376 699012
rect 162832 699068 162896 699072
rect 162832 699012 162836 699068
rect 162836 699012 162892 699068
rect 162892 699012 162896 699068
rect 162832 699008 162896 699012
rect 162912 699068 162976 699072
rect 162912 699012 162916 699068
rect 162916 699012 162972 699068
rect 162972 699012 162976 699068
rect 162912 699008 162976 699012
rect 162992 699068 163056 699072
rect 162992 699012 162996 699068
rect 162996 699012 163052 699068
rect 163052 699012 163056 699068
rect 162992 699008 163056 699012
rect 163072 699068 163136 699072
rect 163072 699012 163076 699068
rect 163076 699012 163132 699068
rect 163132 699012 163136 699068
rect 163072 699008 163136 699012
rect 163152 699068 163216 699072
rect 163152 699012 163156 699068
rect 163156 699012 163212 699068
rect 163212 699012 163216 699068
rect 163152 699008 163216 699012
rect 163232 699068 163296 699072
rect 163232 699012 163236 699068
rect 163236 699012 163292 699068
rect 163292 699012 163296 699068
rect 163232 699008 163296 699012
rect 163312 699068 163376 699072
rect 163312 699012 163316 699068
rect 163316 699012 163372 699068
rect 163372 699012 163376 699068
rect 163312 699008 163376 699012
rect 198832 699068 198896 699072
rect 198832 699012 198836 699068
rect 198836 699012 198892 699068
rect 198892 699012 198896 699068
rect 198832 699008 198896 699012
rect 198912 699068 198976 699072
rect 198912 699012 198916 699068
rect 198916 699012 198972 699068
rect 198972 699012 198976 699068
rect 198912 699008 198976 699012
rect 198992 699068 199056 699072
rect 198992 699012 198996 699068
rect 198996 699012 199052 699068
rect 199052 699012 199056 699068
rect 198992 699008 199056 699012
rect 199072 699068 199136 699072
rect 199072 699012 199076 699068
rect 199076 699012 199132 699068
rect 199132 699012 199136 699068
rect 199072 699008 199136 699012
rect 199152 699068 199216 699072
rect 199152 699012 199156 699068
rect 199156 699012 199212 699068
rect 199212 699012 199216 699068
rect 199152 699008 199216 699012
rect 199232 699068 199296 699072
rect 199232 699012 199236 699068
rect 199236 699012 199292 699068
rect 199292 699012 199296 699068
rect 199232 699008 199296 699012
rect 199312 699068 199376 699072
rect 199312 699012 199316 699068
rect 199316 699012 199372 699068
rect 199372 699012 199376 699068
rect 199312 699008 199376 699012
rect 234832 699068 234896 699072
rect 234832 699012 234836 699068
rect 234836 699012 234892 699068
rect 234892 699012 234896 699068
rect 234832 699008 234896 699012
rect 234912 699068 234976 699072
rect 234912 699012 234916 699068
rect 234916 699012 234972 699068
rect 234972 699012 234976 699068
rect 234912 699008 234976 699012
rect 234992 699068 235056 699072
rect 234992 699012 234996 699068
rect 234996 699012 235052 699068
rect 235052 699012 235056 699068
rect 234992 699008 235056 699012
rect 235072 699068 235136 699072
rect 235072 699012 235076 699068
rect 235076 699012 235132 699068
rect 235132 699012 235136 699068
rect 235072 699008 235136 699012
rect 235152 699068 235216 699072
rect 235152 699012 235156 699068
rect 235156 699012 235212 699068
rect 235212 699012 235216 699068
rect 235152 699008 235216 699012
rect 235232 699068 235296 699072
rect 235232 699012 235236 699068
rect 235236 699012 235292 699068
rect 235292 699012 235296 699068
rect 235232 699008 235296 699012
rect 235312 699068 235376 699072
rect 235312 699012 235316 699068
rect 235316 699012 235372 699068
rect 235372 699012 235376 699068
rect 235312 699008 235376 699012
rect 270832 699068 270896 699072
rect 270832 699012 270836 699068
rect 270836 699012 270892 699068
rect 270892 699012 270896 699068
rect 270832 699008 270896 699012
rect 270912 699068 270976 699072
rect 270912 699012 270916 699068
rect 270916 699012 270972 699068
rect 270972 699012 270976 699068
rect 270912 699008 270976 699012
rect 270992 699068 271056 699072
rect 270992 699012 270996 699068
rect 270996 699012 271052 699068
rect 271052 699012 271056 699068
rect 270992 699008 271056 699012
rect 271072 699068 271136 699072
rect 271072 699012 271076 699068
rect 271076 699012 271132 699068
rect 271132 699012 271136 699068
rect 271072 699008 271136 699012
rect 271152 699068 271216 699072
rect 271152 699012 271156 699068
rect 271156 699012 271212 699068
rect 271212 699012 271216 699068
rect 271152 699008 271216 699012
rect 271232 699068 271296 699072
rect 271232 699012 271236 699068
rect 271236 699012 271292 699068
rect 271292 699012 271296 699068
rect 271232 699008 271296 699012
rect 271312 699068 271376 699072
rect 271312 699012 271316 699068
rect 271316 699012 271372 699068
rect 271372 699012 271376 699068
rect 271312 699008 271376 699012
rect 306832 699068 306896 699072
rect 306832 699012 306836 699068
rect 306836 699012 306892 699068
rect 306892 699012 306896 699068
rect 306832 699008 306896 699012
rect 306912 699068 306976 699072
rect 306912 699012 306916 699068
rect 306916 699012 306972 699068
rect 306972 699012 306976 699068
rect 306912 699008 306976 699012
rect 306992 699068 307056 699072
rect 306992 699012 306996 699068
rect 306996 699012 307052 699068
rect 307052 699012 307056 699068
rect 306992 699008 307056 699012
rect 307072 699068 307136 699072
rect 307072 699012 307076 699068
rect 307076 699012 307132 699068
rect 307132 699012 307136 699068
rect 307072 699008 307136 699012
rect 307152 699068 307216 699072
rect 307152 699012 307156 699068
rect 307156 699012 307212 699068
rect 307212 699012 307216 699068
rect 307152 699008 307216 699012
rect 307232 699068 307296 699072
rect 307232 699012 307236 699068
rect 307236 699012 307292 699068
rect 307292 699012 307296 699068
rect 307232 699008 307296 699012
rect 307312 699068 307376 699072
rect 307312 699012 307316 699068
rect 307316 699012 307372 699068
rect 307372 699012 307376 699068
rect 307312 699008 307376 699012
rect 342832 699068 342896 699072
rect 342832 699012 342836 699068
rect 342836 699012 342892 699068
rect 342892 699012 342896 699068
rect 342832 699008 342896 699012
rect 342912 699068 342976 699072
rect 342912 699012 342916 699068
rect 342916 699012 342972 699068
rect 342972 699012 342976 699068
rect 342912 699008 342976 699012
rect 342992 699068 343056 699072
rect 342992 699012 342996 699068
rect 342996 699012 343052 699068
rect 343052 699012 343056 699068
rect 342992 699008 343056 699012
rect 343072 699068 343136 699072
rect 343072 699012 343076 699068
rect 343076 699012 343132 699068
rect 343132 699012 343136 699068
rect 343072 699008 343136 699012
rect 343152 699068 343216 699072
rect 343152 699012 343156 699068
rect 343156 699012 343212 699068
rect 343212 699012 343216 699068
rect 343152 699008 343216 699012
rect 343232 699068 343296 699072
rect 343232 699012 343236 699068
rect 343236 699012 343292 699068
rect 343292 699012 343296 699068
rect 343232 699008 343296 699012
rect 343312 699068 343376 699072
rect 343312 699012 343316 699068
rect 343316 699012 343372 699068
rect 343372 699012 343376 699068
rect 343312 699008 343376 699012
rect 378832 699068 378896 699072
rect 378832 699012 378836 699068
rect 378836 699012 378892 699068
rect 378892 699012 378896 699068
rect 378832 699008 378896 699012
rect 378912 699068 378976 699072
rect 378912 699012 378916 699068
rect 378916 699012 378972 699068
rect 378972 699012 378976 699068
rect 378912 699008 378976 699012
rect 378992 699068 379056 699072
rect 378992 699012 378996 699068
rect 378996 699012 379052 699068
rect 379052 699012 379056 699068
rect 378992 699008 379056 699012
rect 379072 699068 379136 699072
rect 379072 699012 379076 699068
rect 379076 699012 379132 699068
rect 379132 699012 379136 699068
rect 379072 699008 379136 699012
rect 379152 699068 379216 699072
rect 379152 699012 379156 699068
rect 379156 699012 379212 699068
rect 379212 699012 379216 699068
rect 379152 699008 379216 699012
rect 379232 699068 379296 699072
rect 379232 699012 379236 699068
rect 379236 699012 379292 699068
rect 379292 699012 379296 699068
rect 379232 699008 379296 699012
rect 379312 699068 379376 699072
rect 379312 699012 379316 699068
rect 379316 699012 379372 699068
rect 379372 699012 379376 699068
rect 379312 699008 379376 699012
rect 414832 699068 414896 699072
rect 414832 699012 414836 699068
rect 414836 699012 414892 699068
rect 414892 699012 414896 699068
rect 414832 699008 414896 699012
rect 414912 699068 414976 699072
rect 414912 699012 414916 699068
rect 414916 699012 414972 699068
rect 414972 699012 414976 699068
rect 414912 699008 414976 699012
rect 414992 699068 415056 699072
rect 414992 699012 414996 699068
rect 414996 699012 415052 699068
rect 415052 699012 415056 699068
rect 414992 699008 415056 699012
rect 415072 699068 415136 699072
rect 415072 699012 415076 699068
rect 415076 699012 415132 699068
rect 415132 699012 415136 699068
rect 415072 699008 415136 699012
rect 415152 699068 415216 699072
rect 415152 699012 415156 699068
rect 415156 699012 415212 699068
rect 415212 699012 415216 699068
rect 415152 699008 415216 699012
rect 415232 699068 415296 699072
rect 415232 699012 415236 699068
rect 415236 699012 415292 699068
rect 415292 699012 415296 699068
rect 415232 699008 415296 699012
rect 415312 699068 415376 699072
rect 415312 699012 415316 699068
rect 415316 699012 415372 699068
rect 415372 699012 415376 699068
rect 415312 699008 415376 699012
rect 450832 699068 450896 699072
rect 450832 699012 450836 699068
rect 450836 699012 450892 699068
rect 450892 699012 450896 699068
rect 450832 699008 450896 699012
rect 450912 699068 450976 699072
rect 450912 699012 450916 699068
rect 450916 699012 450972 699068
rect 450972 699012 450976 699068
rect 450912 699008 450976 699012
rect 450992 699068 451056 699072
rect 450992 699012 450996 699068
rect 450996 699012 451052 699068
rect 451052 699012 451056 699068
rect 450992 699008 451056 699012
rect 451072 699068 451136 699072
rect 451072 699012 451076 699068
rect 451076 699012 451132 699068
rect 451132 699012 451136 699068
rect 451072 699008 451136 699012
rect 451152 699068 451216 699072
rect 451152 699012 451156 699068
rect 451156 699012 451212 699068
rect 451212 699012 451216 699068
rect 451152 699008 451216 699012
rect 451232 699068 451296 699072
rect 451232 699012 451236 699068
rect 451236 699012 451292 699068
rect 451292 699012 451296 699068
rect 451232 699008 451296 699012
rect 451312 699068 451376 699072
rect 451312 699012 451316 699068
rect 451316 699012 451372 699068
rect 451372 699012 451376 699068
rect 451312 699008 451376 699012
rect 486832 699068 486896 699072
rect 486832 699012 486836 699068
rect 486836 699012 486892 699068
rect 486892 699012 486896 699068
rect 486832 699008 486896 699012
rect 486912 699068 486976 699072
rect 486912 699012 486916 699068
rect 486916 699012 486972 699068
rect 486972 699012 486976 699068
rect 486912 699008 486976 699012
rect 486992 699068 487056 699072
rect 486992 699012 486996 699068
rect 486996 699012 487052 699068
rect 487052 699012 487056 699068
rect 486992 699008 487056 699012
rect 487072 699068 487136 699072
rect 487072 699012 487076 699068
rect 487076 699012 487132 699068
rect 487132 699012 487136 699068
rect 487072 699008 487136 699012
rect 487152 699068 487216 699072
rect 487152 699012 487156 699068
rect 487156 699012 487212 699068
rect 487212 699012 487216 699068
rect 487152 699008 487216 699012
rect 487232 699068 487296 699072
rect 487232 699012 487236 699068
rect 487236 699012 487292 699068
rect 487292 699012 487296 699068
rect 487232 699008 487296 699012
rect 487312 699068 487376 699072
rect 487312 699012 487316 699068
rect 487316 699012 487372 699068
rect 487372 699012 487376 699068
rect 487312 699008 487376 699012
rect 522832 699068 522896 699072
rect 522832 699012 522836 699068
rect 522836 699012 522892 699068
rect 522892 699012 522896 699068
rect 522832 699008 522896 699012
rect 522912 699068 522976 699072
rect 522912 699012 522916 699068
rect 522916 699012 522972 699068
rect 522972 699012 522976 699068
rect 522912 699008 522976 699012
rect 522992 699068 523056 699072
rect 522992 699012 522996 699068
rect 522996 699012 523052 699068
rect 523052 699012 523056 699068
rect 522992 699008 523056 699012
rect 523072 699068 523136 699072
rect 523072 699012 523076 699068
rect 523076 699012 523132 699068
rect 523132 699012 523136 699068
rect 523072 699008 523136 699012
rect 523152 699068 523216 699072
rect 523152 699012 523156 699068
rect 523156 699012 523212 699068
rect 523212 699012 523216 699068
rect 523152 699008 523216 699012
rect 523232 699068 523296 699072
rect 523232 699012 523236 699068
rect 523236 699012 523292 699068
rect 523292 699012 523296 699068
rect 523232 699008 523296 699012
rect 523312 699068 523376 699072
rect 523312 699012 523316 699068
rect 523316 699012 523372 699068
rect 523372 699012 523376 699068
rect 523312 699008 523376 699012
rect 558832 699068 558896 699072
rect 558832 699012 558836 699068
rect 558836 699012 558892 699068
rect 558892 699012 558896 699068
rect 558832 699008 558896 699012
rect 558912 699068 558976 699072
rect 558912 699012 558916 699068
rect 558916 699012 558972 699068
rect 558972 699012 558976 699068
rect 558912 699008 558976 699012
rect 558992 699068 559056 699072
rect 558992 699012 558996 699068
rect 558996 699012 559052 699068
rect 559052 699012 559056 699068
rect 558992 699008 559056 699012
rect 559072 699068 559136 699072
rect 559072 699012 559076 699068
rect 559076 699012 559132 699068
rect 559132 699012 559136 699068
rect 559072 699008 559136 699012
rect 559152 699068 559216 699072
rect 559152 699012 559156 699068
rect 559156 699012 559212 699068
rect 559212 699012 559216 699068
rect 559152 699008 559216 699012
rect 559232 699068 559296 699072
rect 559232 699012 559236 699068
rect 559236 699012 559292 699068
rect 559292 699012 559296 699068
rect 559232 699008 559296 699012
rect 559312 699068 559376 699072
rect 559312 699012 559316 699068
rect 559316 699012 559372 699068
rect 559372 699012 559376 699068
rect 559312 699008 559376 699012
rect 86724 698804 86788 698868
rect 447180 698804 447244 698868
rect 282868 698532 282932 698596
rect 36832 698524 36896 698528
rect 36832 698468 36836 698524
rect 36836 698468 36892 698524
rect 36892 698468 36896 698524
rect 36832 698464 36896 698468
rect 36912 698524 36976 698528
rect 36912 698468 36916 698524
rect 36916 698468 36972 698524
rect 36972 698468 36976 698524
rect 36912 698464 36976 698468
rect 36992 698524 37056 698528
rect 36992 698468 36996 698524
rect 36996 698468 37052 698524
rect 37052 698468 37056 698524
rect 36992 698464 37056 698468
rect 37072 698524 37136 698528
rect 37072 698468 37076 698524
rect 37076 698468 37132 698524
rect 37132 698468 37136 698524
rect 37072 698464 37136 698468
rect 37152 698524 37216 698528
rect 37152 698468 37156 698524
rect 37156 698468 37212 698524
rect 37212 698468 37216 698524
rect 37152 698464 37216 698468
rect 37232 698524 37296 698528
rect 37232 698468 37236 698524
rect 37236 698468 37292 698524
rect 37292 698468 37296 698524
rect 37232 698464 37296 698468
rect 37312 698524 37376 698528
rect 37312 698468 37316 698524
rect 37316 698468 37372 698524
rect 37372 698468 37376 698524
rect 37312 698464 37376 698468
rect 72832 698524 72896 698528
rect 72832 698468 72836 698524
rect 72836 698468 72892 698524
rect 72892 698468 72896 698524
rect 72832 698464 72896 698468
rect 72912 698524 72976 698528
rect 72912 698468 72916 698524
rect 72916 698468 72972 698524
rect 72972 698468 72976 698524
rect 72912 698464 72976 698468
rect 72992 698524 73056 698528
rect 72992 698468 72996 698524
rect 72996 698468 73052 698524
rect 73052 698468 73056 698524
rect 72992 698464 73056 698468
rect 73072 698524 73136 698528
rect 73072 698468 73076 698524
rect 73076 698468 73132 698524
rect 73132 698468 73136 698524
rect 73072 698464 73136 698468
rect 73152 698524 73216 698528
rect 73152 698468 73156 698524
rect 73156 698468 73212 698524
rect 73212 698468 73216 698524
rect 73152 698464 73216 698468
rect 73232 698524 73296 698528
rect 73232 698468 73236 698524
rect 73236 698468 73292 698524
rect 73292 698468 73296 698524
rect 73232 698464 73296 698468
rect 73312 698524 73376 698528
rect 73312 698468 73316 698524
rect 73316 698468 73372 698524
rect 73372 698468 73376 698524
rect 73312 698464 73376 698468
rect 108832 698524 108896 698528
rect 108832 698468 108836 698524
rect 108836 698468 108892 698524
rect 108892 698468 108896 698524
rect 108832 698464 108896 698468
rect 108912 698524 108976 698528
rect 108912 698468 108916 698524
rect 108916 698468 108972 698524
rect 108972 698468 108976 698524
rect 108912 698464 108976 698468
rect 108992 698524 109056 698528
rect 108992 698468 108996 698524
rect 108996 698468 109052 698524
rect 109052 698468 109056 698524
rect 108992 698464 109056 698468
rect 109072 698524 109136 698528
rect 109072 698468 109076 698524
rect 109076 698468 109132 698524
rect 109132 698468 109136 698524
rect 109072 698464 109136 698468
rect 109152 698524 109216 698528
rect 109152 698468 109156 698524
rect 109156 698468 109212 698524
rect 109212 698468 109216 698524
rect 109152 698464 109216 698468
rect 109232 698524 109296 698528
rect 109232 698468 109236 698524
rect 109236 698468 109292 698524
rect 109292 698468 109296 698524
rect 109232 698464 109296 698468
rect 109312 698524 109376 698528
rect 109312 698468 109316 698524
rect 109316 698468 109372 698524
rect 109372 698468 109376 698524
rect 109312 698464 109376 698468
rect 144832 698524 144896 698528
rect 144832 698468 144836 698524
rect 144836 698468 144892 698524
rect 144892 698468 144896 698524
rect 144832 698464 144896 698468
rect 144912 698524 144976 698528
rect 144912 698468 144916 698524
rect 144916 698468 144972 698524
rect 144972 698468 144976 698524
rect 144912 698464 144976 698468
rect 144992 698524 145056 698528
rect 144992 698468 144996 698524
rect 144996 698468 145052 698524
rect 145052 698468 145056 698524
rect 144992 698464 145056 698468
rect 145072 698524 145136 698528
rect 145072 698468 145076 698524
rect 145076 698468 145132 698524
rect 145132 698468 145136 698524
rect 145072 698464 145136 698468
rect 145152 698524 145216 698528
rect 145152 698468 145156 698524
rect 145156 698468 145212 698524
rect 145212 698468 145216 698524
rect 145152 698464 145216 698468
rect 145232 698524 145296 698528
rect 145232 698468 145236 698524
rect 145236 698468 145292 698524
rect 145292 698468 145296 698524
rect 145232 698464 145296 698468
rect 145312 698524 145376 698528
rect 145312 698468 145316 698524
rect 145316 698468 145372 698524
rect 145372 698468 145376 698524
rect 145312 698464 145376 698468
rect 180832 698524 180896 698528
rect 180832 698468 180836 698524
rect 180836 698468 180892 698524
rect 180892 698468 180896 698524
rect 180832 698464 180896 698468
rect 180912 698524 180976 698528
rect 180912 698468 180916 698524
rect 180916 698468 180972 698524
rect 180972 698468 180976 698524
rect 180912 698464 180976 698468
rect 180992 698524 181056 698528
rect 180992 698468 180996 698524
rect 180996 698468 181052 698524
rect 181052 698468 181056 698524
rect 180992 698464 181056 698468
rect 181072 698524 181136 698528
rect 181072 698468 181076 698524
rect 181076 698468 181132 698524
rect 181132 698468 181136 698524
rect 181072 698464 181136 698468
rect 181152 698524 181216 698528
rect 181152 698468 181156 698524
rect 181156 698468 181212 698524
rect 181212 698468 181216 698524
rect 181152 698464 181216 698468
rect 181232 698524 181296 698528
rect 181232 698468 181236 698524
rect 181236 698468 181292 698524
rect 181292 698468 181296 698524
rect 181232 698464 181296 698468
rect 181312 698524 181376 698528
rect 181312 698468 181316 698524
rect 181316 698468 181372 698524
rect 181372 698468 181376 698524
rect 181312 698464 181376 698468
rect 216832 698524 216896 698528
rect 216832 698468 216836 698524
rect 216836 698468 216892 698524
rect 216892 698468 216896 698524
rect 216832 698464 216896 698468
rect 216912 698524 216976 698528
rect 216912 698468 216916 698524
rect 216916 698468 216972 698524
rect 216972 698468 216976 698524
rect 216912 698464 216976 698468
rect 216992 698524 217056 698528
rect 216992 698468 216996 698524
rect 216996 698468 217052 698524
rect 217052 698468 217056 698524
rect 216992 698464 217056 698468
rect 217072 698524 217136 698528
rect 217072 698468 217076 698524
rect 217076 698468 217132 698524
rect 217132 698468 217136 698524
rect 217072 698464 217136 698468
rect 217152 698524 217216 698528
rect 217152 698468 217156 698524
rect 217156 698468 217212 698524
rect 217212 698468 217216 698524
rect 217152 698464 217216 698468
rect 217232 698524 217296 698528
rect 217232 698468 217236 698524
rect 217236 698468 217292 698524
rect 217292 698468 217296 698524
rect 217232 698464 217296 698468
rect 217312 698524 217376 698528
rect 217312 698468 217316 698524
rect 217316 698468 217372 698524
rect 217372 698468 217376 698524
rect 217312 698464 217376 698468
rect 252832 698524 252896 698528
rect 252832 698468 252836 698524
rect 252836 698468 252892 698524
rect 252892 698468 252896 698524
rect 252832 698464 252896 698468
rect 252912 698524 252976 698528
rect 252912 698468 252916 698524
rect 252916 698468 252972 698524
rect 252972 698468 252976 698524
rect 252912 698464 252976 698468
rect 252992 698524 253056 698528
rect 252992 698468 252996 698524
rect 252996 698468 253052 698524
rect 253052 698468 253056 698524
rect 252992 698464 253056 698468
rect 253072 698524 253136 698528
rect 253072 698468 253076 698524
rect 253076 698468 253132 698524
rect 253132 698468 253136 698524
rect 253072 698464 253136 698468
rect 253152 698524 253216 698528
rect 253152 698468 253156 698524
rect 253156 698468 253212 698524
rect 253212 698468 253216 698524
rect 253152 698464 253216 698468
rect 253232 698524 253296 698528
rect 253232 698468 253236 698524
rect 253236 698468 253292 698524
rect 253292 698468 253296 698524
rect 253232 698464 253296 698468
rect 253312 698524 253376 698528
rect 253312 698468 253316 698524
rect 253316 698468 253372 698524
rect 253372 698468 253376 698524
rect 253312 698464 253376 698468
rect 288832 698524 288896 698528
rect 288832 698468 288836 698524
rect 288836 698468 288892 698524
rect 288892 698468 288896 698524
rect 288832 698464 288896 698468
rect 288912 698524 288976 698528
rect 288912 698468 288916 698524
rect 288916 698468 288972 698524
rect 288972 698468 288976 698524
rect 288912 698464 288976 698468
rect 288992 698524 289056 698528
rect 288992 698468 288996 698524
rect 288996 698468 289052 698524
rect 289052 698468 289056 698524
rect 288992 698464 289056 698468
rect 289072 698524 289136 698528
rect 289072 698468 289076 698524
rect 289076 698468 289132 698524
rect 289132 698468 289136 698524
rect 289072 698464 289136 698468
rect 289152 698524 289216 698528
rect 289152 698468 289156 698524
rect 289156 698468 289212 698524
rect 289212 698468 289216 698524
rect 289152 698464 289216 698468
rect 289232 698524 289296 698528
rect 289232 698468 289236 698524
rect 289236 698468 289292 698524
rect 289292 698468 289296 698524
rect 289232 698464 289296 698468
rect 289312 698524 289376 698528
rect 289312 698468 289316 698524
rect 289316 698468 289372 698524
rect 289372 698468 289376 698524
rect 289312 698464 289376 698468
rect 324832 698524 324896 698528
rect 324832 698468 324836 698524
rect 324836 698468 324892 698524
rect 324892 698468 324896 698524
rect 324832 698464 324896 698468
rect 324912 698524 324976 698528
rect 324912 698468 324916 698524
rect 324916 698468 324972 698524
rect 324972 698468 324976 698524
rect 324912 698464 324976 698468
rect 324992 698524 325056 698528
rect 324992 698468 324996 698524
rect 324996 698468 325052 698524
rect 325052 698468 325056 698524
rect 324992 698464 325056 698468
rect 325072 698524 325136 698528
rect 325072 698468 325076 698524
rect 325076 698468 325132 698524
rect 325132 698468 325136 698524
rect 325072 698464 325136 698468
rect 325152 698524 325216 698528
rect 325152 698468 325156 698524
rect 325156 698468 325212 698524
rect 325212 698468 325216 698524
rect 325152 698464 325216 698468
rect 325232 698524 325296 698528
rect 325232 698468 325236 698524
rect 325236 698468 325292 698524
rect 325292 698468 325296 698524
rect 325232 698464 325296 698468
rect 325312 698524 325376 698528
rect 325312 698468 325316 698524
rect 325316 698468 325372 698524
rect 325372 698468 325376 698524
rect 325312 698464 325376 698468
rect 360832 698524 360896 698528
rect 360832 698468 360836 698524
rect 360836 698468 360892 698524
rect 360892 698468 360896 698524
rect 360832 698464 360896 698468
rect 360912 698524 360976 698528
rect 360912 698468 360916 698524
rect 360916 698468 360972 698524
rect 360972 698468 360976 698524
rect 360912 698464 360976 698468
rect 360992 698524 361056 698528
rect 360992 698468 360996 698524
rect 360996 698468 361052 698524
rect 361052 698468 361056 698524
rect 360992 698464 361056 698468
rect 361072 698524 361136 698528
rect 361072 698468 361076 698524
rect 361076 698468 361132 698524
rect 361132 698468 361136 698524
rect 361072 698464 361136 698468
rect 361152 698524 361216 698528
rect 361152 698468 361156 698524
rect 361156 698468 361212 698524
rect 361212 698468 361216 698524
rect 361152 698464 361216 698468
rect 361232 698524 361296 698528
rect 361232 698468 361236 698524
rect 361236 698468 361292 698524
rect 361292 698468 361296 698524
rect 361232 698464 361296 698468
rect 361312 698524 361376 698528
rect 361312 698468 361316 698524
rect 361316 698468 361372 698524
rect 361372 698468 361376 698524
rect 361312 698464 361376 698468
rect 396832 698524 396896 698528
rect 396832 698468 396836 698524
rect 396836 698468 396892 698524
rect 396892 698468 396896 698524
rect 396832 698464 396896 698468
rect 396912 698524 396976 698528
rect 396912 698468 396916 698524
rect 396916 698468 396972 698524
rect 396972 698468 396976 698524
rect 396912 698464 396976 698468
rect 396992 698524 397056 698528
rect 396992 698468 396996 698524
rect 396996 698468 397052 698524
rect 397052 698468 397056 698524
rect 396992 698464 397056 698468
rect 397072 698524 397136 698528
rect 397072 698468 397076 698524
rect 397076 698468 397132 698524
rect 397132 698468 397136 698524
rect 397072 698464 397136 698468
rect 397152 698524 397216 698528
rect 397152 698468 397156 698524
rect 397156 698468 397212 698524
rect 397212 698468 397216 698524
rect 397152 698464 397216 698468
rect 397232 698524 397296 698528
rect 397232 698468 397236 698524
rect 397236 698468 397292 698524
rect 397292 698468 397296 698524
rect 397232 698464 397296 698468
rect 397312 698524 397376 698528
rect 397312 698468 397316 698524
rect 397316 698468 397372 698524
rect 397372 698468 397376 698524
rect 397312 698464 397376 698468
rect 432832 698524 432896 698528
rect 432832 698468 432836 698524
rect 432836 698468 432892 698524
rect 432892 698468 432896 698524
rect 432832 698464 432896 698468
rect 432912 698524 432976 698528
rect 432912 698468 432916 698524
rect 432916 698468 432972 698524
rect 432972 698468 432976 698524
rect 432912 698464 432976 698468
rect 432992 698524 433056 698528
rect 432992 698468 432996 698524
rect 432996 698468 433052 698524
rect 433052 698468 433056 698524
rect 432992 698464 433056 698468
rect 433072 698524 433136 698528
rect 433072 698468 433076 698524
rect 433076 698468 433132 698524
rect 433132 698468 433136 698524
rect 433072 698464 433136 698468
rect 433152 698524 433216 698528
rect 433152 698468 433156 698524
rect 433156 698468 433212 698524
rect 433212 698468 433216 698524
rect 433152 698464 433216 698468
rect 433232 698524 433296 698528
rect 433232 698468 433236 698524
rect 433236 698468 433292 698524
rect 433292 698468 433296 698524
rect 433232 698464 433296 698468
rect 433312 698524 433376 698528
rect 433312 698468 433316 698524
rect 433316 698468 433372 698524
rect 433372 698468 433376 698524
rect 433312 698464 433376 698468
rect 468832 698524 468896 698528
rect 468832 698468 468836 698524
rect 468836 698468 468892 698524
rect 468892 698468 468896 698524
rect 468832 698464 468896 698468
rect 468912 698524 468976 698528
rect 468912 698468 468916 698524
rect 468916 698468 468972 698524
rect 468972 698468 468976 698524
rect 468912 698464 468976 698468
rect 468992 698524 469056 698528
rect 468992 698468 468996 698524
rect 468996 698468 469052 698524
rect 469052 698468 469056 698524
rect 468992 698464 469056 698468
rect 469072 698524 469136 698528
rect 469072 698468 469076 698524
rect 469076 698468 469132 698524
rect 469132 698468 469136 698524
rect 469072 698464 469136 698468
rect 469152 698524 469216 698528
rect 469152 698468 469156 698524
rect 469156 698468 469212 698524
rect 469212 698468 469216 698524
rect 469152 698464 469216 698468
rect 469232 698524 469296 698528
rect 469232 698468 469236 698524
rect 469236 698468 469292 698524
rect 469292 698468 469296 698524
rect 469232 698464 469296 698468
rect 469312 698524 469376 698528
rect 469312 698468 469316 698524
rect 469316 698468 469372 698524
rect 469372 698468 469376 698524
rect 469312 698464 469376 698468
rect 504832 698524 504896 698528
rect 504832 698468 504836 698524
rect 504836 698468 504892 698524
rect 504892 698468 504896 698524
rect 504832 698464 504896 698468
rect 504912 698524 504976 698528
rect 504912 698468 504916 698524
rect 504916 698468 504972 698524
rect 504972 698468 504976 698524
rect 504912 698464 504976 698468
rect 504992 698524 505056 698528
rect 504992 698468 504996 698524
rect 504996 698468 505052 698524
rect 505052 698468 505056 698524
rect 504992 698464 505056 698468
rect 505072 698524 505136 698528
rect 505072 698468 505076 698524
rect 505076 698468 505132 698524
rect 505132 698468 505136 698524
rect 505072 698464 505136 698468
rect 505152 698524 505216 698528
rect 505152 698468 505156 698524
rect 505156 698468 505212 698524
rect 505212 698468 505216 698524
rect 505152 698464 505216 698468
rect 505232 698524 505296 698528
rect 505232 698468 505236 698524
rect 505236 698468 505292 698524
rect 505292 698468 505296 698524
rect 505232 698464 505296 698468
rect 505312 698524 505376 698528
rect 505312 698468 505316 698524
rect 505316 698468 505372 698524
rect 505372 698468 505376 698524
rect 505312 698464 505376 698468
rect 540832 698524 540896 698528
rect 540832 698468 540836 698524
rect 540836 698468 540892 698524
rect 540892 698468 540896 698524
rect 540832 698464 540896 698468
rect 540912 698524 540976 698528
rect 540912 698468 540916 698524
rect 540916 698468 540972 698524
rect 540972 698468 540976 698524
rect 540912 698464 540976 698468
rect 540992 698524 541056 698528
rect 540992 698468 540996 698524
rect 540996 698468 541052 698524
rect 541052 698468 541056 698524
rect 540992 698464 541056 698468
rect 541072 698524 541136 698528
rect 541072 698468 541076 698524
rect 541076 698468 541132 698524
rect 541132 698468 541136 698524
rect 541072 698464 541136 698468
rect 541152 698524 541216 698528
rect 541152 698468 541156 698524
rect 541156 698468 541212 698524
rect 541212 698468 541216 698524
rect 541152 698464 541216 698468
rect 541232 698524 541296 698528
rect 541232 698468 541236 698524
rect 541236 698468 541292 698524
rect 541292 698468 541296 698524
rect 541232 698464 541296 698468
rect 541312 698524 541376 698528
rect 541312 698468 541316 698524
rect 541316 698468 541372 698524
rect 541372 698468 541376 698524
rect 541312 698464 541376 698468
rect 576832 698524 576896 698528
rect 576832 698468 576836 698524
rect 576836 698468 576892 698524
rect 576892 698468 576896 698524
rect 576832 698464 576896 698468
rect 576912 698524 576976 698528
rect 576912 698468 576916 698524
rect 576916 698468 576972 698524
rect 576972 698468 576976 698524
rect 576912 698464 576976 698468
rect 576992 698524 577056 698528
rect 576992 698468 576996 698524
rect 576996 698468 577052 698524
rect 577052 698468 577056 698524
rect 576992 698464 577056 698468
rect 577072 698524 577136 698528
rect 577072 698468 577076 698524
rect 577076 698468 577132 698524
rect 577132 698468 577136 698524
rect 577072 698464 577136 698468
rect 577152 698524 577216 698528
rect 577152 698468 577156 698524
rect 577156 698468 577212 698524
rect 577212 698468 577216 698524
rect 577152 698464 577216 698468
rect 577232 698524 577296 698528
rect 577232 698468 577236 698524
rect 577236 698468 577292 698524
rect 577292 698468 577296 698524
rect 577232 698464 577296 698468
rect 577312 698524 577376 698528
rect 577312 698468 577316 698524
rect 577316 698468 577372 698524
rect 577372 698468 577376 698524
rect 577312 698464 577376 698468
rect 71820 698260 71884 698324
rect 15332 695328 15396 695332
rect 15332 695272 15346 695328
rect 15346 695272 15396 695328
rect 15332 695268 15396 695272
rect 179644 695268 179708 695332
rect 521332 695328 521396 695332
rect 521332 695272 521382 695328
rect 521382 695272 521396 695328
rect 521332 695268 521396 695272
rect 231900 694996 231964 695060
rect 236868 694996 236932 695060
rect 251220 694996 251284 695060
rect 256188 694996 256252 695060
rect 357388 694996 357452 695060
rect 362172 694996 362236 695060
rect 434668 694996 434732 695060
rect 439452 694996 439516 695060
rect 137324 694860 137388 694924
rect 141924 694860 141988 694924
rect 196204 694860 196268 694924
rect 202460 694860 202524 694924
rect 273116 694860 273180 694924
rect 278820 694860 278884 694924
rect 280108 694860 280172 694924
rect 283236 694860 283300 694924
rect 292804 694860 292868 694924
rect 299060 694860 299124 694924
rect 346348 694860 346412 694924
rect 351316 694860 351380 694924
rect 370084 694860 370148 694924
rect 376340 694860 376404 694924
rect 389404 694860 389468 694924
rect 395660 694860 395724 694924
rect 500908 694860 500972 694924
rect 505692 694860 505756 694924
rect 134932 694724 134996 694788
rect 138244 694724 138308 694788
rect 142108 694724 142172 694788
rect 151676 694724 151740 694788
rect 152780 694724 152844 694788
rect 159404 694724 159468 694788
rect 222148 694724 222212 694788
rect 226932 694724 226996 694788
rect 106228 694588 106292 694652
rect 115796 694588 115860 694652
rect 164188 694588 164252 694652
rect 173572 694588 173636 694652
rect 176700 694588 176764 694652
rect 15332 694452 15396 694516
rect 42012 694452 42076 694516
rect 9628 694180 9692 694244
rect 9628 693908 9692 693972
rect 19012 693908 19076 693972
rect 42012 694180 42076 694244
rect 85252 694452 85316 694516
rect 79916 694316 79980 694380
rect 80100 694316 80164 694380
rect 98316 694316 98380 694380
rect 64828 694180 64892 694244
rect 76972 694180 77036 694244
rect 86724 694180 86788 694244
rect 37228 694044 37292 694108
rect 41276 694044 41340 694108
rect 41460 694044 41524 694108
rect 27292 693908 27356 693972
rect 28948 693908 29012 693972
rect 64828 693908 64892 693972
rect 115980 694452 116044 694516
rect 98868 694316 98932 694380
rect 106228 694316 106292 694380
rect 106412 694316 106476 694380
rect 120580 694316 120644 694380
rect 130332 694452 130396 694516
rect 134932 694452 134996 694516
rect 151676 694452 151740 694516
rect 151860 694452 151924 694516
rect 166948 694452 167012 694516
rect 176884 694452 176948 694516
rect 186268 694588 186332 694652
rect 215340 694588 215404 694652
rect 224356 694588 224420 694652
rect 236684 694724 236748 694788
rect 241100 694724 241164 694788
rect 246068 694724 246132 694788
rect 243860 694588 243924 694652
rect 256004 694724 256068 694788
rect 264284 694724 264348 694788
rect 270356 694724 270420 694788
rect 318748 694724 318812 694788
rect 328316 694724 328380 694788
rect 350580 694724 350644 694788
rect 357388 694724 357452 694788
rect 263180 694588 263244 694652
rect 273116 694588 273180 694652
rect 282684 694588 282748 694652
rect 311940 694588 312004 694652
rect 320956 694588 321020 694652
rect 332916 694588 332980 694652
rect 106228 694044 106292 694108
rect 120580 694044 120644 694108
rect 130332 694044 130396 694108
rect 141924 694316 141988 694380
rect 142108 694316 142172 694380
rect 146892 694316 146956 694380
rect 152780 694316 152844 694380
rect 137324 694044 137388 694108
rect 138244 694044 138308 694108
rect 146892 694044 146956 694108
rect 152044 694044 152108 694108
rect 164188 694316 164252 694380
rect 179644 694316 179708 694380
rect 186084 694316 186148 694380
rect 202644 694452 202708 694516
rect 196204 694316 196268 694380
rect 214972 694452 215036 694516
rect 215524 694452 215588 694516
rect 222148 694316 222212 694380
rect 226932 694316 226996 694380
rect 173756 694180 173820 694244
rect 176700 694180 176764 694244
rect 215708 694180 215772 694244
rect 231900 694316 231964 694380
rect 232084 694316 232148 694380
rect 235948 694316 236012 694380
rect 159404 694044 159468 694108
rect 166948 694044 167012 694108
rect 176884 694044 176948 694108
rect 185900 694044 185964 694108
rect 186084 694044 186148 694108
rect 186268 694044 186332 694108
rect 186452 694044 186516 694108
rect 205404 694044 205468 694108
rect 205956 694044 206020 694108
rect 214972 694044 215036 694108
rect 215340 694044 215404 694108
rect 224356 694044 224420 694108
rect 241100 694316 241164 694380
rect 246068 694316 246132 694380
rect 251220 694316 251284 694380
rect 251404 694316 251468 694380
rect 255268 694316 255332 694380
rect 265572 694452 265636 694516
rect 299244 694452 299308 694516
rect 236868 694180 236932 694244
rect 245700 694180 245764 694244
rect 236684 694044 236748 694108
rect 243860 694044 243924 694108
rect 246436 694180 246500 694244
rect 270724 694316 270788 694380
rect 283052 694316 283116 694380
rect 283236 694316 283300 694380
rect 292804 694316 292868 694380
rect 311572 694452 311636 694516
rect 312124 694452 312188 694516
rect 318748 694316 318812 694380
rect 328316 694316 328380 694380
rect 256188 694180 256252 694244
rect 264284 694180 264348 694244
rect 270356 694180 270420 694244
rect 256004 694044 256068 694108
rect 263180 694044 263244 694108
rect 265572 694044 265636 694108
rect 270540 694044 270604 694108
rect 278820 694180 278884 694244
rect 282684 694180 282748 694244
rect 312308 694180 312372 694244
rect 333100 694452 333164 694516
rect 338620 694588 338684 694652
rect 340460 694588 340524 694652
rect 346348 694588 346412 694652
rect 359964 694588 360028 694652
rect 434668 694724 434732 694788
rect 492812 694588 492876 694652
rect 500908 694588 500972 694652
rect 531268 694588 531332 694652
rect 86908 693908 86972 693972
rect 87092 693908 87156 693972
rect 270540 693908 270604 693972
rect 270724 693908 270788 693972
rect 279924 694044 279988 694108
rect 283236 694044 283300 694108
rect 302004 694044 302068 694108
rect 302556 694044 302620 694108
rect 311572 694044 311636 694108
rect 311940 694044 312004 694108
rect 320956 694044 321020 694108
rect 333100 694180 333164 694244
rect 341564 694452 341628 694516
rect 376524 694452 376588 694516
rect 338620 694316 338684 694380
rect 332916 694044 332980 694108
rect 340460 694044 340524 694108
rect 350396 694316 350460 694380
rect 350764 694316 350828 694380
rect 351132 694316 351196 694380
rect 341564 694180 341628 694244
rect 350580 694180 350644 694244
rect 351316 694180 351380 694244
rect 359964 694180 360028 694244
rect 350396 694044 350460 694108
rect 362172 694316 362236 694380
rect 370084 694316 370148 694380
rect 395844 694452 395908 694516
rect 389404 694316 389468 694380
rect 427676 694452 427740 694516
rect 427860 694452 427924 694516
rect 437244 694452 437308 694516
rect 437428 694452 437492 694516
rect 446996 694452 447060 694516
rect 447180 694452 447244 694516
rect 476068 694452 476132 694516
rect 417556 694316 417620 694380
rect 417740 694316 417804 694380
rect 410564 694180 410628 694244
rect 414980 694180 415044 694244
rect 418476 694316 418540 694380
rect 439452 694316 439516 694380
rect 451228 694316 451292 694380
rect 475884 694316 475948 694380
rect 379284 694044 379348 694108
rect 379836 694044 379900 694108
rect 398604 694044 398668 694108
rect 399156 694044 399220 694108
rect 417740 694044 417804 694108
rect 476068 694180 476132 694244
rect 427676 694044 427740 694108
rect 427860 694044 427924 694108
rect 437244 694044 437308 694108
rect 437428 694044 437492 694108
rect 446996 694044 447060 694108
rect 451412 694044 451476 694108
rect 475884 694044 475948 694108
rect 505692 694316 505756 694380
rect 521700 694452 521764 694516
rect 492628 694180 492692 694244
rect 543596 694316 543660 694380
rect 521700 694180 521764 694244
rect 531268 694180 531332 694244
rect 543780 694180 543844 694244
rect 562916 694316 562980 694380
rect 568620 694316 568684 694380
rect 563100 694180 563164 694244
rect 568620 694180 568684 694244
rect 529244 694044 529308 694108
rect 538812 694044 538876 694108
rect 548564 694044 548628 694108
rect 410564 693908 410628 693972
rect 29132 693772 29196 693836
rect 37228 693772 37292 693836
rect 71820 693772 71884 693836
rect 231900 693772 231964 693836
rect 232636 693772 232700 693836
rect 251220 693772 251284 693836
rect 251956 693772 252020 693836
rect 415164 693908 415228 693972
rect 102732 693636 102796 693700
rect 103284 693636 103348 693700
rect 232084 693636 232148 693700
rect 235948 693636 236012 693700
rect 251404 693636 251468 693700
rect 255268 693636 255332 693700
rect 270908 693636 270972 693700
rect 271276 693636 271340 693700
rect 414428 693636 414492 693700
rect 415164 693636 415228 693700
rect 521332 693636 521396 693700
rect 529244 693636 529308 693700
rect 538812 693636 538876 693700
rect 548564 693636 548628 693700
rect 18832 6012 18896 6016
rect 18832 5956 18836 6012
rect 18836 5956 18892 6012
rect 18892 5956 18896 6012
rect 18832 5952 18896 5956
rect 18912 6012 18976 6016
rect 18912 5956 18916 6012
rect 18916 5956 18972 6012
rect 18972 5956 18976 6012
rect 18912 5952 18976 5956
rect 18992 6012 19056 6016
rect 18992 5956 18996 6012
rect 18996 5956 19052 6012
rect 19052 5956 19056 6012
rect 18992 5952 19056 5956
rect 19072 6012 19136 6016
rect 19072 5956 19076 6012
rect 19076 5956 19132 6012
rect 19132 5956 19136 6012
rect 19072 5952 19136 5956
rect 19152 6012 19216 6016
rect 19152 5956 19156 6012
rect 19156 5956 19212 6012
rect 19212 5956 19216 6012
rect 19152 5952 19216 5956
rect 19232 6012 19296 6016
rect 19232 5956 19236 6012
rect 19236 5956 19292 6012
rect 19292 5956 19296 6012
rect 19232 5952 19296 5956
rect 19312 6012 19376 6016
rect 19312 5956 19316 6012
rect 19316 5956 19372 6012
rect 19372 5956 19376 6012
rect 19312 5952 19376 5956
rect 54832 6012 54896 6016
rect 54832 5956 54836 6012
rect 54836 5956 54892 6012
rect 54892 5956 54896 6012
rect 54832 5952 54896 5956
rect 54912 6012 54976 6016
rect 54912 5956 54916 6012
rect 54916 5956 54972 6012
rect 54972 5956 54976 6012
rect 54912 5952 54976 5956
rect 54992 6012 55056 6016
rect 54992 5956 54996 6012
rect 54996 5956 55052 6012
rect 55052 5956 55056 6012
rect 54992 5952 55056 5956
rect 55072 6012 55136 6016
rect 55072 5956 55076 6012
rect 55076 5956 55132 6012
rect 55132 5956 55136 6012
rect 55072 5952 55136 5956
rect 55152 6012 55216 6016
rect 55152 5956 55156 6012
rect 55156 5956 55212 6012
rect 55212 5956 55216 6012
rect 55152 5952 55216 5956
rect 55232 6012 55296 6016
rect 55232 5956 55236 6012
rect 55236 5956 55292 6012
rect 55292 5956 55296 6012
rect 55232 5952 55296 5956
rect 55312 6012 55376 6016
rect 55312 5956 55316 6012
rect 55316 5956 55372 6012
rect 55372 5956 55376 6012
rect 55312 5952 55376 5956
rect 90832 6012 90896 6016
rect 90832 5956 90836 6012
rect 90836 5956 90892 6012
rect 90892 5956 90896 6012
rect 90832 5952 90896 5956
rect 90912 6012 90976 6016
rect 90912 5956 90916 6012
rect 90916 5956 90972 6012
rect 90972 5956 90976 6012
rect 90912 5952 90976 5956
rect 90992 6012 91056 6016
rect 90992 5956 90996 6012
rect 90996 5956 91052 6012
rect 91052 5956 91056 6012
rect 90992 5952 91056 5956
rect 91072 6012 91136 6016
rect 91072 5956 91076 6012
rect 91076 5956 91132 6012
rect 91132 5956 91136 6012
rect 91072 5952 91136 5956
rect 91152 6012 91216 6016
rect 91152 5956 91156 6012
rect 91156 5956 91212 6012
rect 91212 5956 91216 6012
rect 91152 5952 91216 5956
rect 91232 6012 91296 6016
rect 91232 5956 91236 6012
rect 91236 5956 91292 6012
rect 91292 5956 91296 6012
rect 91232 5952 91296 5956
rect 91312 6012 91376 6016
rect 91312 5956 91316 6012
rect 91316 5956 91372 6012
rect 91372 5956 91376 6012
rect 91312 5952 91376 5956
rect 126832 6012 126896 6016
rect 126832 5956 126836 6012
rect 126836 5956 126892 6012
rect 126892 5956 126896 6012
rect 126832 5952 126896 5956
rect 126912 6012 126976 6016
rect 126912 5956 126916 6012
rect 126916 5956 126972 6012
rect 126972 5956 126976 6012
rect 126912 5952 126976 5956
rect 126992 6012 127056 6016
rect 126992 5956 126996 6012
rect 126996 5956 127052 6012
rect 127052 5956 127056 6012
rect 126992 5952 127056 5956
rect 127072 6012 127136 6016
rect 127072 5956 127076 6012
rect 127076 5956 127132 6012
rect 127132 5956 127136 6012
rect 127072 5952 127136 5956
rect 127152 6012 127216 6016
rect 127152 5956 127156 6012
rect 127156 5956 127212 6012
rect 127212 5956 127216 6012
rect 127152 5952 127216 5956
rect 127232 6012 127296 6016
rect 127232 5956 127236 6012
rect 127236 5956 127292 6012
rect 127292 5956 127296 6012
rect 127232 5952 127296 5956
rect 127312 6012 127376 6016
rect 127312 5956 127316 6012
rect 127316 5956 127372 6012
rect 127372 5956 127376 6012
rect 127312 5952 127376 5956
rect 162832 6012 162896 6016
rect 162832 5956 162836 6012
rect 162836 5956 162892 6012
rect 162892 5956 162896 6012
rect 162832 5952 162896 5956
rect 162912 6012 162976 6016
rect 162912 5956 162916 6012
rect 162916 5956 162972 6012
rect 162972 5956 162976 6012
rect 162912 5952 162976 5956
rect 162992 6012 163056 6016
rect 162992 5956 162996 6012
rect 162996 5956 163052 6012
rect 163052 5956 163056 6012
rect 162992 5952 163056 5956
rect 163072 6012 163136 6016
rect 163072 5956 163076 6012
rect 163076 5956 163132 6012
rect 163132 5956 163136 6012
rect 163072 5952 163136 5956
rect 163152 6012 163216 6016
rect 163152 5956 163156 6012
rect 163156 5956 163212 6012
rect 163212 5956 163216 6012
rect 163152 5952 163216 5956
rect 163232 6012 163296 6016
rect 163232 5956 163236 6012
rect 163236 5956 163292 6012
rect 163292 5956 163296 6012
rect 163232 5952 163296 5956
rect 163312 6012 163376 6016
rect 163312 5956 163316 6012
rect 163316 5956 163372 6012
rect 163372 5956 163376 6012
rect 163312 5952 163376 5956
rect 198832 6012 198896 6016
rect 198832 5956 198836 6012
rect 198836 5956 198892 6012
rect 198892 5956 198896 6012
rect 198832 5952 198896 5956
rect 198912 6012 198976 6016
rect 198912 5956 198916 6012
rect 198916 5956 198972 6012
rect 198972 5956 198976 6012
rect 198912 5952 198976 5956
rect 198992 6012 199056 6016
rect 198992 5956 198996 6012
rect 198996 5956 199052 6012
rect 199052 5956 199056 6012
rect 198992 5952 199056 5956
rect 199072 6012 199136 6016
rect 199072 5956 199076 6012
rect 199076 5956 199132 6012
rect 199132 5956 199136 6012
rect 199072 5952 199136 5956
rect 199152 6012 199216 6016
rect 199152 5956 199156 6012
rect 199156 5956 199212 6012
rect 199212 5956 199216 6012
rect 199152 5952 199216 5956
rect 199232 6012 199296 6016
rect 199232 5956 199236 6012
rect 199236 5956 199292 6012
rect 199292 5956 199296 6012
rect 199232 5952 199296 5956
rect 199312 6012 199376 6016
rect 199312 5956 199316 6012
rect 199316 5956 199372 6012
rect 199372 5956 199376 6012
rect 199312 5952 199376 5956
rect 234832 6012 234896 6016
rect 234832 5956 234836 6012
rect 234836 5956 234892 6012
rect 234892 5956 234896 6012
rect 234832 5952 234896 5956
rect 234912 6012 234976 6016
rect 234912 5956 234916 6012
rect 234916 5956 234972 6012
rect 234972 5956 234976 6012
rect 234912 5952 234976 5956
rect 234992 6012 235056 6016
rect 234992 5956 234996 6012
rect 234996 5956 235052 6012
rect 235052 5956 235056 6012
rect 234992 5952 235056 5956
rect 235072 6012 235136 6016
rect 235072 5956 235076 6012
rect 235076 5956 235132 6012
rect 235132 5956 235136 6012
rect 235072 5952 235136 5956
rect 235152 6012 235216 6016
rect 235152 5956 235156 6012
rect 235156 5956 235212 6012
rect 235212 5956 235216 6012
rect 235152 5952 235216 5956
rect 235232 6012 235296 6016
rect 235232 5956 235236 6012
rect 235236 5956 235292 6012
rect 235292 5956 235296 6012
rect 235232 5952 235296 5956
rect 235312 6012 235376 6016
rect 235312 5956 235316 6012
rect 235316 5956 235372 6012
rect 235372 5956 235376 6012
rect 235312 5952 235376 5956
rect 270832 6012 270896 6016
rect 270832 5956 270836 6012
rect 270836 5956 270892 6012
rect 270892 5956 270896 6012
rect 270832 5952 270896 5956
rect 270912 6012 270976 6016
rect 270912 5956 270916 6012
rect 270916 5956 270972 6012
rect 270972 5956 270976 6012
rect 270912 5952 270976 5956
rect 270992 6012 271056 6016
rect 270992 5956 270996 6012
rect 270996 5956 271052 6012
rect 271052 5956 271056 6012
rect 270992 5952 271056 5956
rect 271072 6012 271136 6016
rect 271072 5956 271076 6012
rect 271076 5956 271132 6012
rect 271132 5956 271136 6012
rect 271072 5952 271136 5956
rect 271152 6012 271216 6016
rect 271152 5956 271156 6012
rect 271156 5956 271212 6012
rect 271212 5956 271216 6012
rect 271152 5952 271216 5956
rect 271232 6012 271296 6016
rect 271232 5956 271236 6012
rect 271236 5956 271292 6012
rect 271292 5956 271296 6012
rect 271232 5952 271296 5956
rect 271312 6012 271376 6016
rect 271312 5956 271316 6012
rect 271316 5956 271372 6012
rect 271372 5956 271376 6012
rect 271312 5952 271376 5956
rect 306832 6012 306896 6016
rect 306832 5956 306836 6012
rect 306836 5956 306892 6012
rect 306892 5956 306896 6012
rect 306832 5952 306896 5956
rect 306912 6012 306976 6016
rect 306912 5956 306916 6012
rect 306916 5956 306972 6012
rect 306972 5956 306976 6012
rect 306912 5952 306976 5956
rect 306992 6012 307056 6016
rect 306992 5956 306996 6012
rect 306996 5956 307052 6012
rect 307052 5956 307056 6012
rect 306992 5952 307056 5956
rect 307072 6012 307136 6016
rect 307072 5956 307076 6012
rect 307076 5956 307132 6012
rect 307132 5956 307136 6012
rect 307072 5952 307136 5956
rect 307152 6012 307216 6016
rect 307152 5956 307156 6012
rect 307156 5956 307212 6012
rect 307212 5956 307216 6012
rect 307152 5952 307216 5956
rect 307232 6012 307296 6016
rect 307232 5956 307236 6012
rect 307236 5956 307292 6012
rect 307292 5956 307296 6012
rect 307232 5952 307296 5956
rect 307312 6012 307376 6016
rect 307312 5956 307316 6012
rect 307316 5956 307372 6012
rect 307372 5956 307376 6012
rect 307312 5952 307376 5956
rect 342832 6012 342896 6016
rect 342832 5956 342836 6012
rect 342836 5956 342892 6012
rect 342892 5956 342896 6012
rect 342832 5952 342896 5956
rect 342912 6012 342976 6016
rect 342912 5956 342916 6012
rect 342916 5956 342972 6012
rect 342972 5956 342976 6012
rect 342912 5952 342976 5956
rect 342992 6012 343056 6016
rect 342992 5956 342996 6012
rect 342996 5956 343052 6012
rect 343052 5956 343056 6012
rect 342992 5952 343056 5956
rect 343072 6012 343136 6016
rect 343072 5956 343076 6012
rect 343076 5956 343132 6012
rect 343132 5956 343136 6012
rect 343072 5952 343136 5956
rect 343152 6012 343216 6016
rect 343152 5956 343156 6012
rect 343156 5956 343212 6012
rect 343212 5956 343216 6012
rect 343152 5952 343216 5956
rect 343232 6012 343296 6016
rect 343232 5956 343236 6012
rect 343236 5956 343292 6012
rect 343292 5956 343296 6012
rect 343232 5952 343296 5956
rect 343312 6012 343376 6016
rect 343312 5956 343316 6012
rect 343316 5956 343372 6012
rect 343372 5956 343376 6012
rect 343312 5952 343376 5956
rect 378832 6012 378896 6016
rect 378832 5956 378836 6012
rect 378836 5956 378892 6012
rect 378892 5956 378896 6012
rect 378832 5952 378896 5956
rect 378912 6012 378976 6016
rect 378912 5956 378916 6012
rect 378916 5956 378972 6012
rect 378972 5956 378976 6012
rect 378912 5952 378976 5956
rect 378992 6012 379056 6016
rect 378992 5956 378996 6012
rect 378996 5956 379052 6012
rect 379052 5956 379056 6012
rect 378992 5952 379056 5956
rect 379072 6012 379136 6016
rect 379072 5956 379076 6012
rect 379076 5956 379132 6012
rect 379132 5956 379136 6012
rect 379072 5952 379136 5956
rect 379152 6012 379216 6016
rect 379152 5956 379156 6012
rect 379156 5956 379212 6012
rect 379212 5956 379216 6012
rect 379152 5952 379216 5956
rect 379232 6012 379296 6016
rect 379232 5956 379236 6012
rect 379236 5956 379292 6012
rect 379292 5956 379296 6012
rect 379232 5952 379296 5956
rect 379312 6012 379376 6016
rect 379312 5956 379316 6012
rect 379316 5956 379372 6012
rect 379372 5956 379376 6012
rect 379312 5952 379376 5956
rect 414832 6012 414896 6016
rect 414832 5956 414836 6012
rect 414836 5956 414892 6012
rect 414892 5956 414896 6012
rect 414832 5952 414896 5956
rect 414912 6012 414976 6016
rect 414912 5956 414916 6012
rect 414916 5956 414972 6012
rect 414972 5956 414976 6012
rect 414912 5952 414976 5956
rect 414992 6012 415056 6016
rect 414992 5956 414996 6012
rect 414996 5956 415052 6012
rect 415052 5956 415056 6012
rect 414992 5952 415056 5956
rect 415072 6012 415136 6016
rect 415072 5956 415076 6012
rect 415076 5956 415132 6012
rect 415132 5956 415136 6012
rect 415072 5952 415136 5956
rect 415152 6012 415216 6016
rect 415152 5956 415156 6012
rect 415156 5956 415212 6012
rect 415212 5956 415216 6012
rect 415152 5952 415216 5956
rect 415232 6012 415296 6016
rect 415232 5956 415236 6012
rect 415236 5956 415292 6012
rect 415292 5956 415296 6012
rect 415232 5952 415296 5956
rect 415312 6012 415376 6016
rect 415312 5956 415316 6012
rect 415316 5956 415372 6012
rect 415372 5956 415376 6012
rect 415312 5952 415376 5956
rect 450832 6012 450896 6016
rect 450832 5956 450836 6012
rect 450836 5956 450892 6012
rect 450892 5956 450896 6012
rect 450832 5952 450896 5956
rect 450912 6012 450976 6016
rect 450912 5956 450916 6012
rect 450916 5956 450972 6012
rect 450972 5956 450976 6012
rect 450912 5952 450976 5956
rect 450992 6012 451056 6016
rect 450992 5956 450996 6012
rect 450996 5956 451052 6012
rect 451052 5956 451056 6012
rect 450992 5952 451056 5956
rect 451072 6012 451136 6016
rect 451072 5956 451076 6012
rect 451076 5956 451132 6012
rect 451132 5956 451136 6012
rect 451072 5952 451136 5956
rect 451152 6012 451216 6016
rect 451152 5956 451156 6012
rect 451156 5956 451212 6012
rect 451212 5956 451216 6012
rect 451152 5952 451216 5956
rect 451232 6012 451296 6016
rect 451232 5956 451236 6012
rect 451236 5956 451292 6012
rect 451292 5956 451296 6012
rect 451232 5952 451296 5956
rect 451312 6012 451376 6016
rect 451312 5956 451316 6012
rect 451316 5956 451372 6012
rect 451372 5956 451376 6012
rect 451312 5952 451376 5956
rect 486832 6012 486896 6016
rect 486832 5956 486836 6012
rect 486836 5956 486892 6012
rect 486892 5956 486896 6012
rect 486832 5952 486896 5956
rect 486912 6012 486976 6016
rect 486912 5956 486916 6012
rect 486916 5956 486972 6012
rect 486972 5956 486976 6012
rect 486912 5952 486976 5956
rect 486992 6012 487056 6016
rect 486992 5956 486996 6012
rect 486996 5956 487052 6012
rect 487052 5956 487056 6012
rect 486992 5952 487056 5956
rect 487072 6012 487136 6016
rect 487072 5956 487076 6012
rect 487076 5956 487132 6012
rect 487132 5956 487136 6012
rect 487072 5952 487136 5956
rect 487152 6012 487216 6016
rect 487152 5956 487156 6012
rect 487156 5956 487212 6012
rect 487212 5956 487216 6012
rect 487152 5952 487216 5956
rect 487232 6012 487296 6016
rect 487232 5956 487236 6012
rect 487236 5956 487292 6012
rect 487292 5956 487296 6012
rect 487232 5952 487296 5956
rect 487312 6012 487376 6016
rect 487312 5956 487316 6012
rect 487316 5956 487372 6012
rect 487372 5956 487376 6012
rect 487312 5952 487376 5956
rect 522832 6012 522896 6016
rect 522832 5956 522836 6012
rect 522836 5956 522892 6012
rect 522892 5956 522896 6012
rect 522832 5952 522896 5956
rect 522912 6012 522976 6016
rect 522912 5956 522916 6012
rect 522916 5956 522972 6012
rect 522972 5956 522976 6012
rect 522912 5952 522976 5956
rect 522992 6012 523056 6016
rect 522992 5956 522996 6012
rect 522996 5956 523052 6012
rect 523052 5956 523056 6012
rect 522992 5952 523056 5956
rect 523072 6012 523136 6016
rect 523072 5956 523076 6012
rect 523076 5956 523132 6012
rect 523132 5956 523136 6012
rect 523072 5952 523136 5956
rect 523152 6012 523216 6016
rect 523152 5956 523156 6012
rect 523156 5956 523212 6012
rect 523212 5956 523216 6012
rect 523152 5952 523216 5956
rect 523232 6012 523296 6016
rect 523232 5956 523236 6012
rect 523236 5956 523292 6012
rect 523292 5956 523296 6012
rect 523232 5952 523296 5956
rect 523312 6012 523376 6016
rect 523312 5956 523316 6012
rect 523316 5956 523372 6012
rect 523372 5956 523376 6012
rect 523312 5952 523376 5956
rect 558832 6012 558896 6016
rect 558832 5956 558836 6012
rect 558836 5956 558892 6012
rect 558892 5956 558896 6012
rect 558832 5952 558896 5956
rect 558912 6012 558976 6016
rect 558912 5956 558916 6012
rect 558916 5956 558972 6012
rect 558972 5956 558976 6012
rect 558912 5952 558976 5956
rect 558992 6012 559056 6016
rect 558992 5956 558996 6012
rect 558996 5956 559052 6012
rect 559052 5956 559056 6012
rect 558992 5952 559056 5956
rect 559072 6012 559136 6016
rect 559072 5956 559076 6012
rect 559076 5956 559132 6012
rect 559132 5956 559136 6012
rect 559072 5952 559136 5956
rect 559152 6012 559216 6016
rect 559152 5956 559156 6012
rect 559156 5956 559212 6012
rect 559212 5956 559216 6012
rect 559152 5952 559216 5956
rect 559232 6012 559296 6016
rect 559232 5956 559236 6012
rect 559236 5956 559292 6012
rect 559292 5956 559296 6012
rect 559232 5952 559296 5956
rect 559312 6012 559376 6016
rect 559312 5956 559316 6012
rect 559316 5956 559372 6012
rect 559372 5956 559376 6012
rect 559312 5952 559376 5956
rect 36832 5468 36896 5472
rect 36832 5412 36836 5468
rect 36836 5412 36892 5468
rect 36892 5412 36896 5468
rect 36832 5408 36896 5412
rect 36912 5468 36976 5472
rect 36912 5412 36916 5468
rect 36916 5412 36972 5468
rect 36972 5412 36976 5468
rect 36912 5408 36976 5412
rect 36992 5468 37056 5472
rect 36992 5412 36996 5468
rect 36996 5412 37052 5468
rect 37052 5412 37056 5468
rect 36992 5408 37056 5412
rect 37072 5468 37136 5472
rect 37072 5412 37076 5468
rect 37076 5412 37132 5468
rect 37132 5412 37136 5468
rect 37072 5408 37136 5412
rect 37152 5468 37216 5472
rect 37152 5412 37156 5468
rect 37156 5412 37212 5468
rect 37212 5412 37216 5468
rect 37152 5408 37216 5412
rect 37232 5468 37296 5472
rect 37232 5412 37236 5468
rect 37236 5412 37292 5468
rect 37292 5412 37296 5468
rect 37232 5408 37296 5412
rect 37312 5468 37376 5472
rect 37312 5412 37316 5468
rect 37316 5412 37372 5468
rect 37372 5412 37376 5468
rect 37312 5408 37376 5412
rect 72832 5468 72896 5472
rect 72832 5412 72836 5468
rect 72836 5412 72892 5468
rect 72892 5412 72896 5468
rect 72832 5408 72896 5412
rect 72912 5468 72976 5472
rect 72912 5412 72916 5468
rect 72916 5412 72972 5468
rect 72972 5412 72976 5468
rect 72912 5408 72976 5412
rect 72992 5468 73056 5472
rect 72992 5412 72996 5468
rect 72996 5412 73052 5468
rect 73052 5412 73056 5468
rect 72992 5408 73056 5412
rect 73072 5468 73136 5472
rect 73072 5412 73076 5468
rect 73076 5412 73132 5468
rect 73132 5412 73136 5468
rect 73072 5408 73136 5412
rect 73152 5468 73216 5472
rect 73152 5412 73156 5468
rect 73156 5412 73212 5468
rect 73212 5412 73216 5468
rect 73152 5408 73216 5412
rect 73232 5468 73296 5472
rect 73232 5412 73236 5468
rect 73236 5412 73292 5468
rect 73292 5412 73296 5468
rect 73232 5408 73296 5412
rect 73312 5468 73376 5472
rect 73312 5412 73316 5468
rect 73316 5412 73372 5468
rect 73372 5412 73376 5468
rect 73312 5408 73376 5412
rect 108832 5468 108896 5472
rect 108832 5412 108836 5468
rect 108836 5412 108892 5468
rect 108892 5412 108896 5468
rect 108832 5408 108896 5412
rect 108912 5468 108976 5472
rect 108912 5412 108916 5468
rect 108916 5412 108972 5468
rect 108972 5412 108976 5468
rect 108912 5408 108976 5412
rect 108992 5468 109056 5472
rect 108992 5412 108996 5468
rect 108996 5412 109052 5468
rect 109052 5412 109056 5468
rect 108992 5408 109056 5412
rect 109072 5468 109136 5472
rect 109072 5412 109076 5468
rect 109076 5412 109132 5468
rect 109132 5412 109136 5468
rect 109072 5408 109136 5412
rect 109152 5468 109216 5472
rect 109152 5412 109156 5468
rect 109156 5412 109212 5468
rect 109212 5412 109216 5468
rect 109152 5408 109216 5412
rect 109232 5468 109296 5472
rect 109232 5412 109236 5468
rect 109236 5412 109292 5468
rect 109292 5412 109296 5468
rect 109232 5408 109296 5412
rect 109312 5468 109376 5472
rect 109312 5412 109316 5468
rect 109316 5412 109372 5468
rect 109372 5412 109376 5468
rect 109312 5408 109376 5412
rect 144832 5468 144896 5472
rect 144832 5412 144836 5468
rect 144836 5412 144892 5468
rect 144892 5412 144896 5468
rect 144832 5408 144896 5412
rect 144912 5468 144976 5472
rect 144912 5412 144916 5468
rect 144916 5412 144972 5468
rect 144972 5412 144976 5468
rect 144912 5408 144976 5412
rect 144992 5468 145056 5472
rect 144992 5412 144996 5468
rect 144996 5412 145052 5468
rect 145052 5412 145056 5468
rect 144992 5408 145056 5412
rect 145072 5468 145136 5472
rect 145072 5412 145076 5468
rect 145076 5412 145132 5468
rect 145132 5412 145136 5468
rect 145072 5408 145136 5412
rect 145152 5468 145216 5472
rect 145152 5412 145156 5468
rect 145156 5412 145212 5468
rect 145212 5412 145216 5468
rect 145152 5408 145216 5412
rect 145232 5468 145296 5472
rect 145232 5412 145236 5468
rect 145236 5412 145292 5468
rect 145292 5412 145296 5468
rect 145232 5408 145296 5412
rect 145312 5468 145376 5472
rect 145312 5412 145316 5468
rect 145316 5412 145372 5468
rect 145372 5412 145376 5468
rect 145312 5408 145376 5412
rect 180832 5468 180896 5472
rect 180832 5412 180836 5468
rect 180836 5412 180892 5468
rect 180892 5412 180896 5468
rect 180832 5408 180896 5412
rect 180912 5468 180976 5472
rect 180912 5412 180916 5468
rect 180916 5412 180972 5468
rect 180972 5412 180976 5468
rect 180912 5408 180976 5412
rect 180992 5468 181056 5472
rect 180992 5412 180996 5468
rect 180996 5412 181052 5468
rect 181052 5412 181056 5468
rect 180992 5408 181056 5412
rect 181072 5468 181136 5472
rect 181072 5412 181076 5468
rect 181076 5412 181132 5468
rect 181132 5412 181136 5468
rect 181072 5408 181136 5412
rect 181152 5468 181216 5472
rect 181152 5412 181156 5468
rect 181156 5412 181212 5468
rect 181212 5412 181216 5468
rect 181152 5408 181216 5412
rect 181232 5468 181296 5472
rect 181232 5412 181236 5468
rect 181236 5412 181292 5468
rect 181292 5412 181296 5468
rect 181232 5408 181296 5412
rect 181312 5468 181376 5472
rect 181312 5412 181316 5468
rect 181316 5412 181372 5468
rect 181372 5412 181376 5468
rect 181312 5408 181376 5412
rect 216832 5468 216896 5472
rect 216832 5412 216836 5468
rect 216836 5412 216892 5468
rect 216892 5412 216896 5468
rect 216832 5408 216896 5412
rect 216912 5468 216976 5472
rect 216912 5412 216916 5468
rect 216916 5412 216972 5468
rect 216972 5412 216976 5468
rect 216912 5408 216976 5412
rect 216992 5468 217056 5472
rect 216992 5412 216996 5468
rect 216996 5412 217052 5468
rect 217052 5412 217056 5468
rect 216992 5408 217056 5412
rect 217072 5468 217136 5472
rect 217072 5412 217076 5468
rect 217076 5412 217132 5468
rect 217132 5412 217136 5468
rect 217072 5408 217136 5412
rect 217152 5468 217216 5472
rect 217152 5412 217156 5468
rect 217156 5412 217212 5468
rect 217212 5412 217216 5468
rect 217152 5408 217216 5412
rect 217232 5468 217296 5472
rect 217232 5412 217236 5468
rect 217236 5412 217292 5468
rect 217292 5412 217296 5468
rect 217232 5408 217296 5412
rect 217312 5468 217376 5472
rect 217312 5412 217316 5468
rect 217316 5412 217372 5468
rect 217372 5412 217376 5468
rect 217312 5408 217376 5412
rect 252832 5468 252896 5472
rect 252832 5412 252836 5468
rect 252836 5412 252892 5468
rect 252892 5412 252896 5468
rect 252832 5408 252896 5412
rect 252912 5468 252976 5472
rect 252912 5412 252916 5468
rect 252916 5412 252972 5468
rect 252972 5412 252976 5468
rect 252912 5408 252976 5412
rect 252992 5468 253056 5472
rect 252992 5412 252996 5468
rect 252996 5412 253052 5468
rect 253052 5412 253056 5468
rect 252992 5408 253056 5412
rect 253072 5468 253136 5472
rect 253072 5412 253076 5468
rect 253076 5412 253132 5468
rect 253132 5412 253136 5468
rect 253072 5408 253136 5412
rect 253152 5468 253216 5472
rect 253152 5412 253156 5468
rect 253156 5412 253212 5468
rect 253212 5412 253216 5468
rect 253152 5408 253216 5412
rect 253232 5468 253296 5472
rect 253232 5412 253236 5468
rect 253236 5412 253292 5468
rect 253292 5412 253296 5468
rect 253232 5408 253296 5412
rect 253312 5468 253376 5472
rect 253312 5412 253316 5468
rect 253316 5412 253372 5468
rect 253372 5412 253376 5468
rect 253312 5408 253376 5412
rect 288832 5468 288896 5472
rect 288832 5412 288836 5468
rect 288836 5412 288892 5468
rect 288892 5412 288896 5468
rect 288832 5408 288896 5412
rect 288912 5468 288976 5472
rect 288912 5412 288916 5468
rect 288916 5412 288972 5468
rect 288972 5412 288976 5468
rect 288912 5408 288976 5412
rect 288992 5468 289056 5472
rect 288992 5412 288996 5468
rect 288996 5412 289052 5468
rect 289052 5412 289056 5468
rect 288992 5408 289056 5412
rect 289072 5468 289136 5472
rect 289072 5412 289076 5468
rect 289076 5412 289132 5468
rect 289132 5412 289136 5468
rect 289072 5408 289136 5412
rect 289152 5468 289216 5472
rect 289152 5412 289156 5468
rect 289156 5412 289212 5468
rect 289212 5412 289216 5468
rect 289152 5408 289216 5412
rect 289232 5468 289296 5472
rect 289232 5412 289236 5468
rect 289236 5412 289292 5468
rect 289292 5412 289296 5468
rect 289232 5408 289296 5412
rect 289312 5468 289376 5472
rect 289312 5412 289316 5468
rect 289316 5412 289372 5468
rect 289372 5412 289376 5468
rect 289312 5408 289376 5412
rect 324832 5468 324896 5472
rect 324832 5412 324836 5468
rect 324836 5412 324892 5468
rect 324892 5412 324896 5468
rect 324832 5408 324896 5412
rect 324912 5468 324976 5472
rect 324912 5412 324916 5468
rect 324916 5412 324972 5468
rect 324972 5412 324976 5468
rect 324912 5408 324976 5412
rect 324992 5468 325056 5472
rect 324992 5412 324996 5468
rect 324996 5412 325052 5468
rect 325052 5412 325056 5468
rect 324992 5408 325056 5412
rect 325072 5468 325136 5472
rect 325072 5412 325076 5468
rect 325076 5412 325132 5468
rect 325132 5412 325136 5468
rect 325072 5408 325136 5412
rect 325152 5468 325216 5472
rect 325152 5412 325156 5468
rect 325156 5412 325212 5468
rect 325212 5412 325216 5468
rect 325152 5408 325216 5412
rect 325232 5468 325296 5472
rect 325232 5412 325236 5468
rect 325236 5412 325292 5468
rect 325292 5412 325296 5468
rect 325232 5408 325296 5412
rect 325312 5468 325376 5472
rect 325312 5412 325316 5468
rect 325316 5412 325372 5468
rect 325372 5412 325376 5468
rect 325312 5408 325376 5412
rect 360832 5468 360896 5472
rect 360832 5412 360836 5468
rect 360836 5412 360892 5468
rect 360892 5412 360896 5468
rect 360832 5408 360896 5412
rect 360912 5468 360976 5472
rect 360912 5412 360916 5468
rect 360916 5412 360972 5468
rect 360972 5412 360976 5468
rect 360912 5408 360976 5412
rect 360992 5468 361056 5472
rect 360992 5412 360996 5468
rect 360996 5412 361052 5468
rect 361052 5412 361056 5468
rect 360992 5408 361056 5412
rect 361072 5468 361136 5472
rect 361072 5412 361076 5468
rect 361076 5412 361132 5468
rect 361132 5412 361136 5468
rect 361072 5408 361136 5412
rect 361152 5468 361216 5472
rect 361152 5412 361156 5468
rect 361156 5412 361212 5468
rect 361212 5412 361216 5468
rect 361152 5408 361216 5412
rect 361232 5468 361296 5472
rect 361232 5412 361236 5468
rect 361236 5412 361292 5468
rect 361292 5412 361296 5468
rect 361232 5408 361296 5412
rect 361312 5468 361376 5472
rect 361312 5412 361316 5468
rect 361316 5412 361372 5468
rect 361372 5412 361376 5468
rect 361312 5408 361376 5412
rect 396832 5468 396896 5472
rect 396832 5412 396836 5468
rect 396836 5412 396892 5468
rect 396892 5412 396896 5468
rect 396832 5408 396896 5412
rect 396912 5468 396976 5472
rect 396912 5412 396916 5468
rect 396916 5412 396972 5468
rect 396972 5412 396976 5468
rect 396912 5408 396976 5412
rect 396992 5468 397056 5472
rect 396992 5412 396996 5468
rect 396996 5412 397052 5468
rect 397052 5412 397056 5468
rect 396992 5408 397056 5412
rect 397072 5468 397136 5472
rect 397072 5412 397076 5468
rect 397076 5412 397132 5468
rect 397132 5412 397136 5468
rect 397072 5408 397136 5412
rect 397152 5468 397216 5472
rect 397152 5412 397156 5468
rect 397156 5412 397212 5468
rect 397212 5412 397216 5468
rect 397152 5408 397216 5412
rect 397232 5468 397296 5472
rect 397232 5412 397236 5468
rect 397236 5412 397292 5468
rect 397292 5412 397296 5468
rect 397232 5408 397296 5412
rect 397312 5468 397376 5472
rect 397312 5412 397316 5468
rect 397316 5412 397372 5468
rect 397372 5412 397376 5468
rect 397312 5408 397376 5412
rect 432832 5468 432896 5472
rect 432832 5412 432836 5468
rect 432836 5412 432892 5468
rect 432892 5412 432896 5468
rect 432832 5408 432896 5412
rect 432912 5468 432976 5472
rect 432912 5412 432916 5468
rect 432916 5412 432972 5468
rect 432972 5412 432976 5468
rect 432912 5408 432976 5412
rect 432992 5468 433056 5472
rect 432992 5412 432996 5468
rect 432996 5412 433052 5468
rect 433052 5412 433056 5468
rect 432992 5408 433056 5412
rect 433072 5468 433136 5472
rect 433072 5412 433076 5468
rect 433076 5412 433132 5468
rect 433132 5412 433136 5468
rect 433072 5408 433136 5412
rect 433152 5468 433216 5472
rect 433152 5412 433156 5468
rect 433156 5412 433212 5468
rect 433212 5412 433216 5468
rect 433152 5408 433216 5412
rect 433232 5468 433296 5472
rect 433232 5412 433236 5468
rect 433236 5412 433292 5468
rect 433292 5412 433296 5468
rect 433232 5408 433296 5412
rect 433312 5468 433376 5472
rect 433312 5412 433316 5468
rect 433316 5412 433372 5468
rect 433372 5412 433376 5468
rect 433312 5408 433376 5412
rect 468832 5468 468896 5472
rect 468832 5412 468836 5468
rect 468836 5412 468892 5468
rect 468892 5412 468896 5468
rect 468832 5408 468896 5412
rect 468912 5468 468976 5472
rect 468912 5412 468916 5468
rect 468916 5412 468972 5468
rect 468972 5412 468976 5468
rect 468912 5408 468976 5412
rect 468992 5468 469056 5472
rect 468992 5412 468996 5468
rect 468996 5412 469052 5468
rect 469052 5412 469056 5468
rect 468992 5408 469056 5412
rect 469072 5468 469136 5472
rect 469072 5412 469076 5468
rect 469076 5412 469132 5468
rect 469132 5412 469136 5468
rect 469072 5408 469136 5412
rect 469152 5468 469216 5472
rect 469152 5412 469156 5468
rect 469156 5412 469212 5468
rect 469212 5412 469216 5468
rect 469152 5408 469216 5412
rect 469232 5468 469296 5472
rect 469232 5412 469236 5468
rect 469236 5412 469292 5468
rect 469292 5412 469296 5468
rect 469232 5408 469296 5412
rect 469312 5468 469376 5472
rect 469312 5412 469316 5468
rect 469316 5412 469372 5468
rect 469372 5412 469376 5468
rect 469312 5408 469376 5412
rect 504832 5468 504896 5472
rect 504832 5412 504836 5468
rect 504836 5412 504892 5468
rect 504892 5412 504896 5468
rect 504832 5408 504896 5412
rect 504912 5468 504976 5472
rect 504912 5412 504916 5468
rect 504916 5412 504972 5468
rect 504972 5412 504976 5468
rect 504912 5408 504976 5412
rect 504992 5468 505056 5472
rect 504992 5412 504996 5468
rect 504996 5412 505052 5468
rect 505052 5412 505056 5468
rect 504992 5408 505056 5412
rect 505072 5468 505136 5472
rect 505072 5412 505076 5468
rect 505076 5412 505132 5468
rect 505132 5412 505136 5468
rect 505072 5408 505136 5412
rect 505152 5468 505216 5472
rect 505152 5412 505156 5468
rect 505156 5412 505212 5468
rect 505212 5412 505216 5468
rect 505152 5408 505216 5412
rect 505232 5468 505296 5472
rect 505232 5412 505236 5468
rect 505236 5412 505292 5468
rect 505292 5412 505296 5468
rect 505232 5408 505296 5412
rect 505312 5468 505376 5472
rect 505312 5412 505316 5468
rect 505316 5412 505372 5468
rect 505372 5412 505376 5468
rect 505312 5408 505376 5412
rect 540832 5468 540896 5472
rect 540832 5412 540836 5468
rect 540836 5412 540892 5468
rect 540892 5412 540896 5468
rect 540832 5408 540896 5412
rect 540912 5468 540976 5472
rect 540912 5412 540916 5468
rect 540916 5412 540972 5468
rect 540972 5412 540976 5468
rect 540912 5408 540976 5412
rect 540992 5468 541056 5472
rect 540992 5412 540996 5468
rect 540996 5412 541052 5468
rect 541052 5412 541056 5468
rect 540992 5408 541056 5412
rect 541072 5468 541136 5472
rect 541072 5412 541076 5468
rect 541076 5412 541132 5468
rect 541132 5412 541136 5468
rect 541072 5408 541136 5412
rect 541152 5468 541216 5472
rect 541152 5412 541156 5468
rect 541156 5412 541212 5468
rect 541212 5412 541216 5468
rect 541152 5408 541216 5412
rect 541232 5468 541296 5472
rect 541232 5412 541236 5468
rect 541236 5412 541292 5468
rect 541292 5412 541296 5468
rect 541232 5408 541296 5412
rect 541312 5468 541376 5472
rect 541312 5412 541316 5468
rect 541316 5412 541372 5468
rect 541372 5412 541376 5468
rect 541312 5408 541376 5412
rect 576832 5468 576896 5472
rect 576832 5412 576836 5468
rect 576836 5412 576892 5468
rect 576892 5412 576896 5468
rect 576832 5408 576896 5412
rect 576912 5468 576976 5472
rect 576912 5412 576916 5468
rect 576916 5412 576972 5468
rect 576972 5412 576976 5468
rect 576912 5408 576976 5412
rect 576992 5468 577056 5472
rect 576992 5412 576996 5468
rect 576996 5412 577052 5468
rect 577052 5412 577056 5468
rect 576992 5408 577056 5412
rect 577072 5468 577136 5472
rect 577072 5412 577076 5468
rect 577076 5412 577132 5468
rect 577132 5412 577136 5468
rect 577072 5408 577136 5412
rect 577152 5468 577216 5472
rect 577152 5412 577156 5468
rect 577156 5412 577212 5468
rect 577212 5412 577216 5468
rect 577152 5408 577216 5412
rect 577232 5468 577296 5472
rect 577232 5412 577236 5468
rect 577236 5412 577292 5468
rect 577292 5412 577296 5468
rect 577232 5408 577296 5412
rect 577312 5468 577376 5472
rect 577312 5412 577316 5468
rect 577316 5412 577372 5468
rect 577372 5412 577376 5468
rect 577312 5408 577376 5412
rect 18832 4924 18896 4928
rect 18832 4868 18836 4924
rect 18836 4868 18892 4924
rect 18892 4868 18896 4924
rect 18832 4864 18896 4868
rect 18912 4924 18976 4928
rect 18912 4868 18916 4924
rect 18916 4868 18972 4924
rect 18972 4868 18976 4924
rect 18912 4864 18976 4868
rect 18992 4924 19056 4928
rect 18992 4868 18996 4924
rect 18996 4868 19052 4924
rect 19052 4868 19056 4924
rect 18992 4864 19056 4868
rect 19072 4924 19136 4928
rect 19072 4868 19076 4924
rect 19076 4868 19132 4924
rect 19132 4868 19136 4924
rect 19072 4864 19136 4868
rect 19152 4924 19216 4928
rect 19152 4868 19156 4924
rect 19156 4868 19212 4924
rect 19212 4868 19216 4924
rect 19152 4864 19216 4868
rect 19232 4924 19296 4928
rect 19232 4868 19236 4924
rect 19236 4868 19292 4924
rect 19292 4868 19296 4924
rect 19232 4864 19296 4868
rect 19312 4924 19376 4928
rect 19312 4868 19316 4924
rect 19316 4868 19372 4924
rect 19372 4868 19376 4924
rect 19312 4864 19376 4868
rect 54832 4924 54896 4928
rect 54832 4868 54836 4924
rect 54836 4868 54892 4924
rect 54892 4868 54896 4924
rect 54832 4864 54896 4868
rect 54912 4924 54976 4928
rect 54912 4868 54916 4924
rect 54916 4868 54972 4924
rect 54972 4868 54976 4924
rect 54912 4864 54976 4868
rect 54992 4924 55056 4928
rect 54992 4868 54996 4924
rect 54996 4868 55052 4924
rect 55052 4868 55056 4924
rect 54992 4864 55056 4868
rect 55072 4924 55136 4928
rect 55072 4868 55076 4924
rect 55076 4868 55132 4924
rect 55132 4868 55136 4924
rect 55072 4864 55136 4868
rect 55152 4924 55216 4928
rect 55152 4868 55156 4924
rect 55156 4868 55212 4924
rect 55212 4868 55216 4924
rect 55152 4864 55216 4868
rect 55232 4924 55296 4928
rect 55232 4868 55236 4924
rect 55236 4868 55292 4924
rect 55292 4868 55296 4924
rect 55232 4864 55296 4868
rect 55312 4924 55376 4928
rect 55312 4868 55316 4924
rect 55316 4868 55372 4924
rect 55372 4868 55376 4924
rect 55312 4864 55376 4868
rect 90832 4924 90896 4928
rect 90832 4868 90836 4924
rect 90836 4868 90892 4924
rect 90892 4868 90896 4924
rect 90832 4864 90896 4868
rect 90912 4924 90976 4928
rect 90912 4868 90916 4924
rect 90916 4868 90972 4924
rect 90972 4868 90976 4924
rect 90912 4864 90976 4868
rect 90992 4924 91056 4928
rect 90992 4868 90996 4924
rect 90996 4868 91052 4924
rect 91052 4868 91056 4924
rect 90992 4864 91056 4868
rect 91072 4924 91136 4928
rect 91072 4868 91076 4924
rect 91076 4868 91132 4924
rect 91132 4868 91136 4924
rect 91072 4864 91136 4868
rect 91152 4924 91216 4928
rect 91152 4868 91156 4924
rect 91156 4868 91212 4924
rect 91212 4868 91216 4924
rect 91152 4864 91216 4868
rect 91232 4924 91296 4928
rect 91232 4868 91236 4924
rect 91236 4868 91292 4924
rect 91292 4868 91296 4924
rect 91232 4864 91296 4868
rect 91312 4924 91376 4928
rect 91312 4868 91316 4924
rect 91316 4868 91372 4924
rect 91372 4868 91376 4924
rect 91312 4864 91376 4868
rect 126832 4924 126896 4928
rect 126832 4868 126836 4924
rect 126836 4868 126892 4924
rect 126892 4868 126896 4924
rect 126832 4864 126896 4868
rect 126912 4924 126976 4928
rect 126912 4868 126916 4924
rect 126916 4868 126972 4924
rect 126972 4868 126976 4924
rect 126912 4864 126976 4868
rect 126992 4924 127056 4928
rect 126992 4868 126996 4924
rect 126996 4868 127052 4924
rect 127052 4868 127056 4924
rect 126992 4864 127056 4868
rect 127072 4924 127136 4928
rect 127072 4868 127076 4924
rect 127076 4868 127132 4924
rect 127132 4868 127136 4924
rect 127072 4864 127136 4868
rect 127152 4924 127216 4928
rect 127152 4868 127156 4924
rect 127156 4868 127212 4924
rect 127212 4868 127216 4924
rect 127152 4864 127216 4868
rect 127232 4924 127296 4928
rect 127232 4868 127236 4924
rect 127236 4868 127292 4924
rect 127292 4868 127296 4924
rect 127232 4864 127296 4868
rect 127312 4924 127376 4928
rect 127312 4868 127316 4924
rect 127316 4868 127372 4924
rect 127372 4868 127376 4924
rect 127312 4864 127376 4868
rect 162832 4924 162896 4928
rect 162832 4868 162836 4924
rect 162836 4868 162892 4924
rect 162892 4868 162896 4924
rect 162832 4864 162896 4868
rect 162912 4924 162976 4928
rect 162912 4868 162916 4924
rect 162916 4868 162972 4924
rect 162972 4868 162976 4924
rect 162912 4864 162976 4868
rect 162992 4924 163056 4928
rect 162992 4868 162996 4924
rect 162996 4868 163052 4924
rect 163052 4868 163056 4924
rect 162992 4864 163056 4868
rect 163072 4924 163136 4928
rect 163072 4868 163076 4924
rect 163076 4868 163132 4924
rect 163132 4868 163136 4924
rect 163072 4864 163136 4868
rect 163152 4924 163216 4928
rect 163152 4868 163156 4924
rect 163156 4868 163212 4924
rect 163212 4868 163216 4924
rect 163152 4864 163216 4868
rect 163232 4924 163296 4928
rect 163232 4868 163236 4924
rect 163236 4868 163292 4924
rect 163292 4868 163296 4924
rect 163232 4864 163296 4868
rect 163312 4924 163376 4928
rect 163312 4868 163316 4924
rect 163316 4868 163372 4924
rect 163372 4868 163376 4924
rect 163312 4864 163376 4868
rect 198832 4924 198896 4928
rect 198832 4868 198836 4924
rect 198836 4868 198892 4924
rect 198892 4868 198896 4924
rect 198832 4864 198896 4868
rect 198912 4924 198976 4928
rect 198912 4868 198916 4924
rect 198916 4868 198972 4924
rect 198972 4868 198976 4924
rect 198912 4864 198976 4868
rect 198992 4924 199056 4928
rect 198992 4868 198996 4924
rect 198996 4868 199052 4924
rect 199052 4868 199056 4924
rect 198992 4864 199056 4868
rect 199072 4924 199136 4928
rect 199072 4868 199076 4924
rect 199076 4868 199132 4924
rect 199132 4868 199136 4924
rect 199072 4864 199136 4868
rect 199152 4924 199216 4928
rect 199152 4868 199156 4924
rect 199156 4868 199212 4924
rect 199212 4868 199216 4924
rect 199152 4864 199216 4868
rect 199232 4924 199296 4928
rect 199232 4868 199236 4924
rect 199236 4868 199292 4924
rect 199292 4868 199296 4924
rect 199232 4864 199296 4868
rect 199312 4924 199376 4928
rect 199312 4868 199316 4924
rect 199316 4868 199372 4924
rect 199372 4868 199376 4924
rect 199312 4864 199376 4868
rect 234832 4924 234896 4928
rect 234832 4868 234836 4924
rect 234836 4868 234892 4924
rect 234892 4868 234896 4924
rect 234832 4864 234896 4868
rect 234912 4924 234976 4928
rect 234912 4868 234916 4924
rect 234916 4868 234972 4924
rect 234972 4868 234976 4924
rect 234912 4864 234976 4868
rect 234992 4924 235056 4928
rect 234992 4868 234996 4924
rect 234996 4868 235052 4924
rect 235052 4868 235056 4924
rect 234992 4864 235056 4868
rect 235072 4924 235136 4928
rect 235072 4868 235076 4924
rect 235076 4868 235132 4924
rect 235132 4868 235136 4924
rect 235072 4864 235136 4868
rect 235152 4924 235216 4928
rect 235152 4868 235156 4924
rect 235156 4868 235212 4924
rect 235212 4868 235216 4924
rect 235152 4864 235216 4868
rect 235232 4924 235296 4928
rect 235232 4868 235236 4924
rect 235236 4868 235292 4924
rect 235292 4868 235296 4924
rect 235232 4864 235296 4868
rect 235312 4924 235376 4928
rect 235312 4868 235316 4924
rect 235316 4868 235372 4924
rect 235372 4868 235376 4924
rect 235312 4864 235376 4868
rect 270832 4924 270896 4928
rect 270832 4868 270836 4924
rect 270836 4868 270892 4924
rect 270892 4868 270896 4924
rect 270832 4864 270896 4868
rect 270912 4924 270976 4928
rect 270912 4868 270916 4924
rect 270916 4868 270972 4924
rect 270972 4868 270976 4924
rect 270912 4864 270976 4868
rect 270992 4924 271056 4928
rect 270992 4868 270996 4924
rect 270996 4868 271052 4924
rect 271052 4868 271056 4924
rect 270992 4864 271056 4868
rect 271072 4924 271136 4928
rect 271072 4868 271076 4924
rect 271076 4868 271132 4924
rect 271132 4868 271136 4924
rect 271072 4864 271136 4868
rect 271152 4924 271216 4928
rect 271152 4868 271156 4924
rect 271156 4868 271212 4924
rect 271212 4868 271216 4924
rect 271152 4864 271216 4868
rect 271232 4924 271296 4928
rect 271232 4868 271236 4924
rect 271236 4868 271292 4924
rect 271292 4868 271296 4924
rect 271232 4864 271296 4868
rect 271312 4924 271376 4928
rect 271312 4868 271316 4924
rect 271316 4868 271372 4924
rect 271372 4868 271376 4924
rect 271312 4864 271376 4868
rect 306832 4924 306896 4928
rect 306832 4868 306836 4924
rect 306836 4868 306892 4924
rect 306892 4868 306896 4924
rect 306832 4864 306896 4868
rect 306912 4924 306976 4928
rect 306912 4868 306916 4924
rect 306916 4868 306972 4924
rect 306972 4868 306976 4924
rect 306912 4864 306976 4868
rect 306992 4924 307056 4928
rect 306992 4868 306996 4924
rect 306996 4868 307052 4924
rect 307052 4868 307056 4924
rect 306992 4864 307056 4868
rect 307072 4924 307136 4928
rect 307072 4868 307076 4924
rect 307076 4868 307132 4924
rect 307132 4868 307136 4924
rect 307072 4864 307136 4868
rect 307152 4924 307216 4928
rect 307152 4868 307156 4924
rect 307156 4868 307212 4924
rect 307212 4868 307216 4924
rect 307152 4864 307216 4868
rect 307232 4924 307296 4928
rect 307232 4868 307236 4924
rect 307236 4868 307292 4924
rect 307292 4868 307296 4924
rect 307232 4864 307296 4868
rect 307312 4924 307376 4928
rect 307312 4868 307316 4924
rect 307316 4868 307372 4924
rect 307372 4868 307376 4924
rect 307312 4864 307376 4868
rect 342832 4924 342896 4928
rect 342832 4868 342836 4924
rect 342836 4868 342892 4924
rect 342892 4868 342896 4924
rect 342832 4864 342896 4868
rect 342912 4924 342976 4928
rect 342912 4868 342916 4924
rect 342916 4868 342972 4924
rect 342972 4868 342976 4924
rect 342912 4864 342976 4868
rect 342992 4924 343056 4928
rect 342992 4868 342996 4924
rect 342996 4868 343052 4924
rect 343052 4868 343056 4924
rect 342992 4864 343056 4868
rect 343072 4924 343136 4928
rect 343072 4868 343076 4924
rect 343076 4868 343132 4924
rect 343132 4868 343136 4924
rect 343072 4864 343136 4868
rect 343152 4924 343216 4928
rect 343152 4868 343156 4924
rect 343156 4868 343212 4924
rect 343212 4868 343216 4924
rect 343152 4864 343216 4868
rect 343232 4924 343296 4928
rect 343232 4868 343236 4924
rect 343236 4868 343292 4924
rect 343292 4868 343296 4924
rect 343232 4864 343296 4868
rect 343312 4924 343376 4928
rect 343312 4868 343316 4924
rect 343316 4868 343372 4924
rect 343372 4868 343376 4924
rect 343312 4864 343376 4868
rect 378832 4924 378896 4928
rect 378832 4868 378836 4924
rect 378836 4868 378892 4924
rect 378892 4868 378896 4924
rect 378832 4864 378896 4868
rect 378912 4924 378976 4928
rect 378912 4868 378916 4924
rect 378916 4868 378972 4924
rect 378972 4868 378976 4924
rect 378912 4864 378976 4868
rect 378992 4924 379056 4928
rect 378992 4868 378996 4924
rect 378996 4868 379052 4924
rect 379052 4868 379056 4924
rect 378992 4864 379056 4868
rect 379072 4924 379136 4928
rect 379072 4868 379076 4924
rect 379076 4868 379132 4924
rect 379132 4868 379136 4924
rect 379072 4864 379136 4868
rect 379152 4924 379216 4928
rect 379152 4868 379156 4924
rect 379156 4868 379212 4924
rect 379212 4868 379216 4924
rect 379152 4864 379216 4868
rect 379232 4924 379296 4928
rect 379232 4868 379236 4924
rect 379236 4868 379292 4924
rect 379292 4868 379296 4924
rect 379232 4864 379296 4868
rect 379312 4924 379376 4928
rect 379312 4868 379316 4924
rect 379316 4868 379372 4924
rect 379372 4868 379376 4924
rect 379312 4864 379376 4868
rect 414832 4924 414896 4928
rect 414832 4868 414836 4924
rect 414836 4868 414892 4924
rect 414892 4868 414896 4924
rect 414832 4864 414896 4868
rect 414912 4924 414976 4928
rect 414912 4868 414916 4924
rect 414916 4868 414972 4924
rect 414972 4868 414976 4924
rect 414912 4864 414976 4868
rect 414992 4924 415056 4928
rect 414992 4868 414996 4924
rect 414996 4868 415052 4924
rect 415052 4868 415056 4924
rect 414992 4864 415056 4868
rect 415072 4924 415136 4928
rect 415072 4868 415076 4924
rect 415076 4868 415132 4924
rect 415132 4868 415136 4924
rect 415072 4864 415136 4868
rect 415152 4924 415216 4928
rect 415152 4868 415156 4924
rect 415156 4868 415212 4924
rect 415212 4868 415216 4924
rect 415152 4864 415216 4868
rect 415232 4924 415296 4928
rect 415232 4868 415236 4924
rect 415236 4868 415292 4924
rect 415292 4868 415296 4924
rect 415232 4864 415296 4868
rect 415312 4924 415376 4928
rect 415312 4868 415316 4924
rect 415316 4868 415372 4924
rect 415372 4868 415376 4924
rect 415312 4864 415376 4868
rect 450832 4924 450896 4928
rect 450832 4868 450836 4924
rect 450836 4868 450892 4924
rect 450892 4868 450896 4924
rect 450832 4864 450896 4868
rect 450912 4924 450976 4928
rect 450912 4868 450916 4924
rect 450916 4868 450972 4924
rect 450972 4868 450976 4924
rect 450912 4864 450976 4868
rect 450992 4924 451056 4928
rect 450992 4868 450996 4924
rect 450996 4868 451052 4924
rect 451052 4868 451056 4924
rect 450992 4864 451056 4868
rect 451072 4924 451136 4928
rect 451072 4868 451076 4924
rect 451076 4868 451132 4924
rect 451132 4868 451136 4924
rect 451072 4864 451136 4868
rect 451152 4924 451216 4928
rect 451152 4868 451156 4924
rect 451156 4868 451212 4924
rect 451212 4868 451216 4924
rect 451152 4864 451216 4868
rect 451232 4924 451296 4928
rect 451232 4868 451236 4924
rect 451236 4868 451292 4924
rect 451292 4868 451296 4924
rect 451232 4864 451296 4868
rect 451312 4924 451376 4928
rect 451312 4868 451316 4924
rect 451316 4868 451372 4924
rect 451372 4868 451376 4924
rect 451312 4864 451376 4868
rect 486832 4924 486896 4928
rect 486832 4868 486836 4924
rect 486836 4868 486892 4924
rect 486892 4868 486896 4924
rect 486832 4864 486896 4868
rect 486912 4924 486976 4928
rect 486912 4868 486916 4924
rect 486916 4868 486972 4924
rect 486972 4868 486976 4924
rect 486912 4864 486976 4868
rect 486992 4924 487056 4928
rect 486992 4868 486996 4924
rect 486996 4868 487052 4924
rect 487052 4868 487056 4924
rect 486992 4864 487056 4868
rect 487072 4924 487136 4928
rect 487072 4868 487076 4924
rect 487076 4868 487132 4924
rect 487132 4868 487136 4924
rect 487072 4864 487136 4868
rect 487152 4924 487216 4928
rect 487152 4868 487156 4924
rect 487156 4868 487212 4924
rect 487212 4868 487216 4924
rect 487152 4864 487216 4868
rect 487232 4924 487296 4928
rect 487232 4868 487236 4924
rect 487236 4868 487292 4924
rect 487292 4868 487296 4924
rect 487232 4864 487296 4868
rect 487312 4924 487376 4928
rect 487312 4868 487316 4924
rect 487316 4868 487372 4924
rect 487372 4868 487376 4924
rect 487312 4864 487376 4868
rect 522832 4924 522896 4928
rect 522832 4868 522836 4924
rect 522836 4868 522892 4924
rect 522892 4868 522896 4924
rect 522832 4864 522896 4868
rect 522912 4924 522976 4928
rect 522912 4868 522916 4924
rect 522916 4868 522972 4924
rect 522972 4868 522976 4924
rect 522912 4864 522976 4868
rect 522992 4924 523056 4928
rect 522992 4868 522996 4924
rect 522996 4868 523052 4924
rect 523052 4868 523056 4924
rect 522992 4864 523056 4868
rect 523072 4924 523136 4928
rect 523072 4868 523076 4924
rect 523076 4868 523132 4924
rect 523132 4868 523136 4924
rect 523072 4864 523136 4868
rect 523152 4924 523216 4928
rect 523152 4868 523156 4924
rect 523156 4868 523212 4924
rect 523212 4868 523216 4924
rect 523152 4864 523216 4868
rect 523232 4924 523296 4928
rect 523232 4868 523236 4924
rect 523236 4868 523292 4924
rect 523292 4868 523296 4924
rect 523232 4864 523296 4868
rect 523312 4924 523376 4928
rect 523312 4868 523316 4924
rect 523316 4868 523372 4924
rect 523372 4868 523376 4924
rect 523312 4864 523376 4868
rect 558832 4924 558896 4928
rect 558832 4868 558836 4924
rect 558836 4868 558892 4924
rect 558892 4868 558896 4924
rect 558832 4864 558896 4868
rect 558912 4924 558976 4928
rect 558912 4868 558916 4924
rect 558916 4868 558972 4924
rect 558972 4868 558976 4924
rect 558912 4864 558976 4868
rect 558992 4924 559056 4928
rect 558992 4868 558996 4924
rect 558996 4868 559052 4924
rect 559052 4868 559056 4924
rect 558992 4864 559056 4868
rect 559072 4924 559136 4928
rect 559072 4868 559076 4924
rect 559076 4868 559132 4924
rect 559132 4868 559136 4924
rect 559072 4864 559136 4868
rect 559152 4924 559216 4928
rect 559152 4868 559156 4924
rect 559156 4868 559212 4924
rect 559212 4868 559216 4924
rect 559152 4864 559216 4868
rect 559232 4924 559296 4928
rect 559232 4868 559236 4924
rect 559236 4868 559292 4924
rect 559292 4868 559296 4924
rect 559232 4864 559296 4868
rect 559312 4924 559376 4928
rect 559312 4868 559316 4924
rect 559316 4868 559372 4924
rect 559372 4868 559376 4924
rect 559312 4864 559376 4868
rect 36832 4380 36896 4384
rect 36832 4324 36836 4380
rect 36836 4324 36892 4380
rect 36892 4324 36896 4380
rect 36832 4320 36896 4324
rect 36912 4380 36976 4384
rect 36912 4324 36916 4380
rect 36916 4324 36972 4380
rect 36972 4324 36976 4380
rect 36912 4320 36976 4324
rect 36992 4380 37056 4384
rect 36992 4324 36996 4380
rect 36996 4324 37052 4380
rect 37052 4324 37056 4380
rect 36992 4320 37056 4324
rect 37072 4380 37136 4384
rect 37072 4324 37076 4380
rect 37076 4324 37132 4380
rect 37132 4324 37136 4380
rect 37072 4320 37136 4324
rect 37152 4380 37216 4384
rect 37152 4324 37156 4380
rect 37156 4324 37212 4380
rect 37212 4324 37216 4380
rect 37152 4320 37216 4324
rect 37232 4380 37296 4384
rect 37232 4324 37236 4380
rect 37236 4324 37292 4380
rect 37292 4324 37296 4380
rect 37232 4320 37296 4324
rect 37312 4380 37376 4384
rect 37312 4324 37316 4380
rect 37316 4324 37372 4380
rect 37372 4324 37376 4380
rect 37312 4320 37376 4324
rect 72832 4380 72896 4384
rect 72832 4324 72836 4380
rect 72836 4324 72892 4380
rect 72892 4324 72896 4380
rect 72832 4320 72896 4324
rect 72912 4380 72976 4384
rect 72912 4324 72916 4380
rect 72916 4324 72972 4380
rect 72972 4324 72976 4380
rect 72912 4320 72976 4324
rect 72992 4380 73056 4384
rect 72992 4324 72996 4380
rect 72996 4324 73052 4380
rect 73052 4324 73056 4380
rect 72992 4320 73056 4324
rect 73072 4380 73136 4384
rect 73072 4324 73076 4380
rect 73076 4324 73132 4380
rect 73132 4324 73136 4380
rect 73072 4320 73136 4324
rect 73152 4380 73216 4384
rect 73152 4324 73156 4380
rect 73156 4324 73212 4380
rect 73212 4324 73216 4380
rect 73152 4320 73216 4324
rect 73232 4380 73296 4384
rect 73232 4324 73236 4380
rect 73236 4324 73292 4380
rect 73292 4324 73296 4380
rect 73232 4320 73296 4324
rect 73312 4380 73376 4384
rect 73312 4324 73316 4380
rect 73316 4324 73372 4380
rect 73372 4324 73376 4380
rect 73312 4320 73376 4324
rect 108832 4380 108896 4384
rect 108832 4324 108836 4380
rect 108836 4324 108892 4380
rect 108892 4324 108896 4380
rect 108832 4320 108896 4324
rect 108912 4380 108976 4384
rect 108912 4324 108916 4380
rect 108916 4324 108972 4380
rect 108972 4324 108976 4380
rect 108912 4320 108976 4324
rect 108992 4380 109056 4384
rect 108992 4324 108996 4380
rect 108996 4324 109052 4380
rect 109052 4324 109056 4380
rect 108992 4320 109056 4324
rect 109072 4380 109136 4384
rect 109072 4324 109076 4380
rect 109076 4324 109132 4380
rect 109132 4324 109136 4380
rect 109072 4320 109136 4324
rect 109152 4380 109216 4384
rect 109152 4324 109156 4380
rect 109156 4324 109212 4380
rect 109212 4324 109216 4380
rect 109152 4320 109216 4324
rect 109232 4380 109296 4384
rect 109232 4324 109236 4380
rect 109236 4324 109292 4380
rect 109292 4324 109296 4380
rect 109232 4320 109296 4324
rect 109312 4380 109376 4384
rect 109312 4324 109316 4380
rect 109316 4324 109372 4380
rect 109372 4324 109376 4380
rect 109312 4320 109376 4324
rect 144832 4380 144896 4384
rect 144832 4324 144836 4380
rect 144836 4324 144892 4380
rect 144892 4324 144896 4380
rect 144832 4320 144896 4324
rect 144912 4380 144976 4384
rect 144912 4324 144916 4380
rect 144916 4324 144972 4380
rect 144972 4324 144976 4380
rect 144912 4320 144976 4324
rect 144992 4380 145056 4384
rect 144992 4324 144996 4380
rect 144996 4324 145052 4380
rect 145052 4324 145056 4380
rect 144992 4320 145056 4324
rect 145072 4380 145136 4384
rect 145072 4324 145076 4380
rect 145076 4324 145132 4380
rect 145132 4324 145136 4380
rect 145072 4320 145136 4324
rect 145152 4380 145216 4384
rect 145152 4324 145156 4380
rect 145156 4324 145212 4380
rect 145212 4324 145216 4380
rect 145152 4320 145216 4324
rect 145232 4380 145296 4384
rect 145232 4324 145236 4380
rect 145236 4324 145292 4380
rect 145292 4324 145296 4380
rect 145232 4320 145296 4324
rect 145312 4380 145376 4384
rect 145312 4324 145316 4380
rect 145316 4324 145372 4380
rect 145372 4324 145376 4380
rect 145312 4320 145376 4324
rect 180832 4380 180896 4384
rect 180832 4324 180836 4380
rect 180836 4324 180892 4380
rect 180892 4324 180896 4380
rect 180832 4320 180896 4324
rect 180912 4380 180976 4384
rect 180912 4324 180916 4380
rect 180916 4324 180972 4380
rect 180972 4324 180976 4380
rect 180912 4320 180976 4324
rect 180992 4380 181056 4384
rect 180992 4324 180996 4380
rect 180996 4324 181052 4380
rect 181052 4324 181056 4380
rect 180992 4320 181056 4324
rect 181072 4380 181136 4384
rect 181072 4324 181076 4380
rect 181076 4324 181132 4380
rect 181132 4324 181136 4380
rect 181072 4320 181136 4324
rect 181152 4380 181216 4384
rect 181152 4324 181156 4380
rect 181156 4324 181212 4380
rect 181212 4324 181216 4380
rect 181152 4320 181216 4324
rect 181232 4380 181296 4384
rect 181232 4324 181236 4380
rect 181236 4324 181292 4380
rect 181292 4324 181296 4380
rect 181232 4320 181296 4324
rect 181312 4380 181376 4384
rect 181312 4324 181316 4380
rect 181316 4324 181372 4380
rect 181372 4324 181376 4380
rect 181312 4320 181376 4324
rect 216832 4380 216896 4384
rect 216832 4324 216836 4380
rect 216836 4324 216892 4380
rect 216892 4324 216896 4380
rect 216832 4320 216896 4324
rect 216912 4380 216976 4384
rect 216912 4324 216916 4380
rect 216916 4324 216972 4380
rect 216972 4324 216976 4380
rect 216912 4320 216976 4324
rect 216992 4380 217056 4384
rect 216992 4324 216996 4380
rect 216996 4324 217052 4380
rect 217052 4324 217056 4380
rect 216992 4320 217056 4324
rect 217072 4380 217136 4384
rect 217072 4324 217076 4380
rect 217076 4324 217132 4380
rect 217132 4324 217136 4380
rect 217072 4320 217136 4324
rect 217152 4380 217216 4384
rect 217152 4324 217156 4380
rect 217156 4324 217212 4380
rect 217212 4324 217216 4380
rect 217152 4320 217216 4324
rect 217232 4380 217296 4384
rect 217232 4324 217236 4380
rect 217236 4324 217292 4380
rect 217292 4324 217296 4380
rect 217232 4320 217296 4324
rect 217312 4380 217376 4384
rect 217312 4324 217316 4380
rect 217316 4324 217372 4380
rect 217372 4324 217376 4380
rect 217312 4320 217376 4324
rect 252832 4380 252896 4384
rect 252832 4324 252836 4380
rect 252836 4324 252892 4380
rect 252892 4324 252896 4380
rect 252832 4320 252896 4324
rect 252912 4380 252976 4384
rect 252912 4324 252916 4380
rect 252916 4324 252972 4380
rect 252972 4324 252976 4380
rect 252912 4320 252976 4324
rect 252992 4380 253056 4384
rect 252992 4324 252996 4380
rect 252996 4324 253052 4380
rect 253052 4324 253056 4380
rect 252992 4320 253056 4324
rect 253072 4380 253136 4384
rect 253072 4324 253076 4380
rect 253076 4324 253132 4380
rect 253132 4324 253136 4380
rect 253072 4320 253136 4324
rect 253152 4380 253216 4384
rect 253152 4324 253156 4380
rect 253156 4324 253212 4380
rect 253212 4324 253216 4380
rect 253152 4320 253216 4324
rect 253232 4380 253296 4384
rect 253232 4324 253236 4380
rect 253236 4324 253292 4380
rect 253292 4324 253296 4380
rect 253232 4320 253296 4324
rect 253312 4380 253376 4384
rect 253312 4324 253316 4380
rect 253316 4324 253372 4380
rect 253372 4324 253376 4380
rect 253312 4320 253376 4324
rect 288832 4380 288896 4384
rect 288832 4324 288836 4380
rect 288836 4324 288892 4380
rect 288892 4324 288896 4380
rect 288832 4320 288896 4324
rect 288912 4380 288976 4384
rect 288912 4324 288916 4380
rect 288916 4324 288972 4380
rect 288972 4324 288976 4380
rect 288912 4320 288976 4324
rect 288992 4380 289056 4384
rect 288992 4324 288996 4380
rect 288996 4324 289052 4380
rect 289052 4324 289056 4380
rect 288992 4320 289056 4324
rect 289072 4380 289136 4384
rect 289072 4324 289076 4380
rect 289076 4324 289132 4380
rect 289132 4324 289136 4380
rect 289072 4320 289136 4324
rect 289152 4380 289216 4384
rect 289152 4324 289156 4380
rect 289156 4324 289212 4380
rect 289212 4324 289216 4380
rect 289152 4320 289216 4324
rect 289232 4380 289296 4384
rect 289232 4324 289236 4380
rect 289236 4324 289292 4380
rect 289292 4324 289296 4380
rect 289232 4320 289296 4324
rect 289312 4380 289376 4384
rect 289312 4324 289316 4380
rect 289316 4324 289372 4380
rect 289372 4324 289376 4380
rect 289312 4320 289376 4324
rect 324832 4380 324896 4384
rect 324832 4324 324836 4380
rect 324836 4324 324892 4380
rect 324892 4324 324896 4380
rect 324832 4320 324896 4324
rect 324912 4380 324976 4384
rect 324912 4324 324916 4380
rect 324916 4324 324972 4380
rect 324972 4324 324976 4380
rect 324912 4320 324976 4324
rect 324992 4380 325056 4384
rect 324992 4324 324996 4380
rect 324996 4324 325052 4380
rect 325052 4324 325056 4380
rect 324992 4320 325056 4324
rect 325072 4380 325136 4384
rect 325072 4324 325076 4380
rect 325076 4324 325132 4380
rect 325132 4324 325136 4380
rect 325072 4320 325136 4324
rect 325152 4380 325216 4384
rect 325152 4324 325156 4380
rect 325156 4324 325212 4380
rect 325212 4324 325216 4380
rect 325152 4320 325216 4324
rect 325232 4380 325296 4384
rect 325232 4324 325236 4380
rect 325236 4324 325292 4380
rect 325292 4324 325296 4380
rect 325232 4320 325296 4324
rect 325312 4380 325376 4384
rect 325312 4324 325316 4380
rect 325316 4324 325372 4380
rect 325372 4324 325376 4380
rect 325312 4320 325376 4324
rect 360832 4380 360896 4384
rect 360832 4324 360836 4380
rect 360836 4324 360892 4380
rect 360892 4324 360896 4380
rect 360832 4320 360896 4324
rect 360912 4380 360976 4384
rect 360912 4324 360916 4380
rect 360916 4324 360972 4380
rect 360972 4324 360976 4380
rect 360912 4320 360976 4324
rect 360992 4380 361056 4384
rect 360992 4324 360996 4380
rect 360996 4324 361052 4380
rect 361052 4324 361056 4380
rect 360992 4320 361056 4324
rect 361072 4380 361136 4384
rect 361072 4324 361076 4380
rect 361076 4324 361132 4380
rect 361132 4324 361136 4380
rect 361072 4320 361136 4324
rect 361152 4380 361216 4384
rect 361152 4324 361156 4380
rect 361156 4324 361212 4380
rect 361212 4324 361216 4380
rect 361152 4320 361216 4324
rect 361232 4380 361296 4384
rect 361232 4324 361236 4380
rect 361236 4324 361292 4380
rect 361292 4324 361296 4380
rect 361232 4320 361296 4324
rect 361312 4380 361376 4384
rect 361312 4324 361316 4380
rect 361316 4324 361372 4380
rect 361372 4324 361376 4380
rect 361312 4320 361376 4324
rect 396832 4380 396896 4384
rect 396832 4324 396836 4380
rect 396836 4324 396892 4380
rect 396892 4324 396896 4380
rect 396832 4320 396896 4324
rect 396912 4380 396976 4384
rect 396912 4324 396916 4380
rect 396916 4324 396972 4380
rect 396972 4324 396976 4380
rect 396912 4320 396976 4324
rect 396992 4380 397056 4384
rect 396992 4324 396996 4380
rect 396996 4324 397052 4380
rect 397052 4324 397056 4380
rect 396992 4320 397056 4324
rect 397072 4380 397136 4384
rect 397072 4324 397076 4380
rect 397076 4324 397132 4380
rect 397132 4324 397136 4380
rect 397072 4320 397136 4324
rect 397152 4380 397216 4384
rect 397152 4324 397156 4380
rect 397156 4324 397212 4380
rect 397212 4324 397216 4380
rect 397152 4320 397216 4324
rect 397232 4380 397296 4384
rect 397232 4324 397236 4380
rect 397236 4324 397292 4380
rect 397292 4324 397296 4380
rect 397232 4320 397296 4324
rect 397312 4380 397376 4384
rect 397312 4324 397316 4380
rect 397316 4324 397372 4380
rect 397372 4324 397376 4380
rect 397312 4320 397376 4324
rect 432832 4380 432896 4384
rect 432832 4324 432836 4380
rect 432836 4324 432892 4380
rect 432892 4324 432896 4380
rect 432832 4320 432896 4324
rect 432912 4380 432976 4384
rect 432912 4324 432916 4380
rect 432916 4324 432972 4380
rect 432972 4324 432976 4380
rect 432912 4320 432976 4324
rect 432992 4380 433056 4384
rect 432992 4324 432996 4380
rect 432996 4324 433052 4380
rect 433052 4324 433056 4380
rect 432992 4320 433056 4324
rect 433072 4380 433136 4384
rect 433072 4324 433076 4380
rect 433076 4324 433132 4380
rect 433132 4324 433136 4380
rect 433072 4320 433136 4324
rect 433152 4380 433216 4384
rect 433152 4324 433156 4380
rect 433156 4324 433212 4380
rect 433212 4324 433216 4380
rect 433152 4320 433216 4324
rect 433232 4380 433296 4384
rect 433232 4324 433236 4380
rect 433236 4324 433292 4380
rect 433292 4324 433296 4380
rect 433232 4320 433296 4324
rect 433312 4380 433376 4384
rect 433312 4324 433316 4380
rect 433316 4324 433372 4380
rect 433372 4324 433376 4380
rect 433312 4320 433376 4324
rect 468832 4380 468896 4384
rect 468832 4324 468836 4380
rect 468836 4324 468892 4380
rect 468892 4324 468896 4380
rect 468832 4320 468896 4324
rect 468912 4380 468976 4384
rect 468912 4324 468916 4380
rect 468916 4324 468972 4380
rect 468972 4324 468976 4380
rect 468912 4320 468976 4324
rect 468992 4380 469056 4384
rect 468992 4324 468996 4380
rect 468996 4324 469052 4380
rect 469052 4324 469056 4380
rect 468992 4320 469056 4324
rect 469072 4380 469136 4384
rect 469072 4324 469076 4380
rect 469076 4324 469132 4380
rect 469132 4324 469136 4380
rect 469072 4320 469136 4324
rect 469152 4380 469216 4384
rect 469152 4324 469156 4380
rect 469156 4324 469212 4380
rect 469212 4324 469216 4380
rect 469152 4320 469216 4324
rect 469232 4380 469296 4384
rect 469232 4324 469236 4380
rect 469236 4324 469292 4380
rect 469292 4324 469296 4380
rect 469232 4320 469296 4324
rect 469312 4380 469376 4384
rect 469312 4324 469316 4380
rect 469316 4324 469372 4380
rect 469372 4324 469376 4380
rect 469312 4320 469376 4324
rect 504832 4380 504896 4384
rect 504832 4324 504836 4380
rect 504836 4324 504892 4380
rect 504892 4324 504896 4380
rect 504832 4320 504896 4324
rect 504912 4380 504976 4384
rect 504912 4324 504916 4380
rect 504916 4324 504972 4380
rect 504972 4324 504976 4380
rect 504912 4320 504976 4324
rect 504992 4380 505056 4384
rect 504992 4324 504996 4380
rect 504996 4324 505052 4380
rect 505052 4324 505056 4380
rect 504992 4320 505056 4324
rect 505072 4380 505136 4384
rect 505072 4324 505076 4380
rect 505076 4324 505132 4380
rect 505132 4324 505136 4380
rect 505072 4320 505136 4324
rect 505152 4380 505216 4384
rect 505152 4324 505156 4380
rect 505156 4324 505212 4380
rect 505212 4324 505216 4380
rect 505152 4320 505216 4324
rect 505232 4380 505296 4384
rect 505232 4324 505236 4380
rect 505236 4324 505292 4380
rect 505292 4324 505296 4380
rect 505232 4320 505296 4324
rect 505312 4380 505376 4384
rect 505312 4324 505316 4380
rect 505316 4324 505372 4380
rect 505372 4324 505376 4380
rect 505312 4320 505376 4324
rect 540832 4380 540896 4384
rect 540832 4324 540836 4380
rect 540836 4324 540892 4380
rect 540892 4324 540896 4380
rect 540832 4320 540896 4324
rect 540912 4380 540976 4384
rect 540912 4324 540916 4380
rect 540916 4324 540972 4380
rect 540972 4324 540976 4380
rect 540912 4320 540976 4324
rect 540992 4380 541056 4384
rect 540992 4324 540996 4380
rect 540996 4324 541052 4380
rect 541052 4324 541056 4380
rect 540992 4320 541056 4324
rect 541072 4380 541136 4384
rect 541072 4324 541076 4380
rect 541076 4324 541132 4380
rect 541132 4324 541136 4380
rect 541072 4320 541136 4324
rect 541152 4380 541216 4384
rect 541152 4324 541156 4380
rect 541156 4324 541212 4380
rect 541212 4324 541216 4380
rect 541152 4320 541216 4324
rect 541232 4380 541296 4384
rect 541232 4324 541236 4380
rect 541236 4324 541292 4380
rect 541292 4324 541296 4380
rect 541232 4320 541296 4324
rect 541312 4380 541376 4384
rect 541312 4324 541316 4380
rect 541316 4324 541372 4380
rect 541372 4324 541376 4380
rect 541312 4320 541376 4324
rect 576832 4380 576896 4384
rect 576832 4324 576836 4380
rect 576836 4324 576892 4380
rect 576892 4324 576896 4380
rect 576832 4320 576896 4324
rect 576912 4380 576976 4384
rect 576912 4324 576916 4380
rect 576916 4324 576972 4380
rect 576972 4324 576976 4380
rect 576912 4320 576976 4324
rect 576992 4380 577056 4384
rect 576992 4324 576996 4380
rect 576996 4324 577052 4380
rect 577052 4324 577056 4380
rect 576992 4320 577056 4324
rect 577072 4380 577136 4384
rect 577072 4324 577076 4380
rect 577076 4324 577132 4380
rect 577132 4324 577136 4380
rect 577072 4320 577136 4324
rect 577152 4380 577216 4384
rect 577152 4324 577156 4380
rect 577156 4324 577212 4380
rect 577212 4324 577216 4380
rect 577152 4320 577216 4324
rect 577232 4380 577296 4384
rect 577232 4324 577236 4380
rect 577236 4324 577292 4380
rect 577292 4324 577296 4380
rect 577232 4320 577296 4324
rect 577312 4380 577376 4384
rect 577312 4324 577316 4380
rect 577316 4324 577372 4380
rect 577372 4324 577376 4380
rect 577312 4320 577376 4324
rect 18832 3836 18896 3840
rect 18832 3780 18836 3836
rect 18836 3780 18892 3836
rect 18892 3780 18896 3836
rect 18832 3776 18896 3780
rect 18912 3836 18976 3840
rect 18912 3780 18916 3836
rect 18916 3780 18972 3836
rect 18972 3780 18976 3836
rect 18912 3776 18976 3780
rect 18992 3836 19056 3840
rect 18992 3780 18996 3836
rect 18996 3780 19052 3836
rect 19052 3780 19056 3836
rect 18992 3776 19056 3780
rect 19072 3836 19136 3840
rect 19072 3780 19076 3836
rect 19076 3780 19132 3836
rect 19132 3780 19136 3836
rect 19072 3776 19136 3780
rect 19152 3836 19216 3840
rect 19152 3780 19156 3836
rect 19156 3780 19212 3836
rect 19212 3780 19216 3836
rect 19152 3776 19216 3780
rect 19232 3836 19296 3840
rect 19232 3780 19236 3836
rect 19236 3780 19292 3836
rect 19292 3780 19296 3836
rect 19232 3776 19296 3780
rect 19312 3836 19376 3840
rect 19312 3780 19316 3836
rect 19316 3780 19372 3836
rect 19372 3780 19376 3836
rect 19312 3776 19376 3780
rect 54832 3836 54896 3840
rect 54832 3780 54836 3836
rect 54836 3780 54892 3836
rect 54892 3780 54896 3836
rect 54832 3776 54896 3780
rect 54912 3836 54976 3840
rect 54912 3780 54916 3836
rect 54916 3780 54972 3836
rect 54972 3780 54976 3836
rect 54912 3776 54976 3780
rect 54992 3836 55056 3840
rect 54992 3780 54996 3836
rect 54996 3780 55052 3836
rect 55052 3780 55056 3836
rect 54992 3776 55056 3780
rect 55072 3836 55136 3840
rect 55072 3780 55076 3836
rect 55076 3780 55132 3836
rect 55132 3780 55136 3836
rect 55072 3776 55136 3780
rect 55152 3836 55216 3840
rect 55152 3780 55156 3836
rect 55156 3780 55212 3836
rect 55212 3780 55216 3836
rect 55152 3776 55216 3780
rect 55232 3836 55296 3840
rect 55232 3780 55236 3836
rect 55236 3780 55292 3836
rect 55292 3780 55296 3836
rect 55232 3776 55296 3780
rect 55312 3836 55376 3840
rect 55312 3780 55316 3836
rect 55316 3780 55372 3836
rect 55372 3780 55376 3836
rect 55312 3776 55376 3780
rect 90832 3836 90896 3840
rect 90832 3780 90836 3836
rect 90836 3780 90892 3836
rect 90892 3780 90896 3836
rect 90832 3776 90896 3780
rect 90912 3836 90976 3840
rect 90912 3780 90916 3836
rect 90916 3780 90972 3836
rect 90972 3780 90976 3836
rect 90912 3776 90976 3780
rect 90992 3836 91056 3840
rect 90992 3780 90996 3836
rect 90996 3780 91052 3836
rect 91052 3780 91056 3836
rect 90992 3776 91056 3780
rect 91072 3836 91136 3840
rect 91072 3780 91076 3836
rect 91076 3780 91132 3836
rect 91132 3780 91136 3836
rect 91072 3776 91136 3780
rect 91152 3836 91216 3840
rect 91152 3780 91156 3836
rect 91156 3780 91212 3836
rect 91212 3780 91216 3836
rect 91152 3776 91216 3780
rect 91232 3836 91296 3840
rect 91232 3780 91236 3836
rect 91236 3780 91292 3836
rect 91292 3780 91296 3836
rect 91232 3776 91296 3780
rect 91312 3836 91376 3840
rect 91312 3780 91316 3836
rect 91316 3780 91372 3836
rect 91372 3780 91376 3836
rect 91312 3776 91376 3780
rect 126832 3836 126896 3840
rect 126832 3780 126836 3836
rect 126836 3780 126892 3836
rect 126892 3780 126896 3836
rect 126832 3776 126896 3780
rect 126912 3836 126976 3840
rect 126912 3780 126916 3836
rect 126916 3780 126972 3836
rect 126972 3780 126976 3836
rect 126912 3776 126976 3780
rect 126992 3836 127056 3840
rect 126992 3780 126996 3836
rect 126996 3780 127052 3836
rect 127052 3780 127056 3836
rect 126992 3776 127056 3780
rect 127072 3836 127136 3840
rect 127072 3780 127076 3836
rect 127076 3780 127132 3836
rect 127132 3780 127136 3836
rect 127072 3776 127136 3780
rect 127152 3836 127216 3840
rect 127152 3780 127156 3836
rect 127156 3780 127212 3836
rect 127212 3780 127216 3836
rect 127152 3776 127216 3780
rect 127232 3836 127296 3840
rect 127232 3780 127236 3836
rect 127236 3780 127292 3836
rect 127292 3780 127296 3836
rect 127232 3776 127296 3780
rect 127312 3836 127376 3840
rect 127312 3780 127316 3836
rect 127316 3780 127372 3836
rect 127372 3780 127376 3836
rect 127312 3776 127376 3780
rect 162832 3836 162896 3840
rect 162832 3780 162836 3836
rect 162836 3780 162892 3836
rect 162892 3780 162896 3836
rect 162832 3776 162896 3780
rect 162912 3836 162976 3840
rect 162912 3780 162916 3836
rect 162916 3780 162972 3836
rect 162972 3780 162976 3836
rect 162912 3776 162976 3780
rect 162992 3836 163056 3840
rect 162992 3780 162996 3836
rect 162996 3780 163052 3836
rect 163052 3780 163056 3836
rect 162992 3776 163056 3780
rect 163072 3836 163136 3840
rect 163072 3780 163076 3836
rect 163076 3780 163132 3836
rect 163132 3780 163136 3836
rect 163072 3776 163136 3780
rect 163152 3836 163216 3840
rect 163152 3780 163156 3836
rect 163156 3780 163212 3836
rect 163212 3780 163216 3836
rect 163152 3776 163216 3780
rect 163232 3836 163296 3840
rect 163232 3780 163236 3836
rect 163236 3780 163292 3836
rect 163292 3780 163296 3836
rect 163232 3776 163296 3780
rect 163312 3836 163376 3840
rect 163312 3780 163316 3836
rect 163316 3780 163372 3836
rect 163372 3780 163376 3836
rect 163312 3776 163376 3780
rect 198832 3836 198896 3840
rect 198832 3780 198836 3836
rect 198836 3780 198892 3836
rect 198892 3780 198896 3836
rect 198832 3776 198896 3780
rect 198912 3836 198976 3840
rect 198912 3780 198916 3836
rect 198916 3780 198972 3836
rect 198972 3780 198976 3836
rect 198912 3776 198976 3780
rect 198992 3836 199056 3840
rect 198992 3780 198996 3836
rect 198996 3780 199052 3836
rect 199052 3780 199056 3836
rect 198992 3776 199056 3780
rect 199072 3836 199136 3840
rect 199072 3780 199076 3836
rect 199076 3780 199132 3836
rect 199132 3780 199136 3836
rect 199072 3776 199136 3780
rect 199152 3836 199216 3840
rect 199152 3780 199156 3836
rect 199156 3780 199212 3836
rect 199212 3780 199216 3836
rect 199152 3776 199216 3780
rect 199232 3836 199296 3840
rect 199232 3780 199236 3836
rect 199236 3780 199292 3836
rect 199292 3780 199296 3836
rect 199232 3776 199296 3780
rect 199312 3836 199376 3840
rect 199312 3780 199316 3836
rect 199316 3780 199372 3836
rect 199372 3780 199376 3836
rect 199312 3776 199376 3780
rect 234832 3836 234896 3840
rect 234832 3780 234836 3836
rect 234836 3780 234892 3836
rect 234892 3780 234896 3836
rect 234832 3776 234896 3780
rect 234912 3836 234976 3840
rect 234912 3780 234916 3836
rect 234916 3780 234972 3836
rect 234972 3780 234976 3836
rect 234912 3776 234976 3780
rect 234992 3836 235056 3840
rect 234992 3780 234996 3836
rect 234996 3780 235052 3836
rect 235052 3780 235056 3836
rect 234992 3776 235056 3780
rect 235072 3836 235136 3840
rect 235072 3780 235076 3836
rect 235076 3780 235132 3836
rect 235132 3780 235136 3836
rect 235072 3776 235136 3780
rect 235152 3836 235216 3840
rect 235152 3780 235156 3836
rect 235156 3780 235212 3836
rect 235212 3780 235216 3836
rect 235152 3776 235216 3780
rect 235232 3836 235296 3840
rect 235232 3780 235236 3836
rect 235236 3780 235292 3836
rect 235292 3780 235296 3836
rect 235232 3776 235296 3780
rect 235312 3836 235376 3840
rect 235312 3780 235316 3836
rect 235316 3780 235372 3836
rect 235372 3780 235376 3836
rect 235312 3776 235376 3780
rect 270832 3836 270896 3840
rect 270832 3780 270836 3836
rect 270836 3780 270892 3836
rect 270892 3780 270896 3836
rect 270832 3776 270896 3780
rect 270912 3836 270976 3840
rect 270912 3780 270916 3836
rect 270916 3780 270972 3836
rect 270972 3780 270976 3836
rect 270912 3776 270976 3780
rect 270992 3836 271056 3840
rect 270992 3780 270996 3836
rect 270996 3780 271052 3836
rect 271052 3780 271056 3836
rect 270992 3776 271056 3780
rect 271072 3836 271136 3840
rect 271072 3780 271076 3836
rect 271076 3780 271132 3836
rect 271132 3780 271136 3836
rect 271072 3776 271136 3780
rect 271152 3836 271216 3840
rect 271152 3780 271156 3836
rect 271156 3780 271212 3836
rect 271212 3780 271216 3836
rect 271152 3776 271216 3780
rect 271232 3836 271296 3840
rect 271232 3780 271236 3836
rect 271236 3780 271292 3836
rect 271292 3780 271296 3836
rect 271232 3776 271296 3780
rect 271312 3836 271376 3840
rect 271312 3780 271316 3836
rect 271316 3780 271372 3836
rect 271372 3780 271376 3836
rect 271312 3776 271376 3780
rect 306832 3836 306896 3840
rect 306832 3780 306836 3836
rect 306836 3780 306892 3836
rect 306892 3780 306896 3836
rect 306832 3776 306896 3780
rect 306912 3836 306976 3840
rect 306912 3780 306916 3836
rect 306916 3780 306972 3836
rect 306972 3780 306976 3836
rect 306912 3776 306976 3780
rect 306992 3836 307056 3840
rect 306992 3780 306996 3836
rect 306996 3780 307052 3836
rect 307052 3780 307056 3836
rect 306992 3776 307056 3780
rect 307072 3836 307136 3840
rect 307072 3780 307076 3836
rect 307076 3780 307132 3836
rect 307132 3780 307136 3836
rect 307072 3776 307136 3780
rect 307152 3836 307216 3840
rect 307152 3780 307156 3836
rect 307156 3780 307212 3836
rect 307212 3780 307216 3836
rect 307152 3776 307216 3780
rect 307232 3836 307296 3840
rect 307232 3780 307236 3836
rect 307236 3780 307292 3836
rect 307292 3780 307296 3836
rect 307232 3776 307296 3780
rect 307312 3836 307376 3840
rect 307312 3780 307316 3836
rect 307316 3780 307372 3836
rect 307372 3780 307376 3836
rect 307312 3776 307376 3780
rect 342832 3836 342896 3840
rect 342832 3780 342836 3836
rect 342836 3780 342892 3836
rect 342892 3780 342896 3836
rect 342832 3776 342896 3780
rect 342912 3836 342976 3840
rect 342912 3780 342916 3836
rect 342916 3780 342972 3836
rect 342972 3780 342976 3836
rect 342912 3776 342976 3780
rect 342992 3836 343056 3840
rect 342992 3780 342996 3836
rect 342996 3780 343052 3836
rect 343052 3780 343056 3836
rect 342992 3776 343056 3780
rect 343072 3836 343136 3840
rect 343072 3780 343076 3836
rect 343076 3780 343132 3836
rect 343132 3780 343136 3836
rect 343072 3776 343136 3780
rect 343152 3836 343216 3840
rect 343152 3780 343156 3836
rect 343156 3780 343212 3836
rect 343212 3780 343216 3836
rect 343152 3776 343216 3780
rect 343232 3836 343296 3840
rect 343232 3780 343236 3836
rect 343236 3780 343292 3836
rect 343292 3780 343296 3836
rect 343232 3776 343296 3780
rect 343312 3836 343376 3840
rect 343312 3780 343316 3836
rect 343316 3780 343372 3836
rect 343372 3780 343376 3836
rect 343312 3776 343376 3780
rect 378832 3836 378896 3840
rect 378832 3780 378836 3836
rect 378836 3780 378892 3836
rect 378892 3780 378896 3836
rect 378832 3776 378896 3780
rect 378912 3836 378976 3840
rect 378912 3780 378916 3836
rect 378916 3780 378972 3836
rect 378972 3780 378976 3836
rect 378912 3776 378976 3780
rect 378992 3836 379056 3840
rect 378992 3780 378996 3836
rect 378996 3780 379052 3836
rect 379052 3780 379056 3836
rect 378992 3776 379056 3780
rect 379072 3836 379136 3840
rect 379072 3780 379076 3836
rect 379076 3780 379132 3836
rect 379132 3780 379136 3836
rect 379072 3776 379136 3780
rect 379152 3836 379216 3840
rect 379152 3780 379156 3836
rect 379156 3780 379212 3836
rect 379212 3780 379216 3836
rect 379152 3776 379216 3780
rect 379232 3836 379296 3840
rect 379232 3780 379236 3836
rect 379236 3780 379292 3836
rect 379292 3780 379296 3836
rect 379232 3776 379296 3780
rect 379312 3836 379376 3840
rect 379312 3780 379316 3836
rect 379316 3780 379372 3836
rect 379372 3780 379376 3836
rect 379312 3776 379376 3780
rect 414832 3836 414896 3840
rect 414832 3780 414836 3836
rect 414836 3780 414892 3836
rect 414892 3780 414896 3836
rect 414832 3776 414896 3780
rect 414912 3836 414976 3840
rect 414912 3780 414916 3836
rect 414916 3780 414972 3836
rect 414972 3780 414976 3836
rect 414912 3776 414976 3780
rect 414992 3836 415056 3840
rect 414992 3780 414996 3836
rect 414996 3780 415052 3836
rect 415052 3780 415056 3836
rect 414992 3776 415056 3780
rect 415072 3836 415136 3840
rect 415072 3780 415076 3836
rect 415076 3780 415132 3836
rect 415132 3780 415136 3836
rect 415072 3776 415136 3780
rect 415152 3836 415216 3840
rect 415152 3780 415156 3836
rect 415156 3780 415212 3836
rect 415212 3780 415216 3836
rect 415152 3776 415216 3780
rect 415232 3836 415296 3840
rect 415232 3780 415236 3836
rect 415236 3780 415292 3836
rect 415292 3780 415296 3836
rect 415232 3776 415296 3780
rect 415312 3836 415376 3840
rect 415312 3780 415316 3836
rect 415316 3780 415372 3836
rect 415372 3780 415376 3836
rect 415312 3776 415376 3780
rect 450832 3836 450896 3840
rect 450832 3780 450836 3836
rect 450836 3780 450892 3836
rect 450892 3780 450896 3836
rect 450832 3776 450896 3780
rect 450912 3836 450976 3840
rect 450912 3780 450916 3836
rect 450916 3780 450972 3836
rect 450972 3780 450976 3836
rect 450912 3776 450976 3780
rect 450992 3836 451056 3840
rect 450992 3780 450996 3836
rect 450996 3780 451052 3836
rect 451052 3780 451056 3836
rect 450992 3776 451056 3780
rect 451072 3836 451136 3840
rect 451072 3780 451076 3836
rect 451076 3780 451132 3836
rect 451132 3780 451136 3836
rect 451072 3776 451136 3780
rect 451152 3836 451216 3840
rect 451152 3780 451156 3836
rect 451156 3780 451212 3836
rect 451212 3780 451216 3836
rect 451152 3776 451216 3780
rect 451232 3836 451296 3840
rect 451232 3780 451236 3836
rect 451236 3780 451292 3836
rect 451292 3780 451296 3836
rect 451232 3776 451296 3780
rect 451312 3836 451376 3840
rect 451312 3780 451316 3836
rect 451316 3780 451372 3836
rect 451372 3780 451376 3836
rect 451312 3776 451376 3780
rect 486832 3836 486896 3840
rect 486832 3780 486836 3836
rect 486836 3780 486892 3836
rect 486892 3780 486896 3836
rect 486832 3776 486896 3780
rect 486912 3836 486976 3840
rect 486912 3780 486916 3836
rect 486916 3780 486972 3836
rect 486972 3780 486976 3836
rect 486912 3776 486976 3780
rect 486992 3836 487056 3840
rect 486992 3780 486996 3836
rect 486996 3780 487052 3836
rect 487052 3780 487056 3836
rect 486992 3776 487056 3780
rect 487072 3836 487136 3840
rect 487072 3780 487076 3836
rect 487076 3780 487132 3836
rect 487132 3780 487136 3836
rect 487072 3776 487136 3780
rect 487152 3836 487216 3840
rect 487152 3780 487156 3836
rect 487156 3780 487212 3836
rect 487212 3780 487216 3836
rect 487152 3776 487216 3780
rect 487232 3836 487296 3840
rect 487232 3780 487236 3836
rect 487236 3780 487292 3836
rect 487292 3780 487296 3836
rect 487232 3776 487296 3780
rect 487312 3836 487376 3840
rect 487312 3780 487316 3836
rect 487316 3780 487372 3836
rect 487372 3780 487376 3836
rect 487312 3776 487376 3780
rect 522832 3836 522896 3840
rect 522832 3780 522836 3836
rect 522836 3780 522892 3836
rect 522892 3780 522896 3836
rect 522832 3776 522896 3780
rect 522912 3836 522976 3840
rect 522912 3780 522916 3836
rect 522916 3780 522972 3836
rect 522972 3780 522976 3836
rect 522912 3776 522976 3780
rect 522992 3836 523056 3840
rect 522992 3780 522996 3836
rect 522996 3780 523052 3836
rect 523052 3780 523056 3836
rect 522992 3776 523056 3780
rect 523072 3836 523136 3840
rect 523072 3780 523076 3836
rect 523076 3780 523132 3836
rect 523132 3780 523136 3836
rect 523072 3776 523136 3780
rect 523152 3836 523216 3840
rect 523152 3780 523156 3836
rect 523156 3780 523212 3836
rect 523212 3780 523216 3836
rect 523152 3776 523216 3780
rect 523232 3836 523296 3840
rect 523232 3780 523236 3836
rect 523236 3780 523292 3836
rect 523292 3780 523296 3836
rect 523232 3776 523296 3780
rect 523312 3836 523376 3840
rect 523312 3780 523316 3836
rect 523316 3780 523372 3836
rect 523372 3780 523376 3836
rect 523312 3776 523376 3780
rect 558832 3836 558896 3840
rect 558832 3780 558836 3836
rect 558836 3780 558892 3836
rect 558892 3780 558896 3836
rect 558832 3776 558896 3780
rect 558912 3836 558976 3840
rect 558912 3780 558916 3836
rect 558916 3780 558972 3836
rect 558972 3780 558976 3836
rect 558912 3776 558976 3780
rect 558992 3836 559056 3840
rect 558992 3780 558996 3836
rect 558996 3780 559052 3836
rect 559052 3780 559056 3836
rect 558992 3776 559056 3780
rect 559072 3836 559136 3840
rect 559072 3780 559076 3836
rect 559076 3780 559132 3836
rect 559132 3780 559136 3836
rect 559072 3776 559136 3780
rect 559152 3836 559216 3840
rect 559152 3780 559156 3836
rect 559156 3780 559212 3836
rect 559212 3780 559216 3836
rect 559152 3776 559216 3780
rect 559232 3836 559296 3840
rect 559232 3780 559236 3836
rect 559236 3780 559292 3836
rect 559292 3780 559296 3836
rect 559232 3776 559296 3780
rect 559312 3836 559376 3840
rect 559312 3780 559316 3836
rect 559316 3780 559372 3836
rect 559372 3780 559376 3836
rect 559312 3776 559376 3780
rect 36832 3292 36896 3296
rect 36832 3236 36836 3292
rect 36836 3236 36892 3292
rect 36892 3236 36896 3292
rect 36832 3232 36896 3236
rect 36912 3292 36976 3296
rect 36912 3236 36916 3292
rect 36916 3236 36972 3292
rect 36972 3236 36976 3292
rect 36912 3232 36976 3236
rect 36992 3292 37056 3296
rect 36992 3236 36996 3292
rect 36996 3236 37052 3292
rect 37052 3236 37056 3292
rect 36992 3232 37056 3236
rect 37072 3292 37136 3296
rect 37072 3236 37076 3292
rect 37076 3236 37132 3292
rect 37132 3236 37136 3292
rect 37072 3232 37136 3236
rect 37152 3292 37216 3296
rect 37152 3236 37156 3292
rect 37156 3236 37212 3292
rect 37212 3236 37216 3292
rect 37152 3232 37216 3236
rect 37232 3292 37296 3296
rect 37232 3236 37236 3292
rect 37236 3236 37292 3292
rect 37292 3236 37296 3292
rect 37232 3232 37296 3236
rect 37312 3292 37376 3296
rect 37312 3236 37316 3292
rect 37316 3236 37372 3292
rect 37372 3236 37376 3292
rect 37312 3232 37376 3236
rect 72832 3292 72896 3296
rect 72832 3236 72836 3292
rect 72836 3236 72892 3292
rect 72892 3236 72896 3292
rect 72832 3232 72896 3236
rect 72912 3292 72976 3296
rect 72912 3236 72916 3292
rect 72916 3236 72972 3292
rect 72972 3236 72976 3292
rect 72912 3232 72976 3236
rect 72992 3292 73056 3296
rect 72992 3236 72996 3292
rect 72996 3236 73052 3292
rect 73052 3236 73056 3292
rect 72992 3232 73056 3236
rect 73072 3292 73136 3296
rect 73072 3236 73076 3292
rect 73076 3236 73132 3292
rect 73132 3236 73136 3292
rect 73072 3232 73136 3236
rect 73152 3292 73216 3296
rect 73152 3236 73156 3292
rect 73156 3236 73212 3292
rect 73212 3236 73216 3292
rect 73152 3232 73216 3236
rect 73232 3292 73296 3296
rect 73232 3236 73236 3292
rect 73236 3236 73292 3292
rect 73292 3236 73296 3292
rect 73232 3232 73296 3236
rect 73312 3292 73376 3296
rect 73312 3236 73316 3292
rect 73316 3236 73372 3292
rect 73372 3236 73376 3292
rect 73312 3232 73376 3236
rect 108832 3292 108896 3296
rect 108832 3236 108836 3292
rect 108836 3236 108892 3292
rect 108892 3236 108896 3292
rect 108832 3232 108896 3236
rect 108912 3292 108976 3296
rect 108912 3236 108916 3292
rect 108916 3236 108972 3292
rect 108972 3236 108976 3292
rect 108912 3232 108976 3236
rect 108992 3292 109056 3296
rect 108992 3236 108996 3292
rect 108996 3236 109052 3292
rect 109052 3236 109056 3292
rect 108992 3232 109056 3236
rect 109072 3292 109136 3296
rect 109072 3236 109076 3292
rect 109076 3236 109132 3292
rect 109132 3236 109136 3292
rect 109072 3232 109136 3236
rect 109152 3292 109216 3296
rect 109152 3236 109156 3292
rect 109156 3236 109212 3292
rect 109212 3236 109216 3292
rect 109152 3232 109216 3236
rect 109232 3292 109296 3296
rect 109232 3236 109236 3292
rect 109236 3236 109292 3292
rect 109292 3236 109296 3292
rect 109232 3232 109296 3236
rect 109312 3292 109376 3296
rect 109312 3236 109316 3292
rect 109316 3236 109372 3292
rect 109372 3236 109376 3292
rect 109312 3232 109376 3236
rect 144832 3292 144896 3296
rect 144832 3236 144836 3292
rect 144836 3236 144892 3292
rect 144892 3236 144896 3292
rect 144832 3232 144896 3236
rect 144912 3292 144976 3296
rect 144912 3236 144916 3292
rect 144916 3236 144972 3292
rect 144972 3236 144976 3292
rect 144912 3232 144976 3236
rect 144992 3292 145056 3296
rect 144992 3236 144996 3292
rect 144996 3236 145052 3292
rect 145052 3236 145056 3292
rect 144992 3232 145056 3236
rect 145072 3292 145136 3296
rect 145072 3236 145076 3292
rect 145076 3236 145132 3292
rect 145132 3236 145136 3292
rect 145072 3232 145136 3236
rect 145152 3292 145216 3296
rect 145152 3236 145156 3292
rect 145156 3236 145212 3292
rect 145212 3236 145216 3292
rect 145152 3232 145216 3236
rect 145232 3292 145296 3296
rect 145232 3236 145236 3292
rect 145236 3236 145292 3292
rect 145292 3236 145296 3292
rect 145232 3232 145296 3236
rect 145312 3292 145376 3296
rect 145312 3236 145316 3292
rect 145316 3236 145372 3292
rect 145372 3236 145376 3292
rect 145312 3232 145376 3236
rect 180832 3292 180896 3296
rect 180832 3236 180836 3292
rect 180836 3236 180892 3292
rect 180892 3236 180896 3292
rect 180832 3232 180896 3236
rect 180912 3292 180976 3296
rect 180912 3236 180916 3292
rect 180916 3236 180972 3292
rect 180972 3236 180976 3292
rect 180912 3232 180976 3236
rect 180992 3292 181056 3296
rect 180992 3236 180996 3292
rect 180996 3236 181052 3292
rect 181052 3236 181056 3292
rect 180992 3232 181056 3236
rect 181072 3292 181136 3296
rect 181072 3236 181076 3292
rect 181076 3236 181132 3292
rect 181132 3236 181136 3292
rect 181072 3232 181136 3236
rect 181152 3292 181216 3296
rect 181152 3236 181156 3292
rect 181156 3236 181212 3292
rect 181212 3236 181216 3292
rect 181152 3232 181216 3236
rect 181232 3292 181296 3296
rect 181232 3236 181236 3292
rect 181236 3236 181292 3292
rect 181292 3236 181296 3292
rect 181232 3232 181296 3236
rect 181312 3292 181376 3296
rect 181312 3236 181316 3292
rect 181316 3236 181372 3292
rect 181372 3236 181376 3292
rect 181312 3232 181376 3236
rect 216832 3292 216896 3296
rect 216832 3236 216836 3292
rect 216836 3236 216892 3292
rect 216892 3236 216896 3292
rect 216832 3232 216896 3236
rect 216912 3292 216976 3296
rect 216912 3236 216916 3292
rect 216916 3236 216972 3292
rect 216972 3236 216976 3292
rect 216912 3232 216976 3236
rect 216992 3292 217056 3296
rect 216992 3236 216996 3292
rect 216996 3236 217052 3292
rect 217052 3236 217056 3292
rect 216992 3232 217056 3236
rect 217072 3292 217136 3296
rect 217072 3236 217076 3292
rect 217076 3236 217132 3292
rect 217132 3236 217136 3292
rect 217072 3232 217136 3236
rect 217152 3292 217216 3296
rect 217152 3236 217156 3292
rect 217156 3236 217212 3292
rect 217212 3236 217216 3292
rect 217152 3232 217216 3236
rect 217232 3292 217296 3296
rect 217232 3236 217236 3292
rect 217236 3236 217292 3292
rect 217292 3236 217296 3292
rect 217232 3232 217296 3236
rect 217312 3292 217376 3296
rect 217312 3236 217316 3292
rect 217316 3236 217372 3292
rect 217372 3236 217376 3292
rect 217312 3232 217376 3236
rect 252832 3292 252896 3296
rect 252832 3236 252836 3292
rect 252836 3236 252892 3292
rect 252892 3236 252896 3292
rect 252832 3232 252896 3236
rect 252912 3292 252976 3296
rect 252912 3236 252916 3292
rect 252916 3236 252972 3292
rect 252972 3236 252976 3292
rect 252912 3232 252976 3236
rect 252992 3292 253056 3296
rect 252992 3236 252996 3292
rect 252996 3236 253052 3292
rect 253052 3236 253056 3292
rect 252992 3232 253056 3236
rect 253072 3292 253136 3296
rect 253072 3236 253076 3292
rect 253076 3236 253132 3292
rect 253132 3236 253136 3292
rect 253072 3232 253136 3236
rect 253152 3292 253216 3296
rect 253152 3236 253156 3292
rect 253156 3236 253212 3292
rect 253212 3236 253216 3292
rect 253152 3232 253216 3236
rect 253232 3292 253296 3296
rect 253232 3236 253236 3292
rect 253236 3236 253292 3292
rect 253292 3236 253296 3292
rect 253232 3232 253296 3236
rect 253312 3292 253376 3296
rect 253312 3236 253316 3292
rect 253316 3236 253372 3292
rect 253372 3236 253376 3292
rect 253312 3232 253376 3236
rect 288832 3292 288896 3296
rect 288832 3236 288836 3292
rect 288836 3236 288892 3292
rect 288892 3236 288896 3292
rect 288832 3232 288896 3236
rect 288912 3292 288976 3296
rect 288912 3236 288916 3292
rect 288916 3236 288972 3292
rect 288972 3236 288976 3292
rect 288912 3232 288976 3236
rect 288992 3292 289056 3296
rect 288992 3236 288996 3292
rect 288996 3236 289052 3292
rect 289052 3236 289056 3292
rect 288992 3232 289056 3236
rect 289072 3292 289136 3296
rect 289072 3236 289076 3292
rect 289076 3236 289132 3292
rect 289132 3236 289136 3292
rect 289072 3232 289136 3236
rect 289152 3292 289216 3296
rect 289152 3236 289156 3292
rect 289156 3236 289212 3292
rect 289212 3236 289216 3292
rect 289152 3232 289216 3236
rect 289232 3292 289296 3296
rect 289232 3236 289236 3292
rect 289236 3236 289292 3292
rect 289292 3236 289296 3292
rect 289232 3232 289296 3236
rect 289312 3292 289376 3296
rect 289312 3236 289316 3292
rect 289316 3236 289372 3292
rect 289372 3236 289376 3292
rect 289312 3232 289376 3236
rect 324832 3292 324896 3296
rect 324832 3236 324836 3292
rect 324836 3236 324892 3292
rect 324892 3236 324896 3292
rect 324832 3232 324896 3236
rect 324912 3292 324976 3296
rect 324912 3236 324916 3292
rect 324916 3236 324972 3292
rect 324972 3236 324976 3292
rect 324912 3232 324976 3236
rect 324992 3292 325056 3296
rect 324992 3236 324996 3292
rect 324996 3236 325052 3292
rect 325052 3236 325056 3292
rect 324992 3232 325056 3236
rect 325072 3292 325136 3296
rect 325072 3236 325076 3292
rect 325076 3236 325132 3292
rect 325132 3236 325136 3292
rect 325072 3232 325136 3236
rect 325152 3292 325216 3296
rect 325152 3236 325156 3292
rect 325156 3236 325212 3292
rect 325212 3236 325216 3292
rect 325152 3232 325216 3236
rect 325232 3292 325296 3296
rect 325232 3236 325236 3292
rect 325236 3236 325292 3292
rect 325292 3236 325296 3292
rect 325232 3232 325296 3236
rect 325312 3292 325376 3296
rect 325312 3236 325316 3292
rect 325316 3236 325372 3292
rect 325372 3236 325376 3292
rect 325312 3232 325376 3236
rect 360832 3292 360896 3296
rect 360832 3236 360836 3292
rect 360836 3236 360892 3292
rect 360892 3236 360896 3292
rect 360832 3232 360896 3236
rect 360912 3292 360976 3296
rect 360912 3236 360916 3292
rect 360916 3236 360972 3292
rect 360972 3236 360976 3292
rect 360912 3232 360976 3236
rect 360992 3292 361056 3296
rect 360992 3236 360996 3292
rect 360996 3236 361052 3292
rect 361052 3236 361056 3292
rect 360992 3232 361056 3236
rect 361072 3292 361136 3296
rect 361072 3236 361076 3292
rect 361076 3236 361132 3292
rect 361132 3236 361136 3292
rect 361072 3232 361136 3236
rect 361152 3292 361216 3296
rect 361152 3236 361156 3292
rect 361156 3236 361212 3292
rect 361212 3236 361216 3292
rect 361152 3232 361216 3236
rect 361232 3292 361296 3296
rect 361232 3236 361236 3292
rect 361236 3236 361292 3292
rect 361292 3236 361296 3292
rect 361232 3232 361296 3236
rect 361312 3292 361376 3296
rect 361312 3236 361316 3292
rect 361316 3236 361372 3292
rect 361372 3236 361376 3292
rect 361312 3232 361376 3236
rect 396832 3292 396896 3296
rect 396832 3236 396836 3292
rect 396836 3236 396892 3292
rect 396892 3236 396896 3292
rect 396832 3232 396896 3236
rect 396912 3292 396976 3296
rect 396912 3236 396916 3292
rect 396916 3236 396972 3292
rect 396972 3236 396976 3292
rect 396912 3232 396976 3236
rect 396992 3292 397056 3296
rect 396992 3236 396996 3292
rect 396996 3236 397052 3292
rect 397052 3236 397056 3292
rect 396992 3232 397056 3236
rect 397072 3292 397136 3296
rect 397072 3236 397076 3292
rect 397076 3236 397132 3292
rect 397132 3236 397136 3292
rect 397072 3232 397136 3236
rect 397152 3292 397216 3296
rect 397152 3236 397156 3292
rect 397156 3236 397212 3292
rect 397212 3236 397216 3292
rect 397152 3232 397216 3236
rect 397232 3292 397296 3296
rect 397232 3236 397236 3292
rect 397236 3236 397292 3292
rect 397292 3236 397296 3292
rect 397232 3232 397296 3236
rect 397312 3292 397376 3296
rect 397312 3236 397316 3292
rect 397316 3236 397372 3292
rect 397372 3236 397376 3292
rect 397312 3232 397376 3236
rect 432832 3292 432896 3296
rect 432832 3236 432836 3292
rect 432836 3236 432892 3292
rect 432892 3236 432896 3292
rect 432832 3232 432896 3236
rect 432912 3292 432976 3296
rect 432912 3236 432916 3292
rect 432916 3236 432972 3292
rect 432972 3236 432976 3292
rect 432912 3232 432976 3236
rect 432992 3292 433056 3296
rect 432992 3236 432996 3292
rect 432996 3236 433052 3292
rect 433052 3236 433056 3292
rect 432992 3232 433056 3236
rect 433072 3292 433136 3296
rect 433072 3236 433076 3292
rect 433076 3236 433132 3292
rect 433132 3236 433136 3292
rect 433072 3232 433136 3236
rect 433152 3292 433216 3296
rect 433152 3236 433156 3292
rect 433156 3236 433212 3292
rect 433212 3236 433216 3292
rect 433152 3232 433216 3236
rect 433232 3292 433296 3296
rect 433232 3236 433236 3292
rect 433236 3236 433292 3292
rect 433292 3236 433296 3292
rect 433232 3232 433296 3236
rect 433312 3292 433376 3296
rect 433312 3236 433316 3292
rect 433316 3236 433372 3292
rect 433372 3236 433376 3292
rect 433312 3232 433376 3236
rect 468832 3292 468896 3296
rect 468832 3236 468836 3292
rect 468836 3236 468892 3292
rect 468892 3236 468896 3292
rect 468832 3232 468896 3236
rect 468912 3292 468976 3296
rect 468912 3236 468916 3292
rect 468916 3236 468972 3292
rect 468972 3236 468976 3292
rect 468912 3232 468976 3236
rect 468992 3292 469056 3296
rect 468992 3236 468996 3292
rect 468996 3236 469052 3292
rect 469052 3236 469056 3292
rect 468992 3232 469056 3236
rect 469072 3292 469136 3296
rect 469072 3236 469076 3292
rect 469076 3236 469132 3292
rect 469132 3236 469136 3292
rect 469072 3232 469136 3236
rect 469152 3292 469216 3296
rect 469152 3236 469156 3292
rect 469156 3236 469212 3292
rect 469212 3236 469216 3292
rect 469152 3232 469216 3236
rect 469232 3292 469296 3296
rect 469232 3236 469236 3292
rect 469236 3236 469292 3292
rect 469292 3236 469296 3292
rect 469232 3232 469296 3236
rect 469312 3292 469376 3296
rect 469312 3236 469316 3292
rect 469316 3236 469372 3292
rect 469372 3236 469376 3292
rect 469312 3232 469376 3236
rect 504832 3292 504896 3296
rect 504832 3236 504836 3292
rect 504836 3236 504892 3292
rect 504892 3236 504896 3292
rect 504832 3232 504896 3236
rect 504912 3292 504976 3296
rect 504912 3236 504916 3292
rect 504916 3236 504972 3292
rect 504972 3236 504976 3292
rect 504912 3232 504976 3236
rect 504992 3292 505056 3296
rect 504992 3236 504996 3292
rect 504996 3236 505052 3292
rect 505052 3236 505056 3292
rect 504992 3232 505056 3236
rect 505072 3292 505136 3296
rect 505072 3236 505076 3292
rect 505076 3236 505132 3292
rect 505132 3236 505136 3292
rect 505072 3232 505136 3236
rect 505152 3292 505216 3296
rect 505152 3236 505156 3292
rect 505156 3236 505212 3292
rect 505212 3236 505216 3292
rect 505152 3232 505216 3236
rect 505232 3292 505296 3296
rect 505232 3236 505236 3292
rect 505236 3236 505292 3292
rect 505292 3236 505296 3292
rect 505232 3232 505296 3236
rect 505312 3292 505376 3296
rect 505312 3236 505316 3292
rect 505316 3236 505372 3292
rect 505372 3236 505376 3292
rect 505312 3232 505376 3236
rect 540832 3292 540896 3296
rect 540832 3236 540836 3292
rect 540836 3236 540892 3292
rect 540892 3236 540896 3292
rect 540832 3232 540896 3236
rect 540912 3292 540976 3296
rect 540912 3236 540916 3292
rect 540916 3236 540972 3292
rect 540972 3236 540976 3292
rect 540912 3232 540976 3236
rect 540992 3292 541056 3296
rect 540992 3236 540996 3292
rect 540996 3236 541052 3292
rect 541052 3236 541056 3292
rect 540992 3232 541056 3236
rect 541072 3292 541136 3296
rect 541072 3236 541076 3292
rect 541076 3236 541132 3292
rect 541132 3236 541136 3292
rect 541072 3232 541136 3236
rect 541152 3292 541216 3296
rect 541152 3236 541156 3292
rect 541156 3236 541212 3292
rect 541212 3236 541216 3292
rect 541152 3232 541216 3236
rect 541232 3292 541296 3296
rect 541232 3236 541236 3292
rect 541236 3236 541292 3292
rect 541292 3236 541296 3292
rect 541232 3232 541296 3236
rect 541312 3292 541376 3296
rect 541312 3236 541316 3292
rect 541316 3236 541372 3292
rect 541372 3236 541376 3292
rect 541312 3232 541376 3236
rect 576832 3292 576896 3296
rect 576832 3236 576836 3292
rect 576836 3236 576892 3292
rect 576892 3236 576896 3292
rect 576832 3232 576896 3236
rect 576912 3292 576976 3296
rect 576912 3236 576916 3292
rect 576916 3236 576972 3292
rect 576972 3236 576976 3292
rect 576912 3232 576976 3236
rect 576992 3292 577056 3296
rect 576992 3236 576996 3292
rect 576996 3236 577052 3292
rect 577052 3236 577056 3292
rect 576992 3232 577056 3236
rect 577072 3292 577136 3296
rect 577072 3236 577076 3292
rect 577076 3236 577132 3292
rect 577132 3236 577136 3292
rect 577072 3232 577136 3236
rect 577152 3292 577216 3296
rect 577152 3236 577156 3292
rect 577156 3236 577212 3292
rect 577212 3236 577216 3292
rect 577152 3232 577216 3236
rect 577232 3292 577296 3296
rect 577232 3236 577236 3292
rect 577236 3236 577292 3292
rect 577292 3236 577296 3292
rect 577232 3232 577296 3236
rect 577312 3292 577376 3296
rect 577312 3236 577316 3292
rect 577316 3236 577372 3292
rect 577372 3236 577376 3292
rect 577312 3232 577376 3236
rect 18832 2748 18896 2752
rect 18832 2692 18836 2748
rect 18836 2692 18892 2748
rect 18892 2692 18896 2748
rect 18832 2688 18896 2692
rect 18912 2748 18976 2752
rect 18912 2692 18916 2748
rect 18916 2692 18972 2748
rect 18972 2692 18976 2748
rect 18912 2688 18976 2692
rect 18992 2748 19056 2752
rect 18992 2692 18996 2748
rect 18996 2692 19052 2748
rect 19052 2692 19056 2748
rect 18992 2688 19056 2692
rect 19072 2748 19136 2752
rect 19072 2692 19076 2748
rect 19076 2692 19132 2748
rect 19132 2692 19136 2748
rect 19072 2688 19136 2692
rect 19152 2748 19216 2752
rect 19152 2692 19156 2748
rect 19156 2692 19212 2748
rect 19212 2692 19216 2748
rect 19152 2688 19216 2692
rect 19232 2748 19296 2752
rect 19232 2692 19236 2748
rect 19236 2692 19292 2748
rect 19292 2692 19296 2748
rect 19232 2688 19296 2692
rect 19312 2748 19376 2752
rect 19312 2692 19316 2748
rect 19316 2692 19372 2748
rect 19372 2692 19376 2748
rect 19312 2688 19376 2692
rect 54832 2748 54896 2752
rect 54832 2692 54836 2748
rect 54836 2692 54892 2748
rect 54892 2692 54896 2748
rect 54832 2688 54896 2692
rect 54912 2748 54976 2752
rect 54912 2692 54916 2748
rect 54916 2692 54972 2748
rect 54972 2692 54976 2748
rect 54912 2688 54976 2692
rect 54992 2748 55056 2752
rect 54992 2692 54996 2748
rect 54996 2692 55052 2748
rect 55052 2692 55056 2748
rect 54992 2688 55056 2692
rect 55072 2748 55136 2752
rect 55072 2692 55076 2748
rect 55076 2692 55132 2748
rect 55132 2692 55136 2748
rect 55072 2688 55136 2692
rect 55152 2748 55216 2752
rect 55152 2692 55156 2748
rect 55156 2692 55212 2748
rect 55212 2692 55216 2748
rect 55152 2688 55216 2692
rect 55232 2748 55296 2752
rect 55232 2692 55236 2748
rect 55236 2692 55292 2748
rect 55292 2692 55296 2748
rect 55232 2688 55296 2692
rect 55312 2748 55376 2752
rect 55312 2692 55316 2748
rect 55316 2692 55372 2748
rect 55372 2692 55376 2748
rect 55312 2688 55376 2692
rect 90832 2748 90896 2752
rect 90832 2692 90836 2748
rect 90836 2692 90892 2748
rect 90892 2692 90896 2748
rect 90832 2688 90896 2692
rect 90912 2748 90976 2752
rect 90912 2692 90916 2748
rect 90916 2692 90972 2748
rect 90972 2692 90976 2748
rect 90912 2688 90976 2692
rect 90992 2748 91056 2752
rect 90992 2692 90996 2748
rect 90996 2692 91052 2748
rect 91052 2692 91056 2748
rect 90992 2688 91056 2692
rect 91072 2748 91136 2752
rect 91072 2692 91076 2748
rect 91076 2692 91132 2748
rect 91132 2692 91136 2748
rect 91072 2688 91136 2692
rect 91152 2748 91216 2752
rect 91152 2692 91156 2748
rect 91156 2692 91212 2748
rect 91212 2692 91216 2748
rect 91152 2688 91216 2692
rect 91232 2748 91296 2752
rect 91232 2692 91236 2748
rect 91236 2692 91292 2748
rect 91292 2692 91296 2748
rect 91232 2688 91296 2692
rect 91312 2748 91376 2752
rect 91312 2692 91316 2748
rect 91316 2692 91372 2748
rect 91372 2692 91376 2748
rect 91312 2688 91376 2692
rect 126832 2748 126896 2752
rect 126832 2692 126836 2748
rect 126836 2692 126892 2748
rect 126892 2692 126896 2748
rect 126832 2688 126896 2692
rect 126912 2748 126976 2752
rect 126912 2692 126916 2748
rect 126916 2692 126972 2748
rect 126972 2692 126976 2748
rect 126912 2688 126976 2692
rect 126992 2748 127056 2752
rect 126992 2692 126996 2748
rect 126996 2692 127052 2748
rect 127052 2692 127056 2748
rect 126992 2688 127056 2692
rect 127072 2748 127136 2752
rect 127072 2692 127076 2748
rect 127076 2692 127132 2748
rect 127132 2692 127136 2748
rect 127072 2688 127136 2692
rect 127152 2748 127216 2752
rect 127152 2692 127156 2748
rect 127156 2692 127212 2748
rect 127212 2692 127216 2748
rect 127152 2688 127216 2692
rect 127232 2748 127296 2752
rect 127232 2692 127236 2748
rect 127236 2692 127292 2748
rect 127292 2692 127296 2748
rect 127232 2688 127296 2692
rect 127312 2748 127376 2752
rect 127312 2692 127316 2748
rect 127316 2692 127372 2748
rect 127372 2692 127376 2748
rect 127312 2688 127376 2692
rect 162832 2748 162896 2752
rect 162832 2692 162836 2748
rect 162836 2692 162892 2748
rect 162892 2692 162896 2748
rect 162832 2688 162896 2692
rect 162912 2748 162976 2752
rect 162912 2692 162916 2748
rect 162916 2692 162972 2748
rect 162972 2692 162976 2748
rect 162912 2688 162976 2692
rect 162992 2748 163056 2752
rect 162992 2692 162996 2748
rect 162996 2692 163052 2748
rect 163052 2692 163056 2748
rect 162992 2688 163056 2692
rect 163072 2748 163136 2752
rect 163072 2692 163076 2748
rect 163076 2692 163132 2748
rect 163132 2692 163136 2748
rect 163072 2688 163136 2692
rect 163152 2748 163216 2752
rect 163152 2692 163156 2748
rect 163156 2692 163212 2748
rect 163212 2692 163216 2748
rect 163152 2688 163216 2692
rect 163232 2748 163296 2752
rect 163232 2692 163236 2748
rect 163236 2692 163292 2748
rect 163292 2692 163296 2748
rect 163232 2688 163296 2692
rect 163312 2748 163376 2752
rect 163312 2692 163316 2748
rect 163316 2692 163372 2748
rect 163372 2692 163376 2748
rect 163312 2688 163376 2692
rect 198832 2748 198896 2752
rect 198832 2692 198836 2748
rect 198836 2692 198892 2748
rect 198892 2692 198896 2748
rect 198832 2688 198896 2692
rect 198912 2748 198976 2752
rect 198912 2692 198916 2748
rect 198916 2692 198972 2748
rect 198972 2692 198976 2748
rect 198912 2688 198976 2692
rect 198992 2748 199056 2752
rect 198992 2692 198996 2748
rect 198996 2692 199052 2748
rect 199052 2692 199056 2748
rect 198992 2688 199056 2692
rect 199072 2748 199136 2752
rect 199072 2692 199076 2748
rect 199076 2692 199132 2748
rect 199132 2692 199136 2748
rect 199072 2688 199136 2692
rect 199152 2748 199216 2752
rect 199152 2692 199156 2748
rect 199156 2692 199212 2748
rect 199212 2692 199216 2748
rect 199152 2688 199216 2692
rect 199232 2748 199296 2752
rect 199232 2692 199236 2748
rect 199236 2692 199292 2748
rect 199292 2692 199296 2748
rect 199232 2688 199296 2692
rect 199312 2748 199376 2752
rect 199312 2692 199316 2748
rect 199316 2692 199372 2748
rect 199372 2692 199376 2748
rect 199312 2688 199376 2692
rect 234832 2748 234896 2752
rect 234832 2692 234836 2748
rect 234836 2692 234892 2748
rect 234892 2692 234896 2748
rect 234832 2688 234896 2692
rect 234912 2748 234976 2752
rect 234912 2692 234916 2748
rect 234916 2692 234972 2748
rect 234972 2692 234976 2748
rect 234912 2688 234976 2692
rect 234992 2748 235056 2752
rect 234992 2692 234996 2748
rect 234996 2692 235052 2748
rect 235052 2692 235056 2748
rect 234992 2688 235056 2692
rect 235072 2748 235136 2752
rect 235072 2692 235076 2748
rect 235076 2692 235132 2748
rect 235132 2692 235136 2748
rect 235072 2688 235136 2692
rect 235152 2748 235216 2752
rect 235152 2692 235156 2748
rect 235156 2692 235212 2748
rect 235212 2692 235216 2748
rect 235152 2688 235216 2692
rect 235232 2748 235296 2752
rect 235232 2692 235236 2748
rect 235236 2692 235292 2748
rect 235292 2692 235296 2748
rect 235232 2688 235296 2692
rect 235312 2748 235376 2752
rect 235312 2692 235316 2748
rect 235316 2692 235372 2748
rect 235372 2692 235376 2748
rect 235312 2688 235376 2692
rect 270832 2748 270896 2752
rect 270832 2692 270836 2748
rect 270836 2692 270892 2748
rect 270892 2692 270896 2748
rect 270832 2688 270896 2692
rect 270912 2748 270976 2752
rect 270912 2692 270916 2748
rect 270916 2692 270972 2748
rect 270972 2692 270976 2748
rect 270912 2688 270976 2692
rect 270992 2748 271056 2752
rect 270992 2692 270996 2748
rect 270996 2692 271052 2748
rect 271052 2692 271056 2748
rect 270992 2688 271056 2692
rect 271072 2748 271136 2752
rect 271072 2692 271076 2748
rect 271076 2692 271132 2748
rect 271132 2692 271136 2748
rect 271072 2688 271136 2692
rect 271152 2748 271216 2752
rect 271152 2692 271156 2748
rect 271156 2692 271212 2748
rect 271212 2692 271216 2748
rect 271152 2688 271216 2692
rect 271232 2748 271296 2752
rect 271232 2692 271236 2748
rect 271236 2692 271292 2748
rect 271292 2692 271296 2748
rect 271232 2688 271296 2692
rect 271312 2748 271376 2752
rect 271312 2692 271316 2748
rect 271316 2692 271372 2748
rect 271372 2692 271376 2748
rect 271312 2688 271376 2692
rect 306832 2748 306896 2752
rect 306832 2692 306836 2748
rect 306836 2692 306892 2748
rect 306892 2692 306896 2748
rect 306832 2688 306896 2692
rect 306912 2748 306976 2752
rect 306912 2692 306916 2748
rect 306916 2692 306972 2748
rect 306972 2692 306976 2748
rect 306912 2688 306976 2692
rect 306992 2748 307056 2752
rect 306992 2692 306996 2748
rect 306996 2692 307052 2748
rect 307052 2692 307056 2748
rect 306992 2688 307056 2692
rect 307072 2748 307136 2752
rect 307072 2692 307076 2748
rect 307076 2692 307132 2748
rect 307132 2692 307136 2748
rect 307072 2688 307136 2692
rect 307152 2748 307216 2752
rect 307152 2692 307156 2748
rect 307156 2692 307212 2748
rect 307212 2692 307216 2748
rect 307152 2688 307216 2692
rect 307232 2748 307296 2752
rect 307232 2692 307236 2748
rect 307236 2692 307292 2748
rect 307292 2692 307296 2748
rect 307232 2688 307296 2692
rect 307312 2748 307376 2752
rect 307312 2692 307316 2748
rect 307316 2692 307372 2748
rect 307372 2692 307376 2748
rect 307312 2688 307376 2692
rect 342832 2748 342896 2752
rect 342832 2692 342836 2748
rect 342836 2692 342892 2748
rect 342892 2692 342896 2748
rect 342832 2688 342896 2692
rect 342912 2748 342976 2752
rect 342912 2692 342916 2748
rect 342916 2692 342972 2748
rect 342972 2692 342976 2748
rect 342912 2688 342976 2692
rect 342992 2748 343056 2752
rect 342992 2692 342996 2748
rect 342996 2692 343052 2748
rect 343052 2692 343056 2748
rect 342992 2688 343056 2692
rect 343072 2748 343136 2752
rect 343072 2692 343076 2748
rect 343076 2692 343132 2748
rect 343132 2692 343136 2748
rect 343072 2688 343136 2692
rect 343152 2748 343216 2752
rect 343152 2692 343156 2748
rect 343156 2692 343212 2748
rect 343212 2692 343216 2748
rect 343152 2688 343216 2692
rect 343232 2748 343296 2752
rect 343232 2692 343236 2748
rect 343236 2692 343292 2748
rect 343292 2692 343296 2748
rect 343232 2688 343296 2692
rect 343312 2748 343376 2752
rect 343312 2692 343316 2748
rect 343316 2692 343372 2748
rect 343372 2692 343376 2748
rect 343312 2688 343376 2692
rect 378832 2748 378896 2752
rect 378832 2692 378836 2748
rect 378836 2692 378892 2748
rect 378892 2692 378896 2748
rect 378832 2688 378896 2692
rect 378912 2748 378976 2752
rect 378912 2692 378916 2748
rect 378916 2692 378972 2748
rect 378972 2692 378976 2748
rect 378912 2688 378976 2692
rect 378992 2748 379056 2752
rect 378992 2692 378996 2748
rect 378996 2692 379052 2748
rect 379052 2692 379056 2748
rect 378992 2688 379056 2692
rect 379072 2748 379136 2752
rect 379072 2692 379076 2748
rect 379076 2692 379132 2748
rect 379132 2692 379136 2748
rect 379072 2688 379136 2692
rect 379152 2748 379216 2752
rect 379152 2692 379156 2748
rect 379156 2692 379212 2748
rect 379212 2692 379216 2748
rect 379152 2688 379216 2692
rect 379232 2748 379296 2752
rect 379232 2692 379236 2748
rect 379236 2692 379292 2748
rect 379292 2692 379296 2748
rect 379232 2688 379296 2692
rect 379312 2748 379376 2752
rect 379312 2692 379316 2748
rect 379316 2692 379372 2748
rect 379372 2692 379376 2748
rect 379312 2688 379376 2692
rect 414832 2748 414896 2752
rect 414832 2692 414836 2748
rect 414836 2692 414892 2748
rect 414892 2692 414896 2748
rect 414832 2688 414896 2692
rect 414912 2748 414976 2752
rect 414912 2692 414916 2748
rect 414916 2692 414972 2748
rect 414972 2692 414976 2748
rect 414912 2688 414976 2692
rect 414992 2748 415056 2752
rect 414992 2692 414996 2748
rect 414996 2692 415052 2748
rect 415052 2692 415056 2748
rect 414992 2688 415056 2692
rect 415072 2748 415136 2752
rect 415072 2692 415076 2748
rect 415076 2692 415132 2748
rect 415132 2692 415136 2748
rect 415072 2688 415136 2692
rect 415152 2748 415216 2752
rect 415152 2692 415156 2748
rect 415156 2692 415212 2748
rect 415212 2692 415216 2748
rect 415152 2688 415216 2692
rect 415232 2748 415296 2752
rect 415232 2692 415236 2748
rect 415236 2692 415292 2748
rect 415292 2692 415296 2748
rect 415232 2688 415296 2692
rect 415312 2748 415376 2752
rect 415312 2692 415316 2748
rect 415316 2692 415372 2748
rect 415372 2692 415376 2748
rect 415312 2688 415376 2692
rect 450832 2748 450896 2752
rect 450832 2692 450836 2748
rect 450836 2692 450892 2748
rect 450892 2692 450896 2748
rect 450832 2688 450896 2692
rect 450912 2748 450976 2752
rect 450912 2692 450916 2748
rect 450916 2692 450972 2748
rect 450972 2692 450976 2748
rect 450912 2688 450976 2692
rect 450992 2748 451056 2752
rect 450992 2692 450996 2748
rect 450996 2692 451052 2748
rect 451052 2692 451056 2748
rect 450992 2688 451056 2692
rect 451072 2748 451136 2752
rect 451072 2692 451076 2748
rect 451076 2692 451132 2748
rect 451132 2692 451136 2748
rect 451072 2688 451136 2692
rect 451152 2748 451216 2752
rect 451152 2692 451156 2748
rect 451156 2692 451212 2748
rect 451212 2692 451216 2748
rect 451152 2688 451216 2692
rect 451232 2748 451296 2752
rect 451232 2692 451236 2748
rect 451236 2692 451292 2748
rect 451292 2692 451296 2748
rect 451232 2688 451296 2692
rect 451312 2748 451376 2752
rect 451312 2692 451316 2748
rect 451316 2692 451372 2748
rect 451372 2692 451376 2748
rect 451312 2688 451376 2692
rect 486832 2748 486896 2752
rect 486832 2692 486836 2748
rect 486836 2692 486892 2748
rect 486892 2692 486896 2748
rect 486832 2688 486896 2692
rect 486912 2748 486976 2752
rect 486912 2692 486916 2748
rect 486916 2692 486972 2748
rect 486972 2692 486976 2748
rect 486912 2688 486976 2692
rect 486992 2748 487056 2752
rect 486992 2692 486996 2748
rect 486996 2692 487052 2748
rect 487052 2692 487056 2748
rect 486992 2688 487056 2692
rect 487072 2748 487136 2752
rect 487072 2692 487076 2748
rect 487076 2692 487132 2748
rect 487132 2692 487136 2748
rect 487072 2688 487136 2692
rect 487152 2748 487216 2752
rect 487152 2692 487156 2748
rect 487156 2692 487212 2748
rect 487212 2692 487216 2748
rect 487152 2688 487216 2692
rect 487232 2748 487296 2752
rect 487232 2692 487236 2748
rect 487236 2692 487292 2748
rect 487292 2692 487296 2748
rect 487232 2688 487296 2692
rect 487312 2748 487376 2752
rect 487312 2692 487316 2748
rect 487316 2692 487372 2748
rect 487372 2692 487376 2748
rect 487312 2688 487376 2692
rect 522832 2748 522896 2752
rect 522832 2692 522836 2748
rect 522836 2692 522892 2748
rect 522892 2692 522896 2748
rect 522832 2688 522896 2692
rect 522912 2748 522976 2752
rect 522912 2692 522916 2748
rect 522916 2692 522972 2748
rect 522972 2692 522976 2748
rect 522912 2688 522976 2692
rect 522992 2748 523056 2752
rect 522992 2692 522996 2748
rect 522996 2692 523052 2748
rect 523052 2692 523056 2748
rect 522992 2688 523056 2692
rect 523072 2748 523136 2752
rect 523072 2692 523076 2748
rect 523076 2692 523132 2748
rect 523132 2692 523136 2748
rect 523072 2688 523136 2692
rect 523152 2748 523216 2752
rect 523152 2692 523156 2748
rect 523156 2692 523212 2748
rect 523212 2692 523216 2748
rect 523152 2688 523216 2692
rect 523232 2748 523296 2752
rect 523232 2692 523236 2748
rect 523236 2692 523292 2748
rect 523292 2692 523296 2748
rect 523232 2688 523296 2692
rect 523312 2748 523376 2752
rect 523312 2692 523316 2748
rect 523316 2692 523372 2748
rect 523372 2692 523376 2748
rect 523312 2688 523376 2692
rect 558832 2748 558896 2752
rect 558832 2692 558836 2748
rect 558836 2692 558892 2748
rect 558892 2692 558896 2748
rect 558832 2688 558896 2692
rect 558912 2748 558976 2752
rect 558912 2692 558916 2748
rect 558916 2692 558972 2748
rect 558972 2692 558976 2748
rect 558912 2688 558976 2692
rect 558992 2748 559056 2752
rect 558992 2692 558996 2748
rect 558996 2692 559052 2748
rect 559052 2692 559056 2748
rect 558992 2688 559056 2692
rect 559072 2748 559136 2752
rect 559072 2692 559076 2748
rect 559076 2692 559132 2748
rect 559132 2692 559136 2748
rect 559072 2688 559136 2692
rect 559152 2748 559216 2752
rect 559152 2692 559156 2748
rect 559156 2692 559212 2748
rect 559212 2692 559216 2748
rect 559152 2688 559216 2692
rect 559232 2748 559296 2752
rect 559232 2692 559236 2748
rect 559236 2692 559292 2748
rect 559292 2692 559296 2748
rect 559232 2688 559296 2692
rect 559312 2748 559376 2752
rect 559312 2692 559316 2748
rect 559316 2692 559372 2748
rect 559372 2692 559376 2748
rect 559312 2688 559376 2692
rect 36832 2204 36896 2208
rect 36832 2148 36836 2204
rect 36836 2148 36892 2204
rect 36892 2148 36896 2204
rect 36832 2144 36896 2148
rect 36912 2204 36976 2208
rect 36912 2148 36916 2204
rect 36916 2148 36972 2204
rect 36972 2148 36976 2204
rect 36912 2144 36976 2148
rect 36992 2204 37056 2208
rect 36992 2148 36996 2204
rect 36996 2148 37052 2204
rect 37052 2148 37056 2204
rect 36992 2144 37056 2148
rect 37072 2204 37136 2208
rect 37072 2148 37076 2204
rect 37076 2148 37132 2204
rect 37132 2148 37136 2204
rect 37072 2144 37136 2148
rect 37152 2204 37216 2208
rect 37152 2148 37156 2204
rect 37156 2148 37212 2204
rect 37212 2148 37216 2204
rect 37152 2144 37216 2148
rect 37232 2204 37296 2208
rect 37232 2148 37236 2204
rect 37236 2148 37292 2204
rect 37292 2148 37296 2204
rect 37232 2144 37296 2148
rect 37312 2204 37376 2208
rect 37312 2148 37316 2204
rect 37316 2148 37372 2204
rect 37372 2148 37376 2204
rect 37312 2144 37376 2148
rect 72832 2204 72896 2208
rect 72832 2148 72836 2204
rect 72836 2148 72892 2204
rect 72892 2148 72896 2204
rect 72832 2144 72896 2148
rect 72912 2204 72976 2208
rect 72912 2148 72916 2204
rect 72916 2148 72972 2204
rect 72972 2148 72976 2204
rect 72912 2144 72976 2148
rect 72992 2204 73056 2208
rect 72992 2148 72996 2204
rect 72996 2148 73052 2204
rect 73052 2148 73056 2204
rect 72992 2144 73056 2148
rect 73072 2204 73136 2208
rect 73072 2148 73076 2204
rect 73076 2148 73132 2204
rect 73132 2148 73136 2204
rect 73072 2144 73136 2148
rect 73152 2204 73216 2208
rect 73152 2148 73156 2204
rect 73156 2148 73212 2204
rect 73212 2148 73216 2204
rect 73152 2144 73216 2148
rect 73232 2204 73296 2208
rect 73232 2148 73236 2204
rect 73236 2148 73292 2204
rect 73292 2148 73296 2204
rect 73232 2144 73296 2148
rect 73312 2204 73376 2208
rect 73312 2148 73316 2204
rect 73316 2148 73372 2204
rect 73372 2148 73376 2204
rect 73312 2144 73376 2148
rect 108832 2204 108896 2208
rect 108832 2148 108836 2204
rect 108836 2148 108892 2204
rect 108892 2148 108896 2204
rect 108832 2144 108896 2148
rect 108912 2204 108976 2208
rect 108912 2148 108916 2204
rect 108916 2148 108972 2204
rect 108972 2148 108976 2204
rect 108912 2144 108976 2148
rect 108992 2204 109056 2208
rect 108992 2148 108996 2204
rect 108996 2148 109052 2204
rect 109052 2148 109056 2204
rect 108992 2144 109056 2148
rect 109072 2204 109136 2208
rect 109072 2148 109076 2204
rect 109076 2148 109132 2204
rect 109132 2148 109136 2204
rect 109072 2144 109136 2148
rect 109152 2204 109216 2208
rect 109152 2148 109156 2204
rect 109156 2148 109212 2204
rect 109212 2148 109216 2204
rect 109152 2144 109216 2148
rect 109232 2204 109296 2208
rect 109232 2148 109236 2204
rect 109236 2148 109292 2204
rect 109292 2148 109296 2204
rect 109232 2144 109296 2148
rect 109312 2204 109376 2208
rect 109312 2148 109316 2204
rect 109316 2148 109372 2204
rect 109372 2148 109376 2204
rect 109312 2144 109376 2148
rect 144832 2204 144896 2208
rect 144832 2148 144836 2204
rect 144836 2148 144892 2204
rect 144892 2148 144896 2204
rect 144832 2144 144896 2148
rect 144912 2204 144976 2208
rect 144912 2148 144916 2204
rect 144916 2148 144972 2204
rect 144972 2148 144976 2204
rect 144912 2144 144976 2148
rect 144992 2204 145056 2208
rect 144992 2148 144996 2204
rect 144996 2148 145052 2204
rect 145052 2148 145056 2204
rect 144992 2144 145056 2148
rect 145072 2204 145136 2208
rect 145072 2148 145076 2204
rect 145076 2148 145132 2204
rect 145132 2148 145136 2204
rect 145072 2144 145136 2148
rect 145152 2204 145216 2208
rect 145152 2148 145156 2204
rect 145156 2148 145212 2204
rect 145212 2148 145216 2204
rect 145152 2144 145216 2148
rect 145232 2204 145296 2208
rect 145232 2148 145236 2204
rect 145236 2148 145292 2204
rect 145292 2148 145296 2204
rect 145232 2144 145296 2148
rect 145312 2204 145376 2208
rect 145312 2148 145316 2204
rect 145316 2148 145372 2204
rect 145372 2148 145376 2204
rect 145312 2144 145376 2148
rect 180832 2204 180896 2208
rect 180832 2148 180836 2204
rect 180836 2148 180892 2204
rect 180892 2148 180896 2204
rect 180832 2144 180896 2148
rect 180912 2204 180976 2208
rect 180912 2148 180916 2204
rect 180916 2148 180972 2204
rect 180972 2148 180976 2204
rect 180912 2144 180976 2148
rect 180992 2204 181056 2208
rect 180992 2148 180996 2204
rect 180996 2148 181052 2204
rect 181052 2148 181056 2204
rect 180992 2144 181056 2148
rect 181072 2204 181136 2208
rect 181072 2148 181076 2204
rect 181076 2148 181132 2204
rect 181132 2148 181136 2204
rect 181072 2144 181136 2148
rect 181152 2204 181216 2208
rect 181152 2148 181156 2204
rect 181156 2148 181212 2204
rect 181212 2148 181216 2204
rect 181152 2144 181216 2148
rect 181232 2204 181296 2208
rect 181232 2148 181236 2204
rect 181236 2148 181292 2204
rect 181292 2148 181296 2204
rect 181232 2144 181296 2148
rect 181312 2204 181376 2208
rect 181312 2148 181316 2204
rect 181316 2148 181372 2204
rect 181372 2148 181376 2204
rect 181312 2144 181376 2148
rect 216832 2204 216896 2208
rect 216832 2148 216836 2204
rect 216836 2148 216892 2204
rect 216892 2148 216896 2204
rect 216832 2144 216896 2148
rect 216912 2204 216976 2208
rect 216912 2148 216916 2204
rect 216916 2148 216972 2204
rect 216972 2148 216976 2204
rect 216912 2144 216976 2148
rect 216992 2204 217056 2208
rect 216992 2148 216996 2204
rect 216996 2148 217052 2204
rect 217052 2148 217056 2204
rect 216992 2144 217056 2148
rect 217072 2204 217136 2208
rect 217072 2148 217076 2204
rect 217076 2148 217132 2204
rect 217132 2148 217136 2204
rect 217072 2144 217136 2148
rect 217152 2204 217216 2208
rect 217152 2148 217156 2204
rect 217156 2148 217212 2204
rect 217212 2148 217216 2204
rect 217152 2144 217216 2148
rect 217232 2204 217296 2208
rect 217232 2148 217236 2204
rect 217236 2148 217292 2204
rect 217292 2148 217296 2204
rect 217232 2144 217296 2148
rect 217312 2204 217376 2208
rect 217312 2148 217316 2204
rect 217316 2148 217372 2204
rect 217372 2148 217376 2204
rect 217312 2144 217376 2148
rect 252832 2204 252896 2208
rect 252832 2148 252836 2204
rect 252836 2148 252892 2204
rect 252892 2148 252896 2204
rect 252832 2144 252896 2148
rect 252912 2204 252976 2208
rect 252912 2148 252916 2204
rect 252916 2148 252972 2204
rect 252972 2148 252976 2204
rect 252912 2144 252976 2148
rect 252992 2204 253056 2208
rect 252992 2148 252996 2204
rect 252996 2148 253052 2204
rect 253052 2148 253056 2204
rect 252992 2144 253056 2148
rect 253072 2204 253136 2208
rect 253072 2148 253076 2204
rect 253076 2148 253132 2204
rect 253132 2148 253136 2204
rect 253072 2144 253136 2148
rect 253152 2204 253216 2208
rect 253152 2148 253156 2204
rect 253156 2148 253212 2204
rect 253212 2148 253216 2204
rect 253152 2144 253216 2148
rect 253232 2204 253296 2208
rect 253232 2148 253236 2204
rect 253236 2148 253292 2204
rect 253292 2148 253296 2204
rect 253232 2144 253296 2148
rect 253312 2204 253376 2208
rect 253312 2148 253316 2204
rect 253316 2148 253372 2204
rect 253372 2148 253376 2204
rect 253312 2144 253376 2148
rect 288832 2204 288896 2208
rect 288832 2148 288836 2204
rect 288836 2148 288892 2204
rect 288892 2148 288896 2204
rect 288832 2144 288896 2148
rect 288912 2204 288976 2208
rect 288912 2148 288916 2204
rect 288916 2148 288972 2204
rect 288972 2148 288976 2204
rect 288912 2144 288976 2148
rect 288992 2204 289056 2208
rect 288992 2148 288996 2204
rect 288996 2148 289052 2204
rect 289052 2148 289056 2204
rect 288992 2144 289056 2148
rect 289072 2204 289136 2208
rect 289072 2148 289076 2204
rect 289076 2148 289132 2204
rect 289132 2148 289136 2204
rect 289072 2144 289136 2148
rect 289152 2204 289216 2208
rect 289152 2148 289156 2204
rect 289156 2148 289212 2204
rect 289212 2148 289216 2204
rect 289152 2144 289216 2148
rect 289232 2204 289296 2208
rect 289232 2148 289236 2204
rect 289236 2148 289292 2204
rect 289292 2148 289296 2204
rect 289232 2144 289296 2148
rect 289312 2204 289376 2208
rect 289312 2148 289316 2204
rect 289316 2148 289372 2204
rect 289372 2148 289376 2204
rect 289312 2144 289376 2148
rect 324832 2204 324896 2208
rect 324832 2148 324836 2204
rect 324836 2148 324892 2204
rect 324892 2148 324896 2204
rect 324832 2144 324896 2148
rect 324912 2204 324976 2208
rect 324912 2148 324916 2204
rect 324916 2148 324972 2204
rect 324972 2148 324976 2204
rect 324912 2144 324976 2148
rect 324992 2204 325056 2208
rect 324992 2148 324996 2204
rect 324996 2148 325052 2204
rect 325052 2148 325056 2204
rect 324992 2144 325056 2148
rect 325072 2204 325136 2208
rect 325072 2148 325076 2204
rect 325076 2148 325132 2204
rect 325132 2148 325136 2204
rect 325072 2144 325136 2148
rect 325152 2204 325216 2208
rect 325152 2148 325156 2204
rect 325156 2148 325212 2204
rect 325212 2148 325216 2204
rect 325152 2144 325216 2148
rect 325232 2204 325296 2208
rect 325232 2148 325236 2204
rect 325236 2148 325292 2204
rect 325292 2148 325296 2204
rect 325232 2144 325296 2148
rect 325312 2204 325376 2208
rect 325312 2148 325316 2204
rect 325316 2148 325372 2204
rect 325372 2148 325376 2204
rect 325312 2144 325376 2148
rect 360832 2204 360896 2208
rect 360832 2148 360836 2204
rect 360836 2148 360892 2204
rect 360892 2148 360896 2204
rect 360832 2144 360896 2148
rect 360912 2204 360976 2208
rect 360912 2148 360916 2204
rect 360916 2148 360972 2204
rect 360972 2148 360976 2204
rect 360912 2144 360976 2148
rect 360992 2204 361056 2208
rect 360992 2148 360996 2204
rect 360996 2148 361052 2204
rect 361052 2148 361056 2204
rect 360992 2144 361056 2148
rect 361072 2204 361136 2208
rect 361072 2148 361076 2204
rect 361076 2148 361132 2204
rect 361132 2148 361136 2204
rect 361072 2144 361136 2148
rect 361152 2204 361216 2208
rect 361152 2148 361156 2204
rect 361156 2148 361212 2204
rect 361212 2148 361216 2204
rect 361152 2144 361216 2148
rect 361232 2204 361296 2208
rect 361232 2148 361236 2204
rect 361236 2148 361292 2204
rect 361292 2148 361296 2204
rect 361232 2144 361296 2148
rect 361312 2204 361376 2208
rect 361312 2148 361316 2204
rect 361316 2148 361372 2204
rect 361372 2148 361376 2204
rect 361312 2144 361376 2148
rect 396832 2204 396896 2208
rect 396832 2148 396836 2204
rect 396836 2148 396892 2204
rect 396892 2148 396896 2204
rect 396832 2144 396896 2148
rect 396912 2204 396976 2208
rect 396912 2148 396916 2204
rect 396916 2148 396972 2204
rect 396972 2148 396976 2204
rect 396912 2144 396976 2148
rect 396992 2204 397056 2208
rect 396992 2148 396996 2204
rect 396996 2148 397052 2204
rect 397052 2148 397056 2204
rect 396992 2144 397056 2148
rect 397072 2204 397136 2208
rect 397072 2148 397076 2204
rect 397076 2148 397132 2204
rect 397132 2148 397136 2204
rect 397072 2144 397136 2148
rect 397152 2204 397216 2208
rect 397152 2148 397156 2204
rect 397156 2148 397212 2204
rect 397212 2148 397216 2204
rect 397152 2144 397216 2148
rect 397232 2204 397296 2208
rect 397232 2148 397236 2204
rect 397236 2148 397292 2204
rect 397292 2148 397296 2204
rect 397232 2144 397296 2148
rect 397312 2204 397376 2208
rect 397312 2148 397316 2204
rect 397316 2148 397372 2204
rect 397372 2148 397376 2204
rect 397312 2144 397376 2148
rect 432832 2204 432896 2208
rect 432832 2148 432836 2204
rect 432836 2148 432892 2204
rect 432892 2148 432896 2204
rect 432832 2144 432896 2148
rect 432912 2204 432976 2208
rect 432912 2148 432916 2204
rect 432916 2148 432972 2204
rect 432972 2148 432976 2204
rect 432912 2144 432976 2148
rect 432992 2204 433056 2208
rect 432992 2148 432996 2204
rect 432996 2148 433052 2204
rect 433052 2148 433056 2204
rect 432992 2144 433056 2148
rect 433072 2204 433136 2208
rect 433072 2148 433076 2204
rect 433076 2148 433132 2204
rect 433132 2148 433136 2204
rect 433072 2144 433136 2148
rect 433152 2204 433216 2208
rect 433152 2148 433156 2204
rect 433156 2148 433212 2204
rect 433212 2148 433216 2204
rect 433152 2144 433216 2148
rect 433232 2204 433296 2208
rect 433232 2148 433236 2204
rect 433236 2148 433292 2204
rect 433292 2148 433296 2204
rect 433232 2144 433296 2148
rect 433312 2204 433376 2208
rect 433312 2148 433316 2204
rect 433316 2148 433372 2204
rect 433372 2148 433376 2204
rect 433312 2144 433376 2148
rect 468832 2204 468896 2208
rect 468832 2148 468836 2204
rect 468836 2148 468892 2204
rect 468892 2148 468896 2204
rect 468832 2144 468896 2148
rect 468912 2204 468976 2208
rect 468912 2148 468916 2204
rect 468916 2148 468972 2204
rect 468972 2148 468976 2204
rect 468912 2144 468976 2148
rect 468992 2204 469056 2208
rect 468992 2148 468996 2204
rect 468996 2148 469052 2204
rect 469052 2148 469056 2204
rect 468992 2144 469056 2148
rect 469072 2204 469136 2208
rect 469072 2148 469076 2204
rect 469076 2148 469132 2204
rect 469132 2148 469136 2204
rect 469072 2144 469136 2148
rect 469152 2204 469216 2208
rect 469152 2148 469156 2204
rect 469156 2148 469212 2204
rect 469212 2148 469216 2204
rect 469152 2144 469216 2148
rect 469232 2204 469296 2208
rect 469232 2148 469236 2204
rect 469236 2148 469292 2204
rect 469292 2148 469296 2204
rect 469232 2144 469296 2148
rect 469312 2204 469376 2208
rect 469312 2148 469316 2204
rect 469316 2148 469372 2204
rect 469372 2148 469376 2204
rect 469312 2144 469376 2148
rect 504832 2204 504896 2208
rect 504832 2148 504836 2204
rect 504836 2148 504892 2204
rect 504892 2148 504896 2204
rect 504832 2144 504896 2148
rect 504912 2204 504976 2208
rect 504912 2148 504916 2204
rect 504916 2148 504972 2204
rect 504972 2148 504976 2204
rect 504912 2144 504976 2148
rect 504992 2204 505056 2208
rect 504992 2148 504996 2204
rect 504996 2148 505052 2204
rect 505052 2148 505056 2204
rect 504992 2144 505056 2148
rect 505072 2204 505136 2208
rect 505072 2148 505076 2204
rect 505076 2148 505132 2204
rect 505132 2148 505136 2204
rect 505072 2144 505136 2148
rect 505152 2204 505216 2208
rect 505152 2148 505156 2204
rect 505156 2148 505212 2204
rect 505212 2148 505216 2204
rect 505152 2144 505216 2148
rect 505232 2204 505296 2208
rect 505232 2148 505236 2204
rect 505236 2148 505292 2204
rect 505292 2148 505296 2204
rect 505232 2144 505296 2148
rect 505312 2204 505376 2208
rect 505312 2148 505316 2204
rect 505316 2148 505372 2204
rect 505372 2148 505376 2204
rect 505312 2144 505376 2148
rect 540832 2204 540896 2208
rect 540832 2148 540836 2204
rect 540836 2148 540892 2204
rect 540892 2148 540896 2204
rect 540832 2144 540896 2148
rect 540912 2204 540976 2208
rect 540912 2148 540916 2204
rect 540916 2148 540972 2204
rect 540972 2148 540976 2204
rect 540912 2144 540976 2148
rect 540992 2204 541056 2208
rect 540992 2148 540996 2204
rect 540996 2148 541052 2204
rect 541052 2148 541056 2204
rect 540992 2144 541056 2148
rect 541072 2204 541136 2208
rect 541072 2148 541076 2204
rect 541076 2148 541132 2204
rect 541132 2148 541136 2204
rect 541072 2144 541136 2148
rect 541152 2204 541216 2208
rect 541152 2148 541156 2204
rect 541156 2148 541212 2204
rect 541212 2148 541216 2204
rect 541152 2144 541216 2148
rect 541232 2204 541296 2208
rect 541232 2148 541236 2204
rect 541236 2148 541292 2204
rect 541292 2148 541296 2204
rect 541232 2144 541296 2148
rect 541312 2204 541376 2208
rect 541312 2148 541316 2204
rect 541316 2148 541372 2204
rect 541372 2148 541376 2204
rect 541312 2144 541376 2148
rect 576832 2204 576896 2208
rect 576832 2148 576836 2204
rect 576836 2148 576892 2204
rect 576892 2148 576896 2204
rect 576832 2144 576896 2148
rect 576912 2204 576976 2208
rect 576912 2148 576916 2204
rect 576916 2148 576972 2204
rect 576972 2148 576976 2204
rect 576912 2144 576976 2148
rect 576992 2204 577056 2208
rect 576992 2148 576996 2204
rect 576996 2148 577052 2204
rect 577052 2148 577056 2204
rect 576992 2144 577056 2148
rect 577072 2204 577136 2208
rect 577072 2148 577076 2204
rect 577076 2148 577132 2204
rect 577132 2148 577136 2204
rect 577072 2144 577136 2148
rect 577152 2204 577216 2208
rect 577152 2148 577156 2204
rect 577156 2148 577212 2204
rect 577212 2148 577216 2204
rect 577152 2144 577216 2148
rect 577232 2204 577296 2208
rect 577232 2148 577236 2204
rect 577236 2148 577292 2204
rect 577292 2148 577296 2204
rect 577232 2144 577296 2148
rect 577312 2204 577376 2208
rect 577312 2148 577316 2204
rect 577316 2148 577372 2204
rect 577372 2148 577376 2204
rect 577312 2144 577376 2148
<< metal4 >>
rect -8576 711418 -7976 711440
rect -8576 711182 -8394 711418
rect -8158 711182 -7976 711418
rect -8576 711098 -7976 711182
rect -8576 710862 -8394 711098
rect -8158 710862 -7976 711098
rect -8576 679254 -7976 710862
rect -8576 679018 -8394 679254
rect -8158 679018 -7976 679254
rect -8576 678934 -7976 679018
rect -8576 678698 -8394 678934
rect -8158 678698 -7976 678934
rect -8576 643254 -7976 678698
rect -8576 643018 -8394 643254
rect -8158 643018 -7976 643254
rect -8576 642934 -7976 643018
rect -8576 642698 -8394 642934
rect -8158 642698 -7976 642934
rect -8576 607254 -7976 642698
rect -8576 607018 -8394 607254
rect -8158 607018 -7976 607254
rect -8576 606934 -7976 607018
rect -8576 606698 -8394 606934
rect -8158 606698 -7976 606934
rect -8576 571254 -7976 606698
rect -8576 571018 -8394 571254
rect -8158 571018 -7976 571254
rect -8576 570934 -7976 571018
rect -8576 570698 -8394 570934
rect -8158 570698 -7976 570934
rect -8576 535254 -7976 570698
rect -8576 535018 -8394 535254
rect -8158 535018 -7976 535254
rect -8576 534934 -7976 535018
rect -8576 534698 -8394 534934
rect -8158 534698 -7976 534934
rect -8576 499254 -7976 534698
rect -8576 499018 -8394 499254
rect -8158 499018 -7976 499254
rect -8576 498934 -7976 499018
rect -8576 498698 -8394 498934
rect -8158 498698 -7976 498934
rect -8576 463254 -7976 498698
rect -8576 463018 -8394 463254
rect -8158 463018 -7976 463254
rect -8576 462934 -7976 463018
rect -8576 462698 -8394 462934
rect -8158 462698 -7976 462934
rect -8576 427254 -7976 462698
rect -8576 427018 -8394 427254
rect -8158 427018 -7976 427254
rect -8576 426934 -7976 427018
rect -8576 426698 -8394 426934
rect -8158 426698 -7976 426934
rect -8576 391254 -7976 426698
rect -8576 391018 -8394 391254
rect -8158 391018 -7976 391254
rect -8576 390934 -7976 391018
rect -8576 390698 -8394 390934
rect -8158 390698 -7976 390934
rect -8576 355254 -7976 390698
rect -8576 355018 -8394 355254
rect -8158 355018 -7976 355254
rect -8576 354934 -7976 355018
rect -8576 354698 -8394 354934
rect -8158 354698 -7976 354934
rect -8576 319254 -7976 354698
rect -8576 319018 -8394 319254
rect -8158 319018 -7976 319254
rect -8576 318934 -7976 319018
rect -8576 318698 -8394 318934
rect -8158 318698 -7976 318934
rect -8576 283254 -7976 318698
rect -8576 283018 -8394 283254
rect -8158 283018 -7976 283254
rect -8576 282934 -7976 283018
rect -8576 282698 -8394 282934
rect -8158 282698 -7976 282934
rect -8576 247254 -7976 282698
rect -8576 247018 -8394 247254
rect -8158 247018 -7976 247254
rect -8576 246934 -7976 247018
rect -8576 246698 -8394 246934
rect -8158 246698 -7976 246934
rect -8576 211254 -7976 246698
rect -8576 211018 -8394 211254
rect -8158 211018 -7976 211254
rect -8576 210934 -7976 211018
rect -8576 210698 -8394 210934
rect -8158 210698 -7976 210934
rect -8576 175254 -7976 210698
rect -8576 175018 -8394 175254
rect -8158 175018 -7976 175254
rect -8576 174934 -7976 175018
rect -8576 174698 -8394 174934
rect -8158 174698 -7976 174934
rect -8576 139254 -7976 174698
rect -8576 139018 -8394 139254
rect -8158 139018 -7976 139254
rect -8576 138934 -7976 139018
rect -8576 138698 -8394 138934
rect -8158 138698 -7976 138934
rect -8576 103254 -7976 138698
rect -8576 103018 -8394 103254
rect -8158 103018 -7976 103254
rect -8576 102934 -7976 103018
rect -8576 102698 -8394 102934
rect -8158 102698 -7976 102934
rect -8576 67254 -7976 102698
rect -8576 67018 -8394 67254
rect -8158 67018 -7976 67254
rect -8576 66934 -7976 67018
rect -8576 66698 -8394 66934
rect -8158 66698 -7976 66934
rect -8576 31254 -7976 66698
rect -8576 31018 -8394 31254
rect -8158 31018 -7976 31254
rect -8576 30934 -7976 31018
rect -8576 30698 -8394 30934
rect -8158 30698 -7976 30934
rect -8576 -6926 -7976 30698
rect -7636 710478 -7036 710500
rect -7636 710242 -7454 710478
rect -7218 710242 -7036 710478
rect -7636 710158 -7036 710242
rect -7636 709922 -7454 710158
rect -7218 709922 -7036 710158
rect -7636 697254 -7036 709922
rect 11604 710478 12204 711440
rect 11604 710242 11786 710478
rect 12022 710242 12204 710478
rect 11604 710158 12204 710242
rect 11604 709922 11786 710158
rect 12022 709922 12204 710158
rect -7636 697018 -7454 697254
rect -7218 697018 -7036 697254
rect -7636 696934 -7036 697018
rect -7636 696698 -7454 696934
rect -7218 696698 -7036 696934
rect -7636 661254 -7036 696698
rect -7636 661018 -7454 661254
rect -7218 661018 -7036 661254
rect -7636 660934 -7036 661018
rect -7636 660698 -7454 660934
rect -7218 660698 -7036 660934
rect -7636 625254 -7036 660698
rect -7636 625018 -7454 625254
rect -7218 625018 -7036 625254
rect -7636 624934 -7036 625018
rect -7636 624698 -7454 624934
rect -7218 624698 -7036 624934
rect -7636 589254 -7036 624698
rect -7636 589018 -7454 589254
rect -7218 589018 -7036 589254
rect -7636 588934 -7036 589018
rect -7636 588698 -7454 588934
rect -7218 588698 -7036 588934
rect -7636 553254 -7036 588698
rect -7636 553018 -7454 553254
rect -7218 553018 -7036 553254
rect -7636 552934 -7036 553018
rect -7636 552698 -7454 552934
rect -7218 552698 -7036 552934
rect -7636 517254 -7036 552698
rect -7636 517018 -7454 517254
rect -7218 517018 -7036 517254
rect -7636 516934 -7036 517018
rect -7636 516698 -7454 516934
rect -7218 516698 -7036 516934
rect -7636 481254 -7036 516698
rect -7636 481018 -7454 481254
rect -7218 481018 -7036 481254
rect -7636 480934 -7036 481018
rect -7636 480698 -7454 480934
rect -7218 480698 -7036 480934
rect -7636 445254 -7036 480698
rect -7636 445018 -7454 445254
rect -7218 445018 -7036 445254
rect -7636 444934 -7036 445018
rect -7636 444698 -7454 444934
rect -7218 444698 -7036 444934
rect -7636 409254 -7036 444698
rect -7636 409018 -7454 409254
rect -7218 409018 -7036 409254
rect -7636 408934 -7036 409018
rect -7636 408698 -7454 408934
rect -7218 408698 -7036 408934
rect -7636 373254 -7036 408698
rect -7636 373018 -7454 373254
rect -7218 373018 -7036 373254
rect -7636 372934 -7036 373018
rect -7636 372698 -7454 372934
rect -7218 372698 -7036 372934
rect -7636 337254 -7036 372698
rect -7636 337018 -7454 337254
rect -7218 337018 -7036 337254
rect -7636 336934 -7036 337018
rect -7636 336698 -7454 336934
rect -7218 336698 -7036 336934
rect -7636 301254 -7036 336698
rect -7636 301018 -7454 301254
rect -7218 301018 -7036 301254
rect -7636 300934 -7036 301018
rect -7636 300698 -7454 300934
rect -7218 300698 -7036 300934
rect -7636 265254 -7036 300698
rect -7636 265018 -7454 265254
rect -7218 265018 -7036 265254
rect -7636 264934 -7036 265018
rect -7636 264698 -7454 264934
rect -7218 264698 -7036 264934
rect -7636 229254 -7036 264698
rect -7636 229018 -7454 229254
rect -7218 229018 -7036 229254
rect -7636 228934 -7036 229018
rect -7636 228698 -7454 228934
rect -7218 228698 -7036 228934
rect -7636 193254 -7036 228698
rect -7636 193018 -7454 193254
rect -7218 193018 -7036 193254
rect -7636 192934 -7036 193018
rect -7636 192698 -7454 192934
rect -7218 192698 -7036 192934
rect -7636 157254 -7036 192698
rect -7636 157018 -7454 157254
rect -7218 157018 -7036 157254
rect -7636 156934 -7036 157018
rect -7636 156698 -7454 156934
rect -7218 156698 -7036 156934
rect -7636 121254 -7036 156698
rect -7636 121018 -7454 121254
rect -7218 121018 -7036 121254
rect -7636 120934 -7036 121018
rect -7636 120698 -7454 120934
rect -7218 120698 -7036 120934
rect -7636 85254 -7036 120698
rect -7636 85018 -7454 85254
rect -7218 85018 -7036 85254
rect -7636 84934 -7036 85018
rect -7636 84698 -7454 84934
rect -7218 84698 -7036 84934
rect -7636 49254 -7036 84698
rect -7636 49018 -7454 49254
rect -7218 49018 -7036 49254
rect -7636 48934 -7036 49018
rect -7636 48698 -7454 48934
rect -7218 48698 -7036 48934
rect -7636 13254 -7036 48698
rect -7636 13018 -7454 13254
rect -7218 13018 -7036 13254
rect -7636 12934 -7036 13018
rect -7636 12698 -7454 12934
rect -7218 12698 -7036 12934
rect -7636 -5986 -7036 12698
rect -6696 709538 -6096 709560
rect -6696 709302 -6514 709538
rect -6278 709302 -6096 709538
rect -6696 709218 -6096 709302
rect -6696 708982 -6514 709218
rect -6278 708982 -6096 709218
rect -6696 675654 -6096 708982
rect -6696 675418 -6514 675654
rect -6278 675418 -6096 675654
rect -6696 675334 -6096 675418
rect -6696 675098 -6514 675334
rect -6278 675098 -6096 675334
rect -6696 639654 -6096 675098
rect -6696 639418 -6514 639654
rect -6278 639418 -6096 639654
rect -6696 639334 -6096 639418
rect -6696 639098 -6514 639334
rect -6278 639098 -6096 639334
rect -6696 603654 -6096 639098
rect -6696 603418 -6514 603654
rect -6278 603418 -6096 603654
rect -6696 603334 -6096 603418
rect -6696 603098 -6514 603334
rect -6278 603098 -6096 603334
rect -6696 567654 -6096 603098
rect -6696 567418 -6514 567654
rect -6278 567418 -6096 567654
rect -6696 567334 -6096 567418
rect -6696 567098 -6514 567334
rect -6278 567098 -6096 567334
rect -6696 531654 -6096 567098
rect -6696 531418 -6514 531654
rect -6278 531418 -6096 531654
rect -6696 531334 -6096 531418
rect -6696 531098 -6514 531334
rect -6278 531098 -6096 531334
rect -6696 495654 -6096 531098
rect -6696 495418 -6514 495654
rect -6278 495418 -6096 495654
rect -6696 495334 -6096 495418
rect -6696 495098 -6514 495334
rect -6278 495098 -6096 495334
rect -6696 459654 -6096 495098
rect -6696 459418 -6514 459654
rect -6278 459418 -6096 459654
rect -6696 459334 -6096 459418
rect -6696 459098 -6514 459334
rect -6278 459098 -6096 459334
rect -6696 423654 -6096 459098
rect -6696 423418 -6514 423654
rect -6278 423418 -6096 423654
rect -6696 423334 -6096 423418
rect -6696 423098 -6514 423334
rect -6278 423098 -6096 423334
rect -6696 387654 -6096 423098
rect -6696 387418 -6514 387654
rect -6278 387418 -6096 387654
rect -6696 387334 -6096 387418
rect -6696 387098 -6514 387334
rect -6278 387098 -6096 387334
rect -6696 351654 -6096 387098
rect -6696 351418 -6514 351654
rect -6278 351418 -6096 351654
rect -6696 351334 -6096 351418
rect -6696 351098 -6514 351334
rect -6278 351098 -6096 351334
rect -6696 315654 -6096 351098
rect -6696 315418 -6514 315654
rect -6278 315418 -6096 315654
rect -6696 315334 -6096 315418
rect -6696 315098 -6514 315334
rect -6278 315098 -6096 315334
rect -6696 279654 -6096 315098
rect -6696 279418 -6514 279654
rect -6278 279418 -6096 279654
rect -6696 279334 -6096 279418
rect -6696 279098 -6514 279334
rect -6278 279098 -6096 279334
rect -6696 243654 -6096 279098
rect -6696 243418 -6514 243654
rect -6278 243418 -6096 243654
rect -6696 243334 -6096 243418
rect -6696 243098 -6514 243334
rect -6278 243098 -6096 243334
rect -6696 207654 -6096 243098
rect -6696 207418 -6514 207654
rect -6278 207418 -6096 207654
rect -6696 207334 -6096 207418
rect -6696 207098 -6514 207334
rect -6278 207098 -6096 207334
rect -6696 171654 -6096 207098
rect -6696 171418 -6514 171654
rect -6278 171418 -6096 171654
rect -6696 171334 -6096 171418
rect -6696 171098 -6514 171334
rect -6278 171098 -6096 171334
rect -6696 135654 -6096 171098
rect -6696 135418 -6514 135654
rect -6278 135418 -6096 135654
rect -6696 135334 -6096 135418
rect -6696 135098 -6514 135334
rect -6278 135098 -6096 135334
rect -6696 99654 -6096 135098
rect -6696 99418 -6514 99654
rect -6278 99418 -6096 99654
rect -6696 99334 -6096 99418
rect -6696 99098 -6514 99334
rect -6278 99098 -6096 99334
rect -6696 63654 -6096 99098
rect -6696 63418 -6514 63654
rect -6278 63418 -6096 63654
rect -6696 63334 -6096 63418
rect -6696 63098 -6514 63334
rect -6278 63098 -6096 63334
rect -6696 27654 -6096 63098
rect -6696 27418 -6514 27654
rect -6278 27418 -6096 27654
rect -6696 27334 -6096 27418
rect -6696 27098 -6514 27334
rect -6278 27098 -6096 27334
rect -6696 -5046 -6096 27098
rect -5756 708598 -5156 708620
rect -5756 708362 -5574 708598
rect -5338 708362 -5156 708598
rect -5756 708278 -5156 708362
rect -5756 708042 -5574 708278
rect -5338 708042 -5156 708278
rect -5756 693654 -5156 708042
rect 8004 708598 8604 709560
rect 8004 708362 8186 708598
rect 8422 708362 8604 708598
rect 8004 708278 8604 708362
rect 8004 708042 8186 708278
rect 8422 708042 8604 708278
rect -5756 693418 -5574 693654
rect -5338 693418 -5156 693654
rect -5756 693334 -5156 693418
rect -5756 693098 -5574 693334
rect -5338 693098 -5156 693334
rect -5756 657654 -5156 693098
rect -5756 657418 -5574 657654
rect -5338 657418 -5156 657654
rect -5756 657334 -5156 657418
rect -5756 657098 -5574 657334
rect -5338 657098 -5156 657334
rect -5756 621654 -5156 657098
rect -5756 621418 -5574 621654
rect -5338 621418 -5156 621654
rect -5756 621334 -5156 621418
rect -5756 621098 -5574 621334
rect -5338 621098 -5156 621334
rect -5756 585654 -5156 621098
rect -5756 585418 -5574 585654
rect -5338 585418 -5156 585654
rect -5756 585334 -5156 585418
rect -5756 585098 -5574 585334
rect -5338 585098 -5156 585334
rect -5756 549654 -5156 585098
rect -5756 549418 -5574 549654
rect -5338 549418 -5156 549654
rect -5756 549334 -5156 549418
rect -5756 549098 -5574 549334
rect -5338 549098 -5156 549334
rect -5756 513654 -5156 549098
rect -5756 513418 -5574 513654
rect -5338 513418 -5156 513654
rect -5756 513334 -5156 513418
rect -5756 513098 -5574 513334
rect -5338 513098 -5156 513334
rect -5756 477654 -5156 513098
rect -5756 477418 -5574 477654
rect -5338 477418 -5156 477654
rect -5756 477334 -5156 477418
rect -5756 477098 -5574 477334
rect -5338 477098 -5156 477334
rect -5756 441654 -5156 477098
rect -5756 441418 -5574 441654
rect -5338 441418 -5156 441654
rect -5756 441334 -5156 441418
rect -5756 441098 -5574 441334
rect -5338 441098 -5156 441334
rect -5756 405654 -5156 441098
rect -5756 405418 -5574 405654
rect -5338 405418 -5156 405654
rect -5756 405334 -5156 405418
rect -5756 405098 -5574 405334
rect -5338 405098 -5156 405334
rect -5756 369654 -5156 405098
rect -5756 369418 -5574 369654
rect -5338 369418 -5156 369654
rect -5756 369334 -5156 369418
rect -5756 369098 -5574 369334
rect -5338 369098 -5156 369334
rect -5756 333654 -5156 369098
rect -5756 333418 -5574 333654
rect -5338 333418 -5156 333654
rect -5756 333334 -5156 333418
rect -5756 333098 -5574 333334
rect -5338 333098 -5156 333334
rect -5756 297654 -5156 333098
rect -5756 297418 -5574 297654
rect -5338 297418 -5156 297654
rect -5756 297334 -5156 297418
rect -5756 297098 -5574 297334
rect -5338 297098 -5156 297334
rect -5756 261654 -5156 297098
rect -5756 261418 -5574 261654
rect -5338 261418 -5156 261654
rect -5756 261334 -5156 261418
rect -5756 261098 -5574 261334
rect -5338 261098 -5156 261334
rect -5756 225654 -5156 261098
rect -5756 225418 -5574 225654
rect -5338 225418 -5156 225654
rect -5756 225334 -5156 225418
rect -5756 225098 -5574 225334
rect -5338 225098 -5156 225334
rect -5756 189654 -5156 225098
rect -5756 189418 -5574 189654
rect -5338 189418 -5156 189654
rect -5756 189334 -5156 189418
rect -5756 189098 -5574 189334
rect -5338 189098 -5156 189334
rect -5756 153654 -5156 189098
rect -5756 153418 -5574 153654
rect -5338 153418 -5156 153654
rect -5756 153334 -5156 153418
rect -5756 153098 -5574 153334
rect -5338 153098 -5156 153334
rect -5756 117654 -5156 153098
rect -5756 117418 -5574 117654
rect -5338 117418 -5156 117654
rect -5756 117334 -5156 117418
rect -5756 117098 -5574 117334
rect -5338 117098 -5156 117334
rect -5756 81654 -5156 117098
rect -5756 81418 -5574 81654
rect -5338 81418 -5156 81654
rect -5756 81334 -5156 81418
rect -5756 81098 -5574 81334
rect -5338 81098 -5156 81334
rect -5756 45654 -5156 81098
rect -5756 45418 -5574 45654
rect -5338 45418 -5156 45654
rect -5756 45334 -5156 45418
rect -5756 45098 -5574 45334
rect -5338 45098 -5156 45334
rect -5756 9654 -5156 45098
rect -5756 9418 -5574 9654
rect -5338 9418 -5156 9654
rect -5756 9334 -5156 9418
rect -5756 9098 -5574 9334
rect -5338 9098 -5156 9334
rect -5756 -4106 -5156 9098
rect -4816 707658 -4216 707680
rect -4816 707422 -4634 707658
rect -4398 707422 -4216 707658
rect -4816 707338 -4216 707422
rect -4816 707102 -4634 707338
rect -4398 707102 -4216 707338
rect -4816 672054 -4216 707102
rect -4816 671818 -4634 672054
rect -4398 671818 -4216 672054
rect -4816 671734 -4216 671818
rect -4816 671498 -4634 671734
rect -4398 671498 -4216 671734
rect -4816 636054 -4216 671498
rect -4816 635818 -4634 636054
rect -4398 635818 -4216 636054
rect -4816 635734 -4216 635818
rect -4816 635498 -4634 635734
rect -4398 635498 -4216 635734
rect -4816 600054 -4216 635498
rect -4816 599818 -4634 600054
rect -4398 599818 -4216 600054
rect -4816 599734 -4216 599818
rect -4816 599498 -4634 599734
rect -4398 599498 -4216 599734
rect -4816 564054 -4216 599498
rect -4816 563818 -4634 564054
rect -4398 563818 -4216 564054
rect -4816 563734 -4216 563818
rect -4816 563498 -4634 563734
rect -4398 563498 -4216 563734
rect -4816 528054 -4216 563498
rect -4816 527818 -4634 528054
rect -4398 527818 -4216 528054
rect -4816 527734 -4216 527818
rect -4816 527498 -4634 527734
rect -4398 527498 -4216 527734
rect -4816 492054 -4216 527498
rect -4816 491818 -4634 492054
rect -4398 491818 -4216 492054
rect -4816 491734 -4216 491818
rect -4816 491498 -4634 491734
rect -4398 491498 -4216 491734
rect -4816 456054 -4216 491498
rect -4816 455818 -4634 456054
rect -4398 455818 -4216 456054
rect -4816 455734 -4216 455818
rect -4816 455498 -4634 455734
rect -4398 455498 -4216 455734
rect -4816 420054 -4216 455498
rect -4816 419818 -4634 420054
rect -4398 419818 -4216 420054
rect -4816 419734 -4216 419818
rect -4816 419498 -4634 419734
rect -4398 419498 -4216 419734
rect -4816 384054 -4216 419498
rect -4816 383818 -4634 384054
rect -4398 383818 -4216 384054
rect -4816 383734 -4216 383818
rect -4816 383498 -4634 383734
rect -4398 383498 -4216 383734
rect -4816 348054 -4216 383498
rect -4816 347818 -4634 348054
rect -4398 347818 -4216 348054
rect -4816 347734 -4216 347818
rect -4816 347498 -4634 347734
rect -4398 347498 -4216 347734
rect -4816 312054 -4216 347498
rect -4816 311818 -4634 312054
rect -4398 311818 -4216 312054
rect -4816 311734 -4216 311818
rect -4816 311498 -4634 311734
rect -4398 311498 -4216 311734
rect -4816 276054 -4216 311498
rect -4816 275818 -4634 276054
rect -4398 275818 -4216 276054
rect -4816 275734 -4216 275818
rect -4816 275498 -4634 275734
rect -4398 275498 -4216 275734
rect -4816 240054 -4216 275498
rect -4816 239818 -4634 240054
rect -4398 239818 -4216 240054
rect -4816 239734 -4216 239818
rect -4816 239498 -4634 239734
rect -4398 239498 -4216 239734
rect -4816 204054 -4216 239498
rect -4816 203818 -4634 204054
rect -4398 203818 -4216 204054
rect -4816 203734 -4216 203818
rect -4816 203498 -4634 203734
rect -4398 203498 -4216 203734
rect -4816 168054 -4216 203498
rect -4816 167818 -4634 168054
rect -4398 167818 -4216 168054
rect -4816 167734 -4216 167818
rect -4816 167498 -4634 167734
rect -4398 167498 -4216 167734
rect -4816 132054 -4216 167498
rect -4816 131818 -4634 132054
rect -4398 131818 -4216 132054
rect -4816 131734 -4216 131818
rect -4816 131498 -4634 131734
rect -4398 131498 -4216 131734
rect -4816 96054 -4216 131498
rect -4816 95818 -4634 96054
rect -4398 95818 -4216 96054
rect -4816 95734 -4216 95818
rect -4816 95498 -4634 95734
rect -4398 95498 -4216 95734
rect -4816 60054 -4216 95498
rect -4816 59818 -4634 60054
rect -4398 59818 -4216 60054
rect -4816 59734 -4216 59818
rect -4816 59498 -4634 59734
rect -4398 59498 -4216 59734
rect -4816 24054 -4216 59498
rect -4816 23818 -4634 24054
rect -4398 23818 -4216 24054
rect -4816 23734 -4216 23818
rect -4816 23498 -4634 23734
rect -4398 23498 -4216 23734
rect -4816 -3166 -4216 23498
rect -3876 706718 -3276 706740
rect -3876 706482 -3694 706718
rect -3458 706482 -3276 706718
rect -3876 706398 -3276 706482
rect -3876 706162 -3694 706398
rect -3458 706162 -3276 706398
rect -3876 690054 -3276 706162
rect 4404 706718 5004 707680
rect 4404 706482 4586 706718
rect 4822 706482 5004 706718
rect 4404 706398 5004 706482
rect 4404 706162 4586 706398
rect 4822 706162 5004 706398
rect -3876 689818 -3694 690054
rect -3458 689818 -3276 690054
rect -3876 689734 -3276 689818
rect -3876 689498 -3694 689734
rect -3458 689498 -3276 689734
rect -3876 654054 -3276 689498
rect -3876 653818 -3694 654054
rect -3458 653818 -3276 654054
rect -3876 653734 -3276 653818
rect -3876 653498 -3694 653734
rect -3458 653498 -3276 653734
rect -3876 618054 -3276 653498
rect -3876 617818 -3694 618054
rect -3458 617818 -3276 618054
rect -3876 617734 -3276 617818
rect -3876 617498 -3694 617734
rect -3458 617498 -3276 617734
rect -3876 582054 -3276 617498
rect -3876 581818 -3694 582054
rect -3458 581818 -3276 582054
rect -3876 581734 -3276 581818
rect -3876 581498 -3694 581734
rect -3458 581498 -3276 581734
rect -3876 546054 -3276 581498
rect -3876 545818 -3694 546054
rect -3458 545818 -3276 546054
rect -3876 545734 -3276 545818
rect -3876 545498 -3694 545734
rect -3458 545498 -3276 545734
rect -3876 510054 -3276 545498
rect -3876 509818 -3694 510054
rect -3458 509818 -3276 510054
rect -3876 509734 -3276 509818
rect -3876 509498 -3694 509734
rect -3458 509498 -3276 509734
rect -3876 474054 -3276 509498
rect -3876 473818 -3694 474054
rect -3458 473818 -3276 474054
rect -3876 473734 -3276 473818
rect -3876 473498 -3694 473734
rect -3458 473498 -3276 473734
rect -3876 438054 -3276 473498
rect -3876 437818 -3694 438054
rect -3458 437818 -3276 438054
rect -3876 437734 -3276 437818
rect -3876 437498 -3694 437734
rect -3458 437498 -3276 437734
rect -3876 402054 -3276 437498
rect -3876 401818 -3694 402054
rect -3458 401818 -3276 402054
rect -3876 401734 -3276 401818
rect -3876 401498 -3694 401734
rect -3458 401498 -3276 401734
rect -3876 366054 -3276 401498
rect -3876 365818 -3694 366054
rect -3458 365818 -3276 366054
rect -3876 365734 -3276 365818
rect -3876 365498 -3694 365734
rect -3458 365498 -3276 365734
rect -3876 330054 -3276 365498
rect -3876 329818 -3694 330054
rect -3458 329818 -3276 330054
rect -3876 329734 -3276 329818
rect -3876 329498 -3694 329734
rect -3458 329498 -3276 329734
rect -3876 294054 -3276 329498
rect -3876 293818 -3694 294054
rect -3458 293818 -3276 294054
rect -3876 293734 -3276 293818
rect -3876 293498 -3694 293734
rect -3458 293498 -3276 293734
rect -3876 258054 -3276 293498
rect -3876 257818 -3694 258054
rect -3458 257818 -3276 258054
rect -3876 257734 -3276 257818
rect -3876 257498 -3694 257734
rect -3458 257498 -3276 257734
rect -3876 222054 -3276 257498
rect -3876 221818 -3694 222054
rect -3458 221818 -3276 222054
rect -3876 221734 -3276 221818
rect -3876 221498 -3694 221734
rect -3458 221498 -3276 221734
rect -3876 186054 -3276 221498
rect -3876 185818 -3694 186054
rect -3458 185818 -3276 186054
rect -3876 185734 -3276 185818
rect -3876 185498 -3694 185734
rect -3458 185498 -3276 185734
rect -3876 150054 -3276 185498
rect -3876 149818 -3694 150054
rect -3458 149818 -3276 150054
rect -3876 149734 -3276 149818
rect -3876 149498 -3694 149734
rect -3458 149498 -3276 149734
rect -3876 114054 -3276 149498
rect -3876 113818 -3694 114054
rect -3458 113818 -3276 114054
rect -3876 113734 -3276 113818
rect -3876 113498 -3694 113734
rect -3458 113498 -3276 113734
rect -3876 78054 -3276 113498
rect -3876 77818 -3694 78054
rect -3458 77818 -3276 78054
rect -3876 77734 -3276 77818
rect -3876 77498 -3694 77734
rect -3458 77498 -3276 77734
rect -3876 42054 -3276 77498
rect -3876 41818 -3694 42054
rect -3458 41818 -3276 42054
rect -3876 41734 -3276 41818
rect -3876 41498 -3694 41734
rect -3458 41498 -3276 41734
rect -3876 6054 -3276 41498
rect -3876 5818 -3694 6054
rect -3458 5818 -3276 6054
rect -3876 5734 -3276 5818
rect -3876 5498 -3694 5734
rect -3458 5498 -3276 5734
rect -3876 -2226 -3276 5498
rect -2936 705778 -2336 705800
rect -2936 705542 -2754 705778
rect -2518 705542 -2336 705778
rect -2936 705458 -2336 705542
rect -2936 705222 -2754 705458
rect -2518 705222 -2336 705458
rect -2936 668406 -2336 705222
rect -2936 668170 -2754 668406
rect -2518 668170 -2336 668406
rect -2936 668086 -2336 668170
rect -2936 667850 -2754 668086
rect -2518 667850 -2336 668086
rect -2936 632406 -2336 667850
rect -2936 632170 -2754 632406
rect -2518 632170 -2336 632406
rect -2936 632086 -2336 632170
rect -2936 631850 -2754 632086
rect -2518 631850 -2336 632086
rect -2936 596406 -2336 631850
rect -2936 596170 -2754 596406
rect -2518 596170 -2336 596406
rect -2936 596086 -2336 596170
rect -2936 595850 -2754 596086
rect -2518 595850 -2336 596086
rect -2936 560406 -2336 595850
rect -2936 560170 -2754 560406
rect -2518 560170 -2336 560406
rect -2936 560086 -2336 560170
rect -2936 559850 -2754 560086
rect -2518 559850 -2336 560086
rect -2936 524406 -2336 559850
rect -2936 524170 -2754 524406
rect -2518 524170 -2336 524406
rect -2936 524086 -2336 524170
rect -2936 523850 -2754 524086
rect -2518 523850 -2336 524086
rect -2936 488406 -2336 523850
rect -2936 488170 -2754 488406
rect -2518 488170 -2336 488406
rect -2936 488086 -2336 488170
rect -2936 487850 -2754 488086
rect -2518 487850 -2336 488086
rect -2936 452406 -2336 487850
rect -2936 452170 -2754 452406
rect -2518 452170 -2336 452406
rect -2936 452086 -2336 452170
rect -2936 451850 -2754 452086
rect -2518 451850 -2336 452086
rect -2936 416406 -2336 451850
rect -2936 416170 -2754 416406
rect -2518 416170 -2336 416406
rect -2936 416086 -2336 416170
rect -2936 415850 -2754 416086
rect -2518 415850 -2336 416086
rect -2936 380406 -2336 415850
rect -2936 380170 -2754 380406
rect -2518 380170 -2336 380406
rect -2936 380086 -2336 380170
rect -2936 379850 -2754 380086
rect -2518 379850 -2336 380086
rect -2936 344406 -2336 379850
rect -2936 344170 -2754 344406
rect -2518 344170 -2336 344406
rect -2936 344086 -2336 344170
rect -2936 343850 -2754 344086
rect -2518 343850 -2336 344086
rect -2936 308406 -2336 343850
rect -2936 308170 -2754 308406
rect -2518 308170 -2336 308406
rect -2936 308086 -2336 308170
rect -2936 307850 -2754 308086
rect -2518 307850 -2336 308086
rect -2936 272406 -2336 307850
rect -2936 272170 -2754 272406
rect -2518 272170 -2336 272406
rect -2936 272086 -2336 272170
rect -2936 271850 -2754 272086
rect -2518 271850 -2336 272086
rect -2936 236406 -2336 271850
rect -2936 236170 -2754 236406
rect -2518 236170 -2336 236406
rect -2936 236086 -2336 236170
rect -2936 235850 -2754 236086
rect -2518 235850 -2336 236086
rect -2936 200406 -2336 235850
rect -2936 200170 -2754 200406
rect -2518 200170 -2336 200406
rect -2936 200086 -2336 200170
rect -2936 199850 -2754 200086
rect -2518 199850 -2336 200086
rect -2936 164406 -2336 199850
rect -2936 164170 -2754 164406
rect -2518 164170 -2336 164406
rect -2936 164086 -2336 164170
rect -2936 163850 -2754 164086
rect -2518 163850 -2336 164086
rect -2936 128406 -2336 163850
rect -2936 128170 -2754 128406
rect -2518 128170 -2336 128406
rect -2936 128086 -2336 128170
rect -2936 127850 -2754 128086
rect -2518 127850 -2336 128086
rect -2936 92406 -2336 127850
rect -2936 92170 -2754 92406
rect -2518 92170 -2336 92406
rect -2936 92086 -2336 92170
rect -2936 91850 -2754 92086
rect -2518 91850 -2336 92086
rect -2936 56406 -2336 91850
rect -2936 56170 -2754 56406
rect -2518 56170 -2336 56406
rect -2936 56086 -2336 56170
rect -2936 55850 -2754 56086
rect -2518 55850 -2336 56086
rect -2936 20406 -2336 55850
rect -2936 20170 -2754 20406
rect -2518 20170 -2336 20406
rect -2936 20086 -2336 20170
rect -2936 19850 -2754 20086
rect -2518 19850 -2336 20086
rect -2936 -1286 -2336 19850
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686406 -1396 704282
rect -1996 686170 -1814 686406
rect -1578 686170 -1396 686406
rect -1996 686086 -1396 686170
rect -1996 685850 -1814 686086
rect -1578 685850 -1396 686086
rect -1996 650406 -1396 685850
rect -1996 650170 -1814 650406
rect -1578 650170 -1396 650406
rect -1996 650086 -1396 650170
rect -1996 649850 -1814 650086
rect -1578 649850 -1396 650086
rect -1996 614406 -1396 649850
rect -1996 614170 -1814 614406
rect -1578 614170 -1396 614406
rect -1996 614086 -1396 614170
rect -1996 613850 -1814 614086
rect -1578 613850 -1396 614086
rect -1996 578406 -1396 613850
rect -1996 578170 -1814 578406
rect -1578 578170 -1396 578406
rect -1996 578086 -1396 578170
rect -1996 577850 -1814 578086
rect -1578 577850 -1396 578086
rect -1996 542406 -1396 577850
rect -1996 542170 -1814 542406
rect -1578 542170 -1396 542406
rect -1996 542086 -1396 542170
rect -1996 541850 -1814 542086
rect -1578 541850 -1396 542086
rect -1996 506406 -1396 541850
rect -1996 506170 -1814 506406
rect -1578 506170 -1396 506406
rect -1996 506086 -1396 506170
rect -1996 505850 -1814 506086
rect -1578 505850 -1396 506086
rect -1996 470406 -1396 505850
rect -1996 470170 -1814 470406
rect -1578 470170 -1396 470406
rect -1996 470086 -1396 470170
rect -1996 469850 -1814 470086
rect -1578 469850 -1396 470086
rect -1996 434406 -1396 469850
rect -1996 434170 -1814 434406
rect -1578 434170 -1396 434406
rect -1996 434086 -1396 434170
rect -1996 433850 -1814 434086
rect -1578 433850 -1396 434086
rect -1996 398406 -1396 433850
rect -1996 398170 -1814 398406
rect -1578 398170 -1396 398406
rect -1996 398086 -1396 398170
rect -1996 397850 -1814 398086
rect -1578 397850 -1396 398086
rect -1996 362406 -1396 397850
rect -1996 362170 -1814 362406
rect -1578 362170 -1396 362406
rect -1996 362086 -1396 362170
rect -1996 361850 -1814 362086
rect -1578 361850 -1396 362086
rect -1996 326406 -1396 361850
rect -1996 326170 -1814 326406
rect -1578 326170 -1396 326406
rect -1996 326086 -1396 326170
rect -1996 325850 -1814 326086
rect -1578 325850 -1396 326086
rect -1996 290406 -1396 325850
rect -1996 290170 -1814 290406
rect -1578 290170 -1396 290406
rect -1996 290086 -1396 290170
rect -1996 289850 -1814 290086
rect -1578 289850 -1396 290086
rect -1996 254406 -1396 289850
rect -1996 254170 -1814 254406
rect -1578 254170 -1396 254406
rect -1996 254086 -1396 254170
rect -1996 253850 -1814 254086
rect -1578 253850 -1396 254086
rect -1996 218406 -1396 253850
rect -1996 218170 -1814 218406
rect -1578 218170 -1396 218406
rect -1996 218086 -1396 218170
rect -1996 217850 -1814 218086
rect -1578 217850 -1396 218086
rect -1996 182406 -1396 217850
rect -1996 182170 -1814 182406
rect -1578 182170 -1396 182406
rect -1996 182086 -1396 182170
rect -1996 181850 -1814 182086
rect -1578 181850 -1396 182086
rect -1996 146406 -1396 181850
rect -1996 146170 -1814 146406
rect -1578 146170 -1396 146406
rect -1996 146086 -1396 146170
rect -1996 145850 -1814 146086
rect -1578 145850 -1396 146086
rect -1996 110406 -1396 145850
rect -1996 110170 -1814 110406
rect -1578 110170 -1396 110406
rect -1996 110086 -1396 110170
rect -1996 109850 -1814 110086
rect -1578 109850 -1396 110086
rect -1996 74406 -1396 109850
rect -1996 74170 -1814 74406
rect -1578 74170 -1396 74406
rect -1996 74086 -1396 74170
rect -1996 73850 -1814 74086
rect -1578 73850 -1396 74086
rect -1996 38406 -1396 73850
rect -1996 38170 -1814 38406
rect -1578 38170 -1396 38406
rect -1996 38086 -1396 38170
rect -1996 37850 -1814 38086
rect -1578 37850 -1396 38086
rect -1996 2406 -1396 37850
rect -1996 2170 -1814 2406
rect -1578 2170 -1396 2406
rect -1996 2086 -1396 2170
rect -1996 1850 -1814 2086
rect -1578 1850 -1396 2086
rect -1996 -346 -1396 1850
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705800
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686406 1404 704282
rect 804 686170 986 686406
rect 1222 686170 1404 686406
rect 804 686086 1404 686170
rect 804 685850 986 686086
rect 1222 685850 1404 686086
rect 804 650406 1404 685850
rect 804 650170 986 650406
rect 1222 650170 1404 650406
rect 804 650086 1404 650170
rect 804 649850 986 650086
rect 1222 649850 1404 650086
rect 804 614406 1404 649850
rect 804 614170 986 614406
rect 1222 614170 1404 614406
rect 804 614086 1404 614170
rect 804 613850 986 614086
rect 1222 613850 1404 614086
rect 804 578406 1404 613850
rect 804 578170 986 578406
rect 1222 578170 1404 578406
rect 804 578086 1404 578170
rect 804 577850 986 578086
rect 1222 577850 1404 578086
rect 804 542406 1404 577850
rect 804 542170 986 542406
rect 1222 542170 1404 542406
rect 804 542086 1404 542170
rect 804 541850 986 542086
rect 1222 541850 1404 542086
rect 804 506406 1404 541850
rect 804 506170 986 506406
rect 1222 506170 1404 506406
rect 804 506086 1404 506170
rect 804 505850 986 506086
rect 1222 505850 1404 506086
rect 804 470406 1404 505850
rect 804 470170 986 470406
rect 1222 470170 1404 470406
rect 804 470086 1404 470170
rect 804 469850 986 470086
rect 1222 469850 1404 470086
rect 804 434406 1404 469850
rect 804 434170 986 434406
rect 1222 434170 1404 434406
rect 804 434086 1404 434170
rect 804 433850 986 434086
rect 1222 433850 1404 434086
rect 804 398406 1404 433850
rect 804 398170 986 398406
rect 1222 398170 1404 398406
rect 804 398086 1404 398170
rect 804 397850 986 398086
rect 1222 397850 1404 398086
rect 804 362406 1404 397850
rect 804 362170 986 362406
rect 1222 362170 1404 362406
rect 804 362086 1404 362170
rect 804 361850 986 362086
rect 1222 361850 1404 362086
rect 804 326406 1404 361850
rect 804 326170 986 326406
rect 1222 326170 1404 326406
rect 804 326086 1404 326170
rect 804 325850 986 326086
rect 1222 325850 1404 326086
rect 804 290406 1404 325850
rect 804 290170 986 290406
rect 1222 290170 1404 290406
rect 804 290086 1404 290170
rect 804 289850 986 290086
rect 1222 289850 1404 290086
rect 804 254406 1404 289850
rect 804 254170 986 254406
rect 1222 254170 1404 254406
rect 804 254086 1404 254170
rect 804 253850 986 254086
rect 1222 253850 1404 254086
rect 804 218406 1404 253850
rect 804 218170 986 218406
rect 1222 218170 1404 218406
rect 804 218086 1404 218170
rect 804 217850 986 218086
rect 1222 217850 1404 218086
rect 804 182406 1404 217850
rect 804 182170 986 182406
rect 1222 182170 1404 182406
rect 804 182086 1404 182170
rect 804 181850 986 182086
rect 1222 181850 1404 182086
rect 804 146406 1404 181850
rect 804 146170 986 146406
rect 1222 146170 1404 146406
rect 804 146086 1404 146170
rect 804 145850 986 146086
rect 1222 145850 1404 146086
rect 804 110406 1404 145850
rect 804 110170 986 110406
rect 1222 110170 1404 110406
rect 804 110086 1404 110170
rect 804 109850 986 110086
rect 1222 109850 1404 110086
rect 804 74406 1404 109850
rect 804 74170 986 74406
rect 1222 74170 1404 74406
rect 804 74086 1404 74170
rect 804 73850 986 74086
rect 1222 73850 1404 74086
rect 804 38406 1404 73850
rect 804 38170 986 38406
rect 1222 38170 1404 38406
rect 804 38086 1404 38170
rect 804 37850 986 38086
rect 1222 37850 1404 38086
rect 804 2406 1404 37850
rect 804 2170 986 2406
rect 1222 2170 1404 2406
rect 804 2086 1404 2170
rect 804 1850 986 2086
rect 1222 1850 1404 2086
rect 804 -346 1404 1850
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2936 -1522 -2754 -1286
rect -2518 -1522 -2336 -1286
rect -2936 -1606 -2336 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 -2336 -1606
rect -2936 -1864 -2336 -1842
rect 804 -1864 1404 -902
rect 4404 690054 5004 706162
rect 8004 698000 8604 708042
rect 11604 698000 12204 709922
rect 29604 711418 30204 711440
rect 29604 711182 29786 711418
rect 30022 711182 30204 711418
rect 29604 711098 30204 711182
rect 29604 710862 29786 711098
rect 30022 710862 30204 711098
rect 26004 709538 26604 709560
rect 26004 709302 26186 709538
rect 26422 709302 26604 709538
rect 26004 709218 26604 709302
rect 26004 708982 26186 709218
rect 26422 708982 26604 709218
rect 22404 707658 23004 707680
rect 22404 707422 22586 707658
rect 22822 707422 23004 707658
rect 22404 707338 23004 707422
rect 22404 707102 22586 707338
rect 22822 707102 23004 707338
rect 18804 705778 19404 705800
rect 18804 705542 18986 705778
rect 19222 705542 19404 705778
rect 18804 705458 19404 705542
rect 18804 705222 18986 705458
rect 19222 705222 19404 705458
rect 18804 701248 19404 705222
rect 18804 701184 18832 701248
rect 18896 701184 18912 701248
rect 18976 701184 18992 701248
rect 19056 701184 19072 701248
rect 19136 701184 19152 701248
rect 19216 701184 19232 701248
rect 19296 701184 19312 701248
rect 19376 701184 19404 701248
rect 18804 700160 19404 701184
rect 18804 700096 18832 700160
rect 18896 700096 18912 700160
rect 18976 700096 18992 700160
rect 19056 700096 19072 700160
rect 19136 700096 19152 700160
rect 19216 700096 19232 700160
rect 19296 700096 19312 700160
rect 19376 700096 19404 700160
rect 18804 699072 19404 700096
rect 18804 699008 18832 699072
rect 18896 699008 18912 699072
rect 18976 699008 18992 699072
rect 19056 699008 19072 699072
rect 19136 699008 19152 699072
rect 19216 699008 19232 699072
rect 19296 699008 19312 699072
rect 19376 699008 19404 699072
rect 18804 697952 19404 699008
rect 22404 698000 23004 707102
rect 26004 698000 26604 708982
rect 29604 698000 30204 710862
rect 47604 710478 48204 711440
rect 47604 710242 47786 710478
rect 48022 710242 48204 710478
rect 47604 710158 48204 710242
rect 47604 709922 47786 710158
rect 48022 709922 48204 710158
rect 44004 708598 44604 709560
rect 44004 708362 44186 708598
rect 44422 708362 44604 708598
rect 44004 708278 44604 708362
rect 44004 708042 44186 708278
rect 44422 708042 44604 708278
rect 40404 706718 41004 707680
rect 40404 706482 40586 706718
rect 40822 706482 41004 706718
rect 40404 706398 41004 706482
rect 40404 706162 40586 706398
rect 40822 706162 41004 706398
rect 36804 704838 37404 705800
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 701792 37404 704282
rect 36804 701728 36832 701792
rect 36896 701728 36912 701792
rect 36976 701728 36992 701792
rect 37056 701728 37072 701792
rect 37136 701728 37152 701792
rect 37216 701728 37232 701792
rect 37296 701728 37312 701792
rect 37376 701728 37404 701792
rect 36804 700704 37404 701728
rect 36804 700640 36832 700704
rect 36896 700640 36912 700704
rect 36976 700640 36992 700704
rect 37056 700640 37072 700704
rect 37136 700640 37152 700704
rect 37216 700640 37232 700704
rect 37296 700640 37312 700704
rect 37376 700640 37404 700704
rect 36804 699616 37404 700640
rect 36804 699552 36832 699616
rect 36896 699552 36912 699616
rect 36976 699552 36992 699616
rect 37056 699552 37072 699616
rect 37136 699552 37152 699616
rect 37216 699552 37232 699616
rect 37296 699552 37312 699616
rect 37376 699552 37404 699616
rect 36804 698528 37404 699552
rect 36804 698464 36832 698528
rect 36896 698464 36912 698528
rect 36976 698464 36992 698528
rect 37056 698464 37072 698528
rect 37136 698464 37152 698528
rect 37216 698464 37232 698528
rect 37296 698464 37312 698528
rect 37376 698464 37404 698528
rect 36804 697952 37404 698464
rect 40404 698000 41004 706162
rect 44004 698000 44604 708042
rect 47604 698000 48204 709922
rect 65604 711418 66204 711440
rect 65604 711182 65786 711418
rect 66022 711182 66204 711418
rect 65604 711098 66204 711182
rect 65604 710862 65786 711098
rect 66022 710862 66204 711098
rect 62004 709538 62604 709560
rect 62004 709302 62186 709538
rect 62422 709302 62604 709538
rect 62004 709218 62604 709302
rect 62004 708982 62186 709218
rect 62422 708982 62604 709218
rect 58404 707658 59004 707680
rect 58404 707422 58586 707658
rect 58822 707422 59004 707658
rect 58404 707338 59004 707422
rect 58404 707102 58586 707338
rect 58822 707102 59004 707338
rect 54804 705778 55404 705800
rect 54804 705542 54986 705778
rect 55222 705542 55404 705778
rect 54804 705458 55404 705542
rect 54804 705222 54986 705458
rect 55222 705222 55404 705458
rect 54804 701248 55404 705222
rect 54804 701184 54832 701248
rect 54896 701184 54912 701248
rect 54976 701184 54992 701248
rect 55056 701184 55072 701248
rect 55136 701184 55152 701248
rect 55216 701184 55232 701248
rect 55296 701184 55312 701248
rect 55376 701184 55404 701248
rect 54804 700160 55404 701184
rect 54804 700096 54832 700160
rect 54896 700096 54912 700160
rect 54976 700096 54992 700160
rect 55056 700096 55072 700160
rect 55136 700096 55152 700160
rect 55216 700096 55232 700160
rect 55296 700096 55312 700160
rect 55376 700096 55404 700160
rect 54804 699072 55404 700096
rect 54804 699008 54832 699072
rect 54896 699008 54912 699072
rect 54976 699008 54992 699072
rect 55056 699008 55072 699072
rect 55136 699008 55152 699072
rect 55216 699008 55232 699072
rect 55296 699008 55312 699072
rect 55376 699008 55404 699072
rect 54804 697952 55404 699008
rect 58404 698000 59004 707102
rect 62004 698000 62604 708982
rect 65604 698000 66204 710862
rect 83604 710478 84204 711440
rect 83604 710242 83786 710478
rect 84022 710242 84204 710478
rect 83604 710158 84204 710242
rect 83604 709922 83786 710158
rect 84022 709922 84204 710158
rect 80004 708598 80604 709560
rect 80004 708362 80186 708598
rect 80422 708362 80604 708598
rect 80004 708278 80604 708362
rect 80004 708042 80186 708278
rect 80422 708042 80604 708278
rect 76404 706718 77004 707680
rect 76404 706482 76586 706718
rect 76822 706482 77004 706718
rect 76404 706398 77004 706482
rect 76404 706162 76586 706398
rect 76822 706162 77004 706398
rect 72804 704838 73404 705800
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 701792 73404 704282
rect 72804 701728 72832 701792
rect 72896 701728 72912 701792
rect 72976 701728 72992 701792
rect 73056 701728 73072 701792
rect 73136 701728 73152 701792
rect 73216 701728 73232 701792
rect 73296 701728 73312 701792
rect 73376 701728 73404 701792
rect 72804 700704 73404 701728
rect 72804 700640 72832 700704
rect 72896 700640 72912 700704
rect 72976 700640 72992 700704
rect 73056 700640 73072 700704
rect 73136 700640 73152 700704
rect 73216 700640 73232 700704
rect 73296 700640 73312 700704
rect 73376 700640 73404 700704
rect 72804 699616 73404 700640
rect 72804 699552 72832 699616
rect 72896 699552 72912 699616
rect 72976 699552 72992 699616
rect 73056 699552 73072 699616
rect 73136 699552 73152 699616
rect 73216 699552 73232 699616
rect 73296 699552 73312 699616
rect 73376 699552 73404 699616
rect 72804 698528 73404 699552
rect 72804 698464 72832 698528
rect 72896 698464 72912 698528
rect 72976 698464 72992 698528
rect 73056 698464 73072 698528
rect 73136 698464 73152 698528
rect 73216 698464 73232 698528
rect 73296 698464 73312 698528
rect 73376 698464 73404 698528
rect 71819 698324 71885 698325
rect 71819 698260 71820 698324
rect 71884 698260 71885 698324
rect 71819 698259 71885 698260
rect 15331 695332 15397 695333
rect 15331 695268 15332 695332
rect 15396 695268 15397 695332
rect 15331 695267 15397 695268
rect 15334 694517 15394 695267
rect 15331 694516 15397 694517
rect 15331 694452 15332 694516
rect 15396 694452 15397 694516
rect 15331 694451 15397 694452
rect 42011 694516 42077 694517
rect 42011 694452 42012 694516
rect 42076 694452 42077 694516
rect 42011 694451 42077 694452
rect 42014 694245 42074 694451
rect 9627 694244 9693 694245
rect 9627 694180 9628 694244
rect 9692 694180 9693 694244
rect 9627 694179 9693 694180
rect 42011 694244 42077 694245
rect 42011 694180 42012 694244
rect 42076 694180 42077 694244
rect 42011 694179 42077 694180
rect 64827 694244 64893 694245
rect 64827 694180 64828 694244
rect 64892 694180 64893 694244
rect 64827 694179 64893 694180
rect 9630 693973 9690 694179
rect 37227 694108 37293 694109
rect 37227 694044 37228 694108
rect 37292 694044 37293 694108
rect 37227 694043 37293 694044
rect 41275 694108 41341 694109
rect 41275 694044 41276 694108
rect 41340 694044 41341 694108
rect 41275 694043 41341 694044
rect 41459 694108 41525 694109
rect 41459 694044 41460 694108
rect 41524 694044 41525 694108
rect 41459 694043 41525 694044
rect 9627 693972 9693 693973
rect 9627 693908 9628 693972
rect 9692 693908 9693 693972
rect 9627 693907 9693 693908
rect 19011 693972 19077 693973
rect 19011 693908 19012 693972
rect 19076 693908 19077 693972
rect 27291 693972 27357 693973
rect 27291 693970 27292 693972
rect 19011 693907 19077 693908
rect 27110 693910 27292 693970
rect 19014 692698 19074 693907
rect 27110 692698 27170 693910
rect 27291 693908 27292 693910
rect 27356 693908 27357 693972
rect 27291 693907 27357 693908
rect 28947 693972 29013 693973
rect 28947 693908 28948 693972
rect 29012 693970 29013 693972
rect 29012 693910 29194 693970
rect 29012 693908 29013 693910
rect 28947 693907 29013 693908
rect 29134 693837 29194 693910
rect 37230 693837 37290 694043
rect 41278 693970 41338 694043
rect 41462 693970 41522 694043
rect 64830 693973 64890 694179
rect 41278 693910 41522 693970
rect 64827 693972 64893 693973
rect 64827 693908 64828 693972
rect 64892 693908 64893 693972
rect 64827 693907 64893 693908
rect 71822 693837 71882 698259
rect 72804 697952 73404 698464
rect 76404 698000 77004 706162
rect 80004 698000 80604 708042
rect 83604 698000 84204 709922
rect 101604 711418 102204 711440
rect 101604 711182 101786 711418
rect 102022 711182 102204 711418
rect 101604 711098 102204 711182
rect 101604 710862 101786 711098
rect 102022 710862 102204 711098
rect 98004 709538 98604 709560
rect 98004 709302 98186 709538
rect 98422 709302 98604 709538
rect 98004 709218 98604 709302
rect 98004 708982 98186 709218
rect 98422 708982 98604 709218
rect 94404 707658 95004 707680
rect 94404 707422 94586 707658
rect 94822 707422 95004 707658
rect 94404 707338 95004 707422
rect 94404 707102 94586 707338
rect 94822 707102 95004 707338
rect 90804 705778 91404 705800
rect 90804 705542 90986 705778
rect 91222 705542 91404 705778
rect 90804 705458 91404 705542
rect 90804 705222 90986 705458
rect 91222 705222 91404 705458
rect 90804 701248 91404 705222
rect 90804 701184 90832 701248
rect 90896 701184 90912 701248
rect 90976 701184 90992 701248
rect 91056 701184 91072 701248
rect 91136 701184 91152 701248
rect 91216 701184 91232 701248
rect 91296 701184 91312 701248
rect 91376 701184 91404 701248
rect 90804 700160 91404 701184
rect 90804 700096 90832 700160
rect 90896 700096 90912 700160
rect 90976 700096 90992 700160
rect 91056 700096 91072 700160
rect 91136 700096 91152 700160
rect 91216 700096 91232 700160
rect 91296 700096 91312 700160
rect 91376 700096 91404 700160
rect 90804 699072 91404 700096
rect 90804 699008 90832 699072
rect 90896 699008 90912 699072
rect 90976 699008 90992 699072
rect 91056 699008 91072 699072
rect 91136 699008 91152 699072
rect 91216 699008 91232 699072
rect 91296 699008 91312 699072
rect 91376 699008 91404 699072
rect 86723 698868 86789 698869
rect 86723 698804 86724 698868
rect 86788 698804 86789 698868
rect 86723 698803 86789 698804
rect 85251 694516 85317 694517
rect 85251 694452 85252 694516
rect 85316 694452 85317 694516
rect 85251 694451 85317 694452
rect 79915 694380 79981 694381
rect 79915 694316 79916 694380
rect 79980 694316 79981 694380
rect 79915 694315 79981 694316
rect 80099 694380 80165 694381
rect 80099 694316 80100 694380
rect 80164 694316 80165 694380
rect 80099 694315 80165 694316
rect 76971 694244 77037 694245
rect 76971 694180 76972 694244
rect 77036 694180 77037 694244
rect 79918 694242 79978 694315
rect 80102 694242 80162 694315
rect 79918 694182 80162 694242
rect 76971 694179 77037 694180
rect 29131 693836 29197 693837
rect 29131 693772 29132 693836
rect 29196 693772 29197 693836
rect 29131 693771 29197 693772
rect 37227 693836 37293 693837
rect 37227 693772 37228 693836
rect 37292 693772 37293 693836
rect 37227 693771 37293 693772
rect 71819 693836 71885 693837
rect 71819 693772 71820 693836
rect 71884 693772 71885 693836
rect 71819 693771 71885 693772
rect 76974 692698 77034 694179
rect 85254 692698 85314 694451
rect 86726 694245 86786 698803
rect 90804 697952 91404 699008
rect 94404 698000 95004 707102
rect 98004 698000 98604 708982
rect 101604 698000 102204 710862
rect 119604 710478 120204 711440
rect 119604 710242 119786 710478
rect 120022 710242 120204 710478
rect 119604 710158 120204 710242
rect 119604 709922 119786 710158
rect 120022 709922 120204 710158
rect 116004 708598 116604 709560
rect 116004 708362 116186 708598
rect 116422 708362 116604 708598
rect 116004 708278 116604 708362
rect 116004 708042 116186 708278
rect 116422 708042 116604 708278
rect 112404 706718 113004 707680
rect 112404 706482 112586 706718
rect 112822 706482 113004 706718
rect 112404 706398 113004 706482
rect 112404 706162 112586 706398
rect 112822 706162 113004 706398
rect 108804 704838 109404 705800
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 701792 109404 704282
rect 108804 701728 108832 701792
rect 108896 701728 108912 701792
rect 108976 701728 108992 701792
rect 109056 701728 109072 701792
rect 109136 701728 109152 701792
rect 109216 701728 109232 701792
rect 109296 701728 109312 701792
rect 109376 701728 109404 701792
rect 108804 700704 109404 701728
rect 108804 700640 108832 700704
rect 108896 700640 108912 700704
rect 108976 700640 108992 700704
rect 109056 700640 109072 700704
rect 109136 700640 109152 700704
rect 109216 700640 109232 700704
rect 109296 700640 109312 700704
rect 109376 700640 109404 700704
rect 108804 699616 109404 700640
rect 108804 699552 108832 699616
rect 108896 699552 108912 699616
rect 108976 699552 108992 699616
rect 109056 699552 109072 699616
rect 109136 699552 109152 699616
rect 109216 699552 109232 699616
rect 109296 699552 109312 699616
rect 109376 699552 109404 699616
rect 108804 698528 109404 699552
rect 108804 698464 108832 698528
rect 108896 698464 108912 698528
rect 108976 698464 108992 698528
rect 109056 698464 109072 698528
rect 109136 698464 109152 698528
rect 109216 698464 109232 698528
rect 109296 698464 109312 698528
rect 109376 698464 109404 698528
rect 108804 697952 109404 698464
rect 112404 698000 113004 706162
rect 116004 698000 116604 708042
rect 119604 698000 120204 709922
rect 137604 711418 138204 711440
rect 137604 711182 137786 711418
rect 138022 711182 138204 711418
rect 137604 711098 138204 711182
rect 137604 710862 137786 711098
rect 138022 710862 138204 711098
rect 134004 709538 134604 709560
rect 134004 709302 134186 709538
rect 134422 709302 134604 709538
rect 134004 709218 134604 709302
rect 134004 708982 134186 709218
rect 134422 708982 134604 709218
rect 130404 707658 131004 707680
rect 130404 707422 130586 707658
rect 130822 707422 131004 707658
rect 130404 707338 131004 707422
rect 130404 707102 130586 707338
rect 130822 707102 131004 707338
rect 126804 705778 127404 705800
rect 126804 705542 126986 705778
rect 127222 705542 127404 705778
rect 126804 705458 127404 705542
rect 126804 705222 126986 705458
rect 127222 705222 127404 705458
rect 126804 701248 127404 705222
rect 126804 701184 126832 701248
rect 126896 701184 126912 701248
rect 126976 701184 126992 701248
rect 127056 701184 127072 701248
rect 127136 701184 127152 701248
rect 127216 701184 127232 701248
rect 127296 701184 127312 701248
rect 127376 701184 127404 701248
rect 126804 700160 127404 701184
rect 126804 700096 126832 700160
rect 126896 700096 126912 700160
rect 126976 700096 126992 700160
rect 127056 700096 127072 700160
rect 127136 700096 127152 700160
rect 127216 700096 127232 700160
rect 127296 700096 127312 700160
rect 127376 700096 127404 700160
rect 126804 699072 127404 700096
rect 126804 699008 126832 699072
rect 126896 699008 126912 699072
rect 126976 699008 126992 699072
rect 127056 699008 127072 699072
rect 127136 699008 127152 699072
rect 127216 699008 127232 699072
rect 127296 699008 127312 699072
rect 127376 699008 127404 699072
rect 126804 697952 127404 699008
rect 130404 698000 131004 707102
rect 134004 698000 134604 708982
rect 137604 698000 138204 710862
rect 155604 710478 156204 711440
rect 155604 710242 155786 710478
rect 156022 710242 156204 710478
rect 155604 710158 156204 710242
rect 155604 709922 155786 710158
rect 156022 709922 156204 710158
rect 152004 708598 152604 709560
rect 152004 708362 152186 708598
rect 152422 708362 152604 708598
rect 152004 708278 152604 708362
rect 152004 708042 152186 708278
rect 152422 708042 152604 708278
rect 148404 706718 149004 707680
rect 148404 706482 148586 706718
rect 148822 706482 149004 706718
rect 148404 706398 149004 706482
rect 148404 706162 148586 706398
rect 148822 706162 149004 706398
rect 144804 704838 145404 705800
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 701792 145404 704282
rect 144804 701728 144832 701792
rect 144896 701728 144912 701792
rect 144976 701728 144992 701792
rect 145056 701728 145072 701792
rect 145136 701728 145152 701792
rect 145216 701728 145232 701792
rect 145296 701728 145312 701792
rect 145376 701728 145404 701792
rect 144804 700704 145404 701728
rect 144804 700640 144832 700704
rect 144896 700640 144912 700704
rect 144976 700640 144992 700704
rect 145056 700640 145072 700704
rect 145136 700640 145152 700704
rect 145216 700640 145232 700704
rect 145296 700640 145312 700704
rect 145376 700640 145404 700704
rect 144804 699616 145404 700640
rect 144804 699552 144832 699616
rect 144896 699552 144912 699616
rect 144976 699552 144992 699616
rect 145056 699552 145072 699616
rect 145136 699552 145152 699616
rect 145216 699552 145232 699616
rect 145296 699552 145312 699616
rect 145376 699552 145404 699616
rect 144804 698528 145404 699552
rect 144804 698464 144832 698528
rect 144896 698464 144912 698528
rect 144976 698464 144992 698528
rect 145056 698464 145072 698528
rect 145136 698464 145152 698528
rect 145216 698464 145232 698528
rect 145296 698464 145312 698528
rect 145376 698464 145404 698528
rect 144804 697952 145404 698464
rect 148404 698000 149004 706162
rect 152004 698000 152604 708042
rect 155604 698000 156204 709922
rect 173604 711418 174204 711440
rect 173604 711182 173786 711418
rect 174022 711182 174204 711418
rect 173604 711098 174204 711182
rect 173604 710862 173786 711098
rect 174022 710862 174204 711098
rect 170004 709538 170604 709560
rect 170004 709302 170186 709538
rect 170422 709302 170604 709538
rect 170004 709218 170604 709302
rect 170004 708982 170186 709218
rect 170422 708982 170604 709218
rect 166404 707658 167004 707680
rect 166404 707422 166586 707658
rect 166822 707422 167004 707658
rect 166404 707338 167004 707422
rect 166404 707102 166586 707338
rect 166822 707102 167004 707338
rect 162804 705778 163404 705800
rect 162804 705542 162986 705778
rect 163222 705542 163404 705778
rect 162804 705458 163404 705542
rect 162804 705222 162986 705458
rect 163222 705222 163404 705458
rect 162804 701248 163404 705222
rect 162804 701184 162832 701248
rect 162896 701184 162912 701248
rect 162976 701184 162992 701248
rect 163056 701184 163072 701248
rect 163136 701184 163152 701248
rect 163216 701184 163232 701248
rect 163296 701184 163312 701248
rect 163376 701184 163404 701248
rect 162804 700160 163404 701184
rect 162804 700096 162832 700160
rect 162896 700096 162912 700160
rect 162976 700096 162992 700160
rect 163056 700096 163072 700160
rect 163136 700096 163152 700160
rect 163216 700096 163232 700160
rect 163296 700096 163312 700160
rect 163376 700096 163404 700160
rect 162804 699072 163404 700096
rect 162804 699008 162832 699072
rect 162896 699008 162912 699072
rect 162976 699008 162992 699072
rect 163056 699008 163072 699072
rect 163136 699008 163152 699072
rect 163216 699008 163232 699072
rect 163296 699008 163312 699072
rect 163376 699008 163404 699072
rect 162804 697952 163404 699008
rect 166404 698000 167004 707102
rect 170004 698000 170604 708982
rect 173604 698000 174204 710862
rect 191604 710478 192204 711440
rect 191604 710242 191786 710478
rect 192022 710242 192204 710478
rect 191604 710158 192204 710242
rect 191604 709922 191786 710158
rect 192022 709922 192204 710158
rect 188004 708598 188604 709560
rect 188004 708362 188186 708598
rect 188422 708362 188604 708598
rect 188004 708278 188604 708362
rect 188004 708042 188186 708278
rect 188422 708042 188604 708278
rect 184404 706718 185004 707680
rect 184404 706482 184586 706718
rect 184822 706482 185004 706718
rect 184404 706398 185004 706482
rect 184404 706162 184586 706398
rect 184822 706162 185004 706398
rect 180804 704838 181404 705800
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 701792 181404 704282
rect 180804 701728 180832 701792
rect 180896 701728 180912 701792
rect 180976 701728 180992 701792
rect 181056 701728 181072 701792
rect 181136 701728 181152 701792
rect 181216 701728 181232 701792
rect 181296 701728 181312 701792
rect 181376 701728 181404 701792
rect 180804 700704 181404 701728
rect 180804 700640 180832 700704
rect 180896 700640 180912 700704
rect 180976 700640 180992 700704
rect 181056 700640 181072 700704
rect 181136 700640 181152 700704
rect 181216 700640 181232 700704
rect 181296 700640 181312 700704
rect 181376 700640 181404 700704
rect 180804 699616 181404 700640
rect 180804 699552 180832 699616
rect 180896 699552 180912 699616
rect 180976 699552 180992 699616
rect 181056 699552 181072 699616
rect 181136 699552 181152 699616
rect 181216 699552 181232 699616
rect 181296 699552 181312 699616
rect 181376 699552 181404 699616
rect 180804 698528 181404 699552
rect 180804 698464 180832 698528
rect 180896 698464 180912 698528
rect 180976 698464 180992 698528
rect 181056 698464 181072 698528
rect 181136 698464 181152 698528
rect 181216 698464 181232 698528
rect 181296 698464 181312 698528
rect 181376 698464 181404 698528
rect 180804 697952 181404 698464
rect 184404 698000 185004 706162
rect 188004 698000 188604 708042
rect 191604 698000 192204 709922
rect 209604 711418 210204 711440
rect 209604 711182 209786 711418
rect 210022 711182 210204 711418
rect 209604 711098 210204 711182
rect 209604 710862 209786 711098
rect 210022 710862 210204 711098
rect 206004 709538 206604 709560
rect 206004 709302 206186 709538
rect 206422 709302 206604 709538
rect 206004 709218 206604 709302
rect 206004 708982 206186 709218
rect 206422 708982 206604 709218
rect 202404 707658 203004 707680
rect 202404 707422 202586 707658
rect 202822 707422 203004 707658
rect 202404 707338 203004 707422
rect 202404 707102 202586 707338
rect 202822 707102 203004 707338
rect 198804 705778 199404 705800
rect 198804 705542 198986 705778
rect 199222 705542 199404 705778
rect 198804 705458 199404 705542
rect 198804 705222 198986 705458
rect 199222 705222 199404 705458
rect 198804 701248 199404 705222
rect 198804 701184 198832 701248
rect 198896 701184 198912 701248
rect 198976 701184 198992 701248
rect 199056 701184 199072 701248
rect 199136 701184 199152 701248
rect 199216 701184 199232 701248
rect 199296 701184 199312 701248
rect 199376 701184 199404 701248
rect 198804 700160 199404 701184
rect 198804 700096 198832 700160
rect 198896 700096 198912 700160
rect 198976 700096 198992 700160
rect 199056 700096 199072 700160
rect 199136 700096 199152 700160
rect 199216 700096 199232 700160
rect 199296 700096 199312 700160
rect 199376 700096 199404 700160
rect 198804 699072 199404 700096
rect 198804 699008 198832 699072
rect 198896 699008 198912 699072
rect 198976 699008 198992 699072
rect 199056 699008 199072 699072
rect 199136 699008 199152 699072
rect 199216 699008 199232 699072
rect 199296 699008 199312 699072
rect 199376 699008 199404 699072
rect 198804 697952 199404 699008
rect 202404 698000 203004 707102
rect 206004 698000 206604 708982
rect 209604 698000 210204 710862
rect 227604 710478 228204 711440
rect 227604 710242 227786 710478
rect 228022 710242 228204 710478
rect 227604 710158 228204 710242
rect 227604 709922 227786 710158
rect 228022 709922 228204 710158
rect 224004 708598 224604 709560
rect 224004 708362 224186 708598
rect 224422 708362 224604 708598
rect 224004 708278 224604 708362
rect 224004 708042 224186 708278
rect 224422 708042 224604 708278
rect 220404 706718 221004 707680
rect 220404 706482 220586 706718
rect 220822 706482 221004 706718
rect 220404 706398 221004 706482
rect 220404 706162 220586 706398
rect 220822 706162 221004 706398
rect 216804 704838 217404 705800
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 701792 217404 704282
rect 216804 701728 216832 701792
rect 216896 701728 216912 701792
rect 216976 701728 216992 701792
rect 217056 701728 217072 701792
rect 217136 701728 217152 701792
rect 217216 701728 217232 701792
rect 217296 701728 217312 701792
rect 217376 701728 217404 701792
rect 216804 700704 217404 701728
rect 216804 700640 216832 700704
rect 216896 700640 216912 700704
rect 216976 700640 216992 700704
rect 217056 700640 217072 700704
rect 217136 700640 217152 700704
rect 217216 700640 217232 700704
rect 217296 700640 217312 700704
rect 217376 700640 217404 700704
rect 216804 699616 217404 700640
rect 216804 699552 216832 699616
rect 216896 699552 216912 699616
rect 216976 699552 216992 699616
rect 217056 699552 217072 699616
rect 217136 699552 217152 699616
rect 217216 699552 217232 699616
rect 217296 699552 217312 699616
rect 217376 699552 217404 699616
rect 216804 698528 217404 699552
rect 216804 698464 216832 698528
rect 216896 698464 216912 698528
rect 216976 698464 216992 698528
rect 217056 698464 217072 698528
rect 217136 698464 217152 698528
rect 217216 698464 217232 698528
rect 217296 698464 217312 698528
rect 217376 698464 217404 698528
rect 216804 697952 217404 698464
rect 220404 698000 221004 706162
rect 224004 698000 224604 708042
rect 227604 698000 228204 709922
rect 245604 711418 246204 711440
rect 245604 711182 245786 711418
rect 246022 711182 246204 711418
rect 245604 711098 246204 711182
rect 245604 710862 245786 711098
rect 246022 710862 246204 711098
rect 242004 709538 242604 709560
rect 242004 709302 242186 709538
rect 242422 709302 242604 709538
rect 242004 709218 242604 709302
rect 242004 708982 242186 709218
rect 242422 708982 242604 709218
rect 238404 707658 239004 707680
rect 238404 707422 238586 707658
rect 238822 707422 239004 707658
rect 238404 707338 239004 707422
rect 238404 707102 238586 707338
rect 238822 707102 239004 707338
rect 234804 705778 235404 705800
rect 234804 705542 234986 705778
rect 235222 705542 235404 705778
rect 234804 705458 235404 705542
rect 234804 705222 234986 705458
rect 235222 705222 235404 705458
rect 234804 701248 235404 705222
rect 234804 701184 234832 701248
rect 234896 701184 234912 701248
rect 234976 701184 234992 701248
rect 235056 701184 235072 701248
rect 235136 701184 235152 701248
rect 235216 701184 235232 701248
rect 235296 701184 235312 701248
rect 235376 701184 235404 701248
rect 234804 700160 235404 701184
rect 234804 700096 234832 700160
rect 234896 700096 234912 700160
rect 234976 700096 234992 700160
rect 235056 700096 235072 700160
rect 235136 700096 235152 700160
rect 235216 700096 235232 700160
rect 235296 700096 235312 700160
rect 235376 700096 235404 700160
rect 234804 699072 235404 700096
rect 234804 699008 234832 699072
rect 234896 699008 234912 699072
rect 234976 699008 234992 699072
rect 235056 699008 235072 699072
rect 235136 699008 235152 699072
rect 235216 699008 235232 699072
rect 235296 699008 235312 699072
rect 235376 699008 235404 699072
rect 234804 697952 235404 699008
rect 238404 698000 239004 707102
rect 242004 698000 242604 708982
rect 245604 698000 246204 710862
rect 263604 710478 264204 711440
rect 263604 710242 263786 710478
rect 264022 710242 264204 710478
rect 263604 710158 264204 710242
rect 263604 709922 263786 710158
rect 264022 709922 264204 710158
rect 260004 708598 260604 709560
rect 260004 708362 260186 708598
rect 260422 708362 260604 708598
rect 260004 708278 260604 708362
rect 260004 708042 260186 708278
rect 260422 708042 260604 708278
rect 256404 706718 257004 707680
rect 256404 706482 256586 706718
rect 256822 706482 257004 706718
rect 256404 706398 257004 706482
rect 256404 706162 256586 706398
rect 256822 706162 257004 706398
rect 252804 704838 253404 705800
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 701792 253404 704282
rect 252804 701728 252832 701792
rect 252896 701728 252912 701792
rect 252976 701728 252992 701792
rect 253056 701728 253072 701792
rect 253136 701728 253152 701792
rect 253216 701728 253232 701792
rect 253296 701728 253312 701792
rect 253376 701728 253404 701792
rect 252804 700704 253404 701728
rect 252804 700640 252832 700704
rect 252896 700640 252912 700704
rect 252976 700640 252992 700704
rect 253056 700640 253072 700704
rect 253136 700640 253152 700704
rect 253216 700640 253232 700704
rect 253296 700640 253312 700704
rect 253376 700640 253404 700704
rect 252804 699616 253404 700640
rect 252804 699552 252832 699616
rect 252896 699552 252912 699616
rect 252976 699552 252992 699616
rect 253056 699552 253072 699616
rect 253136 699552 253152 699616
rect 253216 699552 253232 699616
rect 253296 699552 253312 699616
rect 253376 699552 253404 699616
rect 252804 698528 253404 699552
rect 252804 698464 252832 698528
rect 252896 698464 252912 698528
rect 252976 698464 252992 698528
rect 253056 698464 253072 698528
rect 253136 698464 253152 698528
rect 253216 698464 253232 698528
rect 253296 698464 253312 698528
rect 253376 698464 253404 698528
rect 252804 697952 253404 698464
rect 256404 698000 257004 706162
rect 260004 698000 260604 708042
rect 263604 698000 264204 709922
rect 281604 711418 282204 711440
rect 281604 711182 281786 711418
rect 282022 711182 282204 711418
rect 281604 711098 282204 711182
rect 281604 710862 281786 711098
rect 282022 710862 282204 711098
rect 278004 709538 278604 709560
rect 278004 709302 278186 709538
rect 278422 709302 278604 709538
rect 278004 709218 278604 709302
rect 278004 708982 278186 709218
rect 278422 708982 278604 709218
rect 274404 707658 275004 707680
rect 274404 707422 274586 707658
rect 274822 707422 275004 707658
rect 274404 707338 275004 707422
rect 274404 707102 274586 707338
rect 274822 707102 275004 707338
rect 270804 705778 271404 705800
rect 270804 705542 270986 705778
rect 271222 705542 271404 705778
rect 270804 705458 271404 705542
rect 270804 705222 270986 705458
rect 271222 705222 271404 705458
rect 270804 701248 271404 705222
rect 270804 701184 270832 701248
rect 270896 701184 270912 701248
rect 270976 701184 270992 701248
rect 271056 701184 271072 701248
rect 271136 701184 271152 701248
rect 271216 701184 271232 701248
rect 271296 701184 271312 701248
rect 271376 701184 271404 701248
rect 270804 700160 271404 701184
rect 270804 700096 270832 700160
rect 270896 700096 270912 700160
rect 270976 700096 270992 700160
rect 271056 700096 271072 700160
rect 271136 700096 271152 700160
rect 271216 700096 271232 700160
rect 271296 700096 271312 700160
rect 271376 700096 271404 700160
rect 270804 699072 271404 700096
rect 270804 699008 270832 699072
rect 270896 699008 270912 699072
rect 270976 699008 270992 699072
rect 271056 699008 271072 699072
rect 271136 699008 271152 699072
rect 271216 699008 271232 699072
rect 271296 699008 271312 699072
rect 271376 699008 271404 699072
rect 270804 697952 271404 699008
rect 274404 698000 275004 707102
rect 278004 698000 278604 708982
rect 281604 698000 282204 710862
rect 299604 710478 300204 711440
rect 299604 710242 299786 710478
rect 300022 710242 300204 710478
rect 299604 710158 300204 710242
rect 299604 709922 299786 710158
rect 300022 709922 300204 710158
rect 296004 708598 296604 709560
rect 296004 708362 296186 708598
rect 296422 708362 296604 708598
rect 296004 708278 296604 708362
rect 296004 708042 296186 708278
rect 296422 708042 296604 708278
rect 292404 706718 293004 707680
rect 292404 706482 292586 706718
rect 292822 706482 293004 706718
rect 292404 706398 293004 706482
rect 292404 706162 292586 706398
rect 292822 706162 293004 706398
rect 288804 704838 289404 705800
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 701792 289404 704282
rect 288804 701728 288832 701792
rect 288896 701728 288912 701792
rect 288976 701728 288992 701792
rect 289056 701728 289072 701792
rect 289136 701728 289152 701792
rect 289216 701728 289232 701792
rect 289296 701728 289312 701792
rect 289376 701728 289404 701792
rect 288804 700704 289404 701728
rect 288804 700640 288832 700704
rect 288896 700640 288912 700704
rect 288976 700640 288992 700704
rect 289056 700640 289072 700704
rect 289136 700640 289152 700704
rect 289216 700640 289232 700704
rect 289296 700640 289312 700704
rect 289376 700640 289404 700704
rect 288804 699616 289404 700640
rect 288804 699552 288832 699616
rect 288896 699552 288912 699616
rect 288976 699552 288992 699616
rect 289056 699552 289072 699616
rect 289136 699552 289152 699616
rect 289216 699552 289232 699616
rect 289296 699552 289312 699616
rect 289376 699552 289404 699616
rect 282867 699140 282933 699141
rect 282867 699076 282868 699140
rect 282932 699076 282933 699140
rect 282867 699075 282933 699076
rect 282870 698597 282930 699075
rect 282867 698596 282933 698597
rect 282867 698532 282868 698596
rect 282932 698532 282933 698596
rect 282867 698531 282933 698532
rect 288804 698528 289404 699552
rect 288804 698464 288832 698528
rect 288896 698464 288912 698528
rect 288976 698464 288992 698528
rect 289056 698464 289072 698528
rect 289136 698464 289152 698528
rect 289216 698464 289232 698528
rect 289296 698464 289312 698528
rect 289376 698464 289404 698528
rect 288804 697952 289404 698464
rect 292404 698000 293004 706162
rect 296004 698000 296604 708042
rect 299604 698000 300204 709922
rect 317604 711418 318204 711440
rect 317604 711182 317786 711418
rect 318022 711182 318204 711418
rect 317604 711098 318204 711182
rect 317604 710862 317786 711098
rect 318022 710862 318204 711098
rect 314004 709538 314604 709560
rect 314004 709302 314186 709538
rect 314422 709302 314604 709538
rect 314004 709218 314604 709302
rect 314004 708982 314186 709218
rect 314422 708982 314604 709218
rect 310404 707658 311004 707680
rect 310404 707422 310586 707658
rect 310822 707422 311004 707658
rect 310404 707338 311004 707422
rect 310404 707102 310586 707338
rect 310822 707102 311004 707338
rect 306804 705778 307404 705800
rect 306804 705542 306986 705778
rect 307222 705542 307404 705778
rect 306804 705458 307404 705542
rect 306804 705222 306986 705458
rect 307222 705222 307404 705458
rect 306804 701248 307404 705222
rect 306804 701184 306832 701248
rect 306896 701184 306912 701248
rect 306976 701184 306992 701248
rect 307056 701184 307072 701248
rect 307136 701184 307152 701248
rect 307216 701184 307232 701248
rect 307296 701184 307312 701248
rect 307376 701184 307404 701248
rect 306804 700160 307404 701184
rect 306804 700096 306832 700160
rect 306896 700096 306912 700160
rect 306976 700096 306992 700160
rect 307056 700096 307072 700160
rect 307136 700096 307152 700160
rect 307216 700096 307232 700160
rect 307296 700096 307312 700160
rect 307376 700096 307404 700160
rect 306804 699072 307404 700096
rect 306804 699008 306832 699072
rect 306896 699008 306912 699072
rect 306976 699008 306992 699072
rect 307056 699008 307072 699072
rect 307136 699008 307152 699072
rect 307216 699008 307232 699072
rect 307296 699008 307312 699072
rect 307376 699008 307404 699072
rect 306804 697952 307404 699008
rect 310404 698000 311004 707102
rect 314004 698000 314604 708982
rect 317604 698000 318204 710862
rect 335604 710478 336204 711440
rect 335604 710242 335786 710478
rect 336022 710242 336204 710478
rect 335604 710158 336204 710242
rect 335604 709922 335786 710158
rect 336022 709922 336204 710158
rect 332004 708598 332604 709560
rect 332004 708362 332186 708598
rect 332422 708362 332604 708598
rect 332004 708278 332604 708362
rect 332004 708042 332186 708278
rect 332422 708042 332604 708278
rect 328404 706718 329004 707680
rect 328404 706482 328586 706718
rect 328822 706482 329004 706718
rect 328404 706398 329004 706482
rect 328404 706162 328586 706398
rect 328822 706162 329004 706398
rect 324804 704838 325404 705800
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 701792 325404 704282
rect 324804 701728 324832 701792
rect 324896 701728 324912 701792
rect 324976 701728 324992 701792
rect 325056 701728 325072 701792
rect 325136 701728 325152 701792
rect 325216 701728 325232 701792
rect 325296 701728 325312 701792
rect 325376 701728 325404 701792
rect 324804 700704 325404 701728
rect 324804 700640 324832 700704
rect 324896 700640 324912 700704
rect 324976 700640 324992 700704
rect 325056 700640 325072 700704
rect 325136 700640 325152 700704
rect 325216 700640 325232 700704
rect 325296 700640 325312 700704
rect 325376 700640 325404 700704
rect 324804 699616 325404 700640
rect 324804 699552 324832 699616
rect 324896 699552 324912 699616
rect 324976 699552 324992 699616
rect 325056 699552 325072 699616
rect 325136 699552 325152 699616
rect 325216 699552 325232 699616
rect 325296 699552 325312 699616
rect 325376 699552 325404 699616
rect 324804 698528 325404 699552
rect 324804 698464 324832 698528
rect 324896 698464 324912 698528
rect 324976 698464 324992 698528
rect 325056 698464 325072 698528
rect 325136 698464 325152 698528
rect 325216 698464 325232 698528
rect 325296 698464 325312 698528
rect 325376 698464 325404 698528
rect 324804 697952 325404 698464
rect 328404 698000 329004 706162
rect 332004 698000 332604 708042
rect 335604 698000 336204 709922
rect 353604 711418 354204 711440
rect 353604 711182 353786 711418
rect 354022 711182 354204 711418
rect 353604 711098 354204 711182
rect 353604 710862 353786 711098
rect 354022 710862 354204 711098
rect 350004 709538 350604 709560
rect 350004 709302 350186 709538
rect 350422 709302 350604 709538
rect 350004 709218 350604 709302
rect 350004 708982 350186 709218
rect 350422 708982 350604 709218
rect 346404 707658 347004 707680
rect 346404 707422 346586 707658
rect 346822 707422 347004 707658
rect 346404 707338 347004 707422
rect 346404 707102 346586 707338
rect 346822 707102 347004 707338
rect 342804 705778 343404 705800
rect 342804 705542 342986 705778
rect 343222 705542 343404 705778
rect 342804 705458 343404 705542
rect 342804 705222 342986 705458
rect 343222 705222 343404 705458
rect 342804 701248 343404 705222
rect 342804 701184 342832 701248
rect 342896 701184 342912 701248
rect 342976 701184 342992 701248
rect 343056 701184 343072 701248
rect 343136 701184 343152 701248
rect 343216 701184 343232 701248
rect 343296 701184 343312 701248
rect 343376 701184 343404 701248
rect 342804 700160 343404 701184
rect 342804 700096 342832 700160
rect 342896 700096 342912 700160
rect 342976 700096 342992 700160
rect 343056 700096 343072 700160
rect 343136 700096 343152 700160
rect 343216 700096 343232 700160
rect 343296 700096 343312 700160
rect 343376 700096 343404 700160
rect 342804 699072 343404 700096
rect 342804 699008 342832 699072
rect 342896 699008 342912 699072
rect 342976 699008 342992 699072
rect 343056 699008 343072 699072
rect 343136 699008 343152 699072
rect 343216 699008 343232 699072
rect 343296 699008 343312 699072
rect 343376 699008 343404 699072
rect 342804 697952 343404 699008
rect 346404 698000 347004 707102
rect 350004 698000 350604 708982
rect 353604 698000 354204 710862
rect 371604 710478 372204 711440
rect 371604 710242 371786 710478
rect 372022 710242 372204 710478
rect 371604 710158 372204 710242
rect 371604 709922 371786 710158
rect 372022 709922 372204 710158
rect 368004 708598 368604 709560
rect 368004 708362 368186 708598
rect 368422 708362 368604 708598
rect 368004 708278 368604 708362
rect 368004 708042 368186 708278
rect 368422 708042 368604 708278
rect 364404 706718 365004 707680
rect 364404 706482 364586 706718
rect 364822 706482 365004 706718
rect 364404 706398 365004 706482
rect 364404 706162 364586 706398
rect 364822 706162 365004 706398
rect 360804 704838 361404 705800
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 701792 361404 704282
rect 360804 701728 360832 701792
rect 360896 701728 360912 701792
rect 360976 701728 360992 701792
rect 361056 701728 361072 701792
rect 361136 701728 361152 701792
rect 361216 701728 361232 701792
rect 361296 701728 361312 701792
rect 361376 701728 361404 701792
rect 360804 700704 361404 701728
rect 360804 700640 360832 700704
rect 360896 700640 360912 700704
rect 360976 700640 360992 700704
rect 361056 700640 361072 700704
rect 361136 700640 361152 700704
rect 361216 700640 361232 700704
rect 361296 700640 361312 700704
rect 361376 700640 361404 700704
rect 360804 699616 361404 700640
rect 360804 699552 360832 699616
rect 360896 699552 360912 699616
rect 360976 699552 360992 699616
rect 361056 699552 361072 699616
rect 361136 699552 361152 699616
rect 361216 699552 361232 699616
rect 361296 699552 361312 699616
rect 361376 699552 361404 699616
rect 360804 698528 361404 699552
rect 360804 698464 360832 698528
rect 360896 698464 360912 698528
rect 360976 698464 360992 698528
rect 361056 698464 361072 698528
rect 361136 698464 361152 698528
rect 361216 698464 361232 698528
rect 361296 698464 361312 698528
rect 361376 698464 361404 698528
rect 360804 697952 361404 698464
rect 364404 698000 365004 706162
rect 368004 698000 368604 708042
rect 371604 698000 372204 709922
rect 389604 711418 390204 711440
rect 389604 711182 389786 711418
rect 390022 711182 390204 711418
rect 389604 711098 390204 711182
rect 389604 710862 389786 711098
rect 390022 710862 390204 711098
rect 386004 709538 386604 709560
rect 386004 709302 386186 709538
rect 386422 709302 386604 709538
rect 386004 709218 386604 709302
rect 386004 708982 386186 709218
rect 386422 708982 386604 709218
rect 382404 707658 383004 707680
rect 382404 707422 382586 707658
rect 382822 707422 383004 707658
rect 382404 707338 383004 707422
rect 382404 707102 382586 707338
rect 382822 707102 383004 707338
rect 378804 705778 379404 705800
rect 378804 705542 378986 705778
rect 379222 705542 379404 705778
rect 378804 705458 379404 705542
rect 378804 705222 378986 705458
rect 379222 705222 379404 705458
rect 378804 701248 379404 705222
rect 378804 701184 378832 701248
rect 378896 701184 378912 701248
rect 378976 701184 378992 701248
rect 379056 701184 379072 701248
rect 379136 701184 379152 701248
rect 379216 701184 379232 701248
rect 379296 701184 379312 701248
rect 379376 701184 379404 701248
rect 378804 700160 379404 701184
rect 378804 700096 378832 700160
rect 378896 700096 378912 700160
rect 378976 700096 378992 700160
rect 379056 700096 379072 700160
rect 379136 700096 379152 700160
rect 379216 700096 379232 700160
rect 379296 700096 379312 700160
rect 379376 700096 379404 700160
rect 378804 699072 379404 700096
rect 378804 699008 378832 699072
rect 378896 699008 378912 699072
rect 378976 699008 378992 699072
rect 379056 699008 379072 699072
rect 379136 699008 379152 699072
rect 379216 699008 379232 699072
rect 379296 699008 379312 699072
rect 379376 699008 379404 699072
rect 378804 697952 379404 699008
rect 382404 698000 383004 707102
rect 386004 698000 386604 708982
rect 389604 698000 390204 710862
rect 407604 710478 408204 711440
rect 407604 710242 407786 710478
rect 408022 710242 408204 710478
rect 407604 710158 408204 710242
rect 407604 709922 407786 710158
rect 408022 709922 408204 710158
rect 404004 708598 404604 709560
rect 404004 708362 404186 708598
rect 404422 708362 404604 708598
rect 404004 708278 404604 708362
rect 404004 708042 404186 708278
rect 404422 708042 404604 708278
rect 400404 706718 401004 707680
rect 400404 706482 400586 706718
rect 400822 706482 401004 706718
rect 400404 706398 401004 706482
rect 400404 706162 400586 706398
rect 400822 706162 401004 706398
rect 396804 704838 397404 705800
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 701792 397404 704282
rect 396804 701728 396832 701792
rect 396896 701728 396912 701792
rect 396976 701728 396992 701792
rect 397056 701728 397072 701792
rect 397136 701728 397152 701792
rect 397216 701728 397232 701792
rect 397296 701728 397312 701792
rect 397376 701728 397404 701792
rect 396804 700704 397404 701728
rect 396804 700640 396832 700704
rect 396896 700640 396912 700704
rect 396976 700640 396992 700704
rect 397056 700640 397072 700704
rect 397136 700640 397152 700704
rect 397216 700640 397232 700704
rect 397296 700640 397312 700704
rect 397376 700640 397404 700704
rect 396804 699616 397404 700640
rect 396804 699552 396832 699616
rect 396896 699552 396912 699616
rect 396976 699552 396992 699616
rect 397056 699552 397072 699616
rect 397136 699552 397152 699616
rect 397216 699552 397232 699616
rect 397296 699552 397312 699616
rect 397376 699552 397404 699616
rect 396804 698528 397404 699552
rect 396804 698464 396832 698528
rect 396896 698464 396912 698528
rect 396976 698464 396992 698528
rect 397056 698464 397072 698528
rect 397136 698464 397152 698528
rect 397216 698464 397232 698528
rect 397296 698464 397312 698528
rect 397376 698464 397404 698528
rect 396804 697952 397404 698464
rect 400404 698000 401004 706162
rect 404004 698000 404604 708042
rect 407604 698000 408204 709922
rect 425604 711418 426204 711440
rect 425604 711182 425786 711418
rect 426022 711182 426204 711418
rect 425604 711098 426204 711182
rect 425604 710862 425786 711098
rect 426022 710862 426204 711098
rect 422004 709538 422604 709560
rect 422004 709302 422186 709538
rect 422422 709302 422604 709538
rect 422004 709218 422604 709302
rect 422004 708982 422186 709218
rect 422422 708982 422604 709218
rect 418404 707658 419004 707680
rect 418404 707422 418586 707658
rect 418822 707422 419004 707658
rect 418404 707338 419004 707422
rect 418404 707102 418586 707338
rect 418822 707102 419004 707338
rect 414804 705778 415404 705800
rect 414804 705542 414986 705778
rect 415222 705542 415404 705778
rect 414804 705458 415404 705542
rect 414804 705222 414986 705458
rect 415222 705222 415404 705458
rect 414804 701248 415404 705222
rect 414804 701184 414832 701248
rect 414896 701184 414912 701248
rect 414976 701184 414992 701248
rect 415056 701184 415072 701248
rect 415136 701184 415152 701248
rect 415216 701184 415232 701248
rect 415296 701184 415312 701248
rect 415376 701184 415404 701248
rect 414804 700160 415404 701184
rect 414804 700096 414832 700160
rect 414896 700096 414912 700160
rect 414976 700096 414992 700160
rect 415056 700096 415072 700160
rect 415136 700096 415152 700160
rect 415216 700096 415232 700160
rect 415296 700096 415312 700160
rect 415376 700096 415404 700160
rect 414804 699072 415404 700096
rect 414804 699008 414832 699072
rect 414896 699008 414912 699072
rect 414976 699008 414992 699072
rect 415056 699008 415072 699072
rect 415136 699008 415152 699072
rect 415216 699008 415232 699072
rect 415296 699008 415312 699072
rect 415376 699008 415404 699072
rect 414804 697952 415404 699008
rect 418404 698000 419004 707102
rect 422004 698000 422604 708982
rect 425604 698000 426204 710862
rect 443604 710478 444204 711440
rect 443604 710242 443786 710478
rect 444022 710242 444204 710478
rect 443604 710158 444204 710242
rect 443604 709922 443786 710158
rect 444022 709922 444204 710158
rect 440004 708598 440604 709560
rect 440004 708362 440186 708598
rect 440422 708362 440604 708598
rect 440004 708278 440604 708362
rect 440004 708042 440186 708278
rect 440422 708042 440604 708278
rect 436404 706718 437004 707680
rect 436404 706482 436586 706718
rect 436822 706482 437004 706718
rect 436404 706398 437004 706482
rect 436404 706162 436586 706398
rect 436822 706162 437004 706398
rect 432804 704838 433404 705800
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 701792 433404 704282
rect 432804 701728 432832 701792
rect 432896 701728 432912 701792
rect 432976 701728 432992 701792
rect 433056 701728 433072 701792
rect 433136 701728 433152 701792
rect 433216 701728 433232 701792
rect 433296 701728 433312 701792
rect 433376 701728 433404 701792
rect 432804 700704 433404 701728
rect 432804 700640 432832 700704
rect 432896 700640 432912 700704
rect 432976 700640 432992 700704
rect 433056 700640 433072 700704
rect 433136 700640 433152 700704
rect 433216 700640 433232 700704
rect 433296 700640 433312 700704
rect 433376 700640 433404 700704
rect 432804 699616 433404 700640
rect 432804 699552 432832 699616
rect 432896 699552 432912 699616
rect 432976 699552 432992 699616
rect 433056 699552 433072 699616
rect 433136 699552 433152 699616
rect 433216 699552 433232 699616
rect 433296 699552 433312 699616
rect 433376 699552 433404 699616
rect 432804 698528 433404 699552
rect 432804 698464 432832 698528
rect 432896 698464 432912 698528
rect 432976 698464 432992 698528
rect 433056 698464 433072 698528
rect 433136 698464 433152 698528
rect 433216 698464 433232 698528
rect 433296 698464 433312 698528
rect 433376 698464 433404 698528
rect 432804 697952 433404 698464
rect 436404 698000 437004 706162
rect 440004 698000 440604 708042
rect 443604 698000 444204 709922
rect 461604 711418 462204 711440
rect 461604 711182 461786 711418
rect 462022 711182 462204 711418
rect 461604 711098 462204 711182
rect 461604 710862 461786 711098
rect 462022 710862 462204 711098
rect 458004 709538 458604 709560
rect 458004 709302 458186 709538
rect 458422 709302 458604 709538
rect 458004 709218 458604 709302
rect 458004 708982 458186 709218
rect 458422 708982 458604 709218
rect 454404 707658 455004 707680
rect 454404 707422 454586 707658
rect 454822 707422 455004 707658
rect 454404 707338 455004 707422
rect 454404 707102 454586 707338
rect 454822 707102 455004 707338
rect 450804 705778 451404 705800
rect 450804 705542 450986 705778
rect 451222 705542 451404 705778
rect 450804 705458 451404 705542
rect 450804 705222 450986 705458
rect 451222 705222 451404 705458
rect 450804 701248 451404 705222
rect 450804 701184 450832 701248
rect 450896 701184 450912 701248
rect 450976 701184 450992 701248
rect 451056 701184 451072 701248
rect 451136 701184 451152 701248
rect 451216 701184 451232 701248
rect 451296 701184 451312 701248
rect 451376 701184 451404 701248
rect 450804 700160 451404 701184
rect 450804 700096 450832 700160
rect 450896 700096 450912 700160
rect 450976 700096 450992 700160
rect 451056 700096 451072 700160
rect 451136 700096 451152 700160
rect 451216 700096 451232 700160
rect 451296 700096 451312 700160
rect 451376 700096 451404 700160
rect 450804 699072 451404 700096
rect 450804 699008 450832 699072
rect 450896 699008 450912 699072
rect 450976 699008 450992 699072
rect 451056 699008 451072 699072
rect 451136 699008 451152 699072
rect 451216 699008 451232 699072
rect 451296 699008 451312 699072
rect 451376 699008 451404 699072
rect 447179 698868 447245 698869
rect 447179 698804 447180 698868
rect 447244 698804 447245 698868
rect 447179 698803 447245 698804
rect 179643 695332 179709 695333
rect 179643 695268 179644 695332
rect 179708 695268 179709 695332
rect 179643 695267 179709 695268
rect 137323 694924 137389 694925
rect 137323 694860 137324 694924
rect 137388 694860 137389 694924
rect 137323 694859 137389 694860
rect 141923 694924 141989 694925
rect 141923 694860 141924 694924
rect 141988 694860 141989 694924
rect 141923 694859 141989 694860
rect 134931 694788 134997 694789
rect 134931 694724 134932 694788
rect 134996 694724 134997 694788
rect 134931 694723 134997 694724
rect 106227 694652 106293 694653
rect 106227 694588 106228 694652
rect 106292 694588 106293 694652
rect 106227 694587 106293 694588
rect 115795 694652 115861 694653
rect 115795 694588 115796 694652
rect 115860 694588 115861 694652
rect 115795 694587 115861 694588
rect 106230 694381 106290 694587
rect 98315 694380 98381 694381
rect 98315 694316 98316 694380
rect 98380 694378 98381 694380
rect 98867 694380 98933 694381
rect 98867 694378 98868 694380
rect 98380 694318 98868 694378
rect 98380 694316 98381 694318
rect 98315 694315 98381 694316
rect 98867 694316 98868 694318
rect 98932 694316 98933 694380
rect 98867 694315 98933 694316
rect 106227 694380 106293 694381
rect 106227 694316 106228 694380
rect 106292 694316 106293 694380
rect 106227 694315 106293 694316
rect 106411 694380 106477 694381
rect 106411 694316 106412 694380
rect 106476 694316 106477 694380
rect 106411 694315 106477 694316
rect 86723 694244 86789 694245
rect 86723 694180 86724 694244
rect 86788 694180 86789 694244
rect 86723 694179 86789 694180
rect 106227 694108 106293 694109
rect 102734 694046 103346 694106
rect 86907 693972 86973 693973
rect 86907 693908 86908 693972
rect 86972 693970 86973 693972
rect 87091 693972 87157 693973
rect 87091 693970 87092 693972
rect 86972 693910 87092 693970
rect 86972 693908 86973 693910
rect 86907 693907 86973 693908
rect 87091 693908 87092 693910
rect 87156 693908 87157 693972
rect 87091 693907 87157 693908
rect 102734 693701 102794 694046
rect 103286 693701 103346 694046
rect 106227 694044 106228 694108
rect 106292 694106 106293 694108
rect 106414 694106 106474 694315
rect 106292 694046 106474 694106
rect 106292 694044 106293 694046
rect 106227 694043 106293 694044
rect 115798 693970 115858 694587
rect 134934 694517 134994 694723
rect 115979 694516 116045 694517
rect 115979 694452 115980 694516
rect 116044 694452 116045 694516
rect 115979 694451 116045 694452
rect 130331 694516 130397 694517
rect 130331 694452 130332 694516
rect 130396 694452 130397 694516
rect 130331 694451 130397 694452
rect 134931 694516 134997 694517
rect 134931 694452 134932 694516
rect 134996 694452 134997 694516
rect 134931 694451 134997 694452
rect 115982 693970 116042 694451
rect 120579 694380 120645 694381
rect 120579 694316 120580 694380
rect 120644 694316 120645 694380
rect 120579 694315 120645 694316
rect 120582 694109 120642 694315
rect 130334 694109 130394 694451
rect 137326 694109 137386 694859
rect 138243 694788 138309 694789
rect 138243 694724 138244 694788
rect 138308 694724 138309 694788
rect 138243 694723 138309 694724
rect 138246 694109 138306 694723
rect 141926 694381 141986 694859
rect 142107 694788 142173 694789
rect 142107 694724 142108 694788
rect 142172 694724 142173 694788
rect 142107 694723 142173 694724
rect 151675 694788 151741 694789
rect 151675 694724 151676 694788
rect 151740 694724 151741 694788
rect 151675 694723 151741 694724
rect 152779 694788 152845 694789
rect 152779 694724 152780 694788
rect 152844 694724 152845 694788
rect 152779 694723 152845 694724
rect 159403 694788 159469 694789
rect 159403 694724 159404 694788
rect 159468 694724 159469 694788
rect 159403 694723 159469 694724
rect 142110 694381 142170 694723
rect 151678 694517 151738 694723
rect 151862 694590 152106 694650
rect 151862 694517 151922 694590
rect 151675 694516 151741 694517
rect 151675 694452 151676 694516
rect 151740 694452 151741 694516
rect 151675 694451 151741 694452
rect 151859 694516 151925 694517
rect 151859 694452 151860 694516
rect 151924 694452 151925 694516
rect 151859 694451 151925 694452
rect 141923 694380 141989 694381
rect 141923 694316 141924 694380
rect 141988 694316 141989 694380
rect 141923 694315 141989 694316
rect 142107 694380 142173 694381
rect 142107 694316 142108 694380
rect 142172 694316 142173 694380
rect 142107 694315 142173 694316
rect 146891 694380 146957 694381
rect 146891 694316 146892 694380
rect 146956 694316 146957 694380
rect 146891 694315 146957 694316
rect 146894 694109 146954 694315
rect 152046 694109 152106 694590
rect 152782 694381 152842 694723
rect 152779 694380 152845 694381
rect 152779 694316 152780 694380
rect 152844 694316 152845 694380
rect 152779 694315 152845 694316
rect 159406 694109 159466 694723
rect 164187 694652 164253 694653
rect 164187 694588 164188 694652
rect 164252 694588 164253 694652
rect 164187 694587 164253 694588
rect 173571 694652 173637 694653
rect 173571 694588 173572 694652
rect 173636 694588 173637 694652
rect 173571 694587 173637 694588
rect 176699 694652 176765 694653
rect 176699 694588 176700 694652
rect 176764 694588 176765 694652
rect 176699 694587 176765 694588
rect 164190 694381 164250 694587
rect 166947 694516 167013 694517
rect 166947 694452 166948 694516
rect 167012 694452 167013 694516
rect 173574 694514 173634 694587
rect 173574 694454 173818 694514
rect 166947 694451 167013 694452
rect 164187 694380 164253 694381
rect 164187 694316 164188 694380
rect 164252 694316 164253 694380
rect 164187 694315 164253 694316
rect 166950 694109 167010 694451
rect 173758 694245 173818 694454
rect 176702 694245 176762 694587
rect 176883 694516 176949 694517
rect 176883 694452 176884 694516
rect 176948 694452 176949 694516
rect 176883 694451 176949 694452
rect 173755 694244 173821 694245
rect 173755 694180 173756 694244
rect 173820 694180 173821 694244
rect 173755 694179 173821 694180
rect 176699 694244 176765 694245
rect 176699 694180 176700 694244
rect 176764 694180 176765 694244
rect 176699 694179 176765 694180
rect 176886 694109 176946 694451
rect 179646 694381 179706 695267
rect 231899 695060 231965 695061
rect 231899 694996 231900 695060
rect 231964 694996 231965 695060
rect 231899 694995 231965 694996
rect 236867 695060 236933 695061
rect 236867 694996 236868 695060
rect 236932 694996 236933 695060
rect 236867 694995 236933 694996
rect 251219 695060 251285 695061
rect 251219 694996 251220 695060
rect 251284 694996 251285 695060
rect 251219 694995 251285 694996
rect 256187 695060 256253 695061
rect 256187 694996 256188 695060
rect 256252 694996 256253 695060
rect 256187 694995 256253 694996
rect 357387 695060 357453 695061
rect 357387 694996 357388 695060
rect 357452 694996 357453 695060
rect 357387 694995 357453 694996
rect 362171 695060 362237 695061
rect 362171 694996 362172 695060
rect 362236 694996 362237 695060
rect 362171 694995 362237 694996
rect 434667 695060 434733 695061
rect 434667 694996 434668 695060
rect 434732 694996 434733 695060
rect 434667 694995 434733 694996
rect 439451 695060 439517 695061
rect 439451 694996 439452 695060
rect 439516 694996 439517 695060
rect 439451 694995 439517 694996
rect 196203 694924 196269 694925
rect 196203 694860 196204 694924
rect 196268 694860 196269 694924
rect 196203 694859 196269 694860
rect 202459 694924 202525 694925
rect 202459 694860 202460 694924
rect 202524 694860 202525 694924
rect 202459 694859 202525 694860
rect 186267 694652 186333 694653
rect 186267 694588 186268 694652
rect 186332 694588 186333 694652
rect 186267 694587 186333 694588
rect 179643 694380 179709 694381
rect 179643 694316 179644 694380
rect 179708 694316 179709 694380
rect 179643 694315 179709 694316
rect 186083 694380 186149 694381
rect 186083 694316 186084 694380
rect 186148 694316 186149 694380
rect 186083 694315 186149 694316
rect 186086 694109 186146 694315
rect 186270 694109 186330 694587
rect 196206 694381 196266 694859
rect 202462 694514 202522 694859
rect 222147 694788 222213 694789
rect 222147 694724 222148 694788
rect 222212 694724 222213 694788
rect 222147 694723 222213 694724
rect 226931 694788 226997 694789
rect 226931 694724 226932 694788
rect 226996 694724 226997 694788
rect 226931 694723 226997 694724
rect 215339 694652 215405 694653
rect 215339 694588 215340 694652
rect 215404 694588 215405 694652
rect 215339 694587 215405 694588
rect 202643 694516 202709 694517
rect 202643 694514 202644 694516
rect 202462 694454 202644 694514
rect 202643 694452 202644 694454
rect 202708 694452 202709 694516
rect 202643 694451 202709 694452
rect 214971 694516 215037 694517
rect 214971 694452 214972 694516
rect 215036 694452 215037 694516
rect 214971 694451 215037 694452
rect 196203 694380 196269 694381
rect 196203 694316 196204 694380
rect 196268 694316 196269 694380
rect 196203 694315 196269 694316
rect 214974 694109 215034 694451
rect 215342 694109 215402 694587
rect 215523 694516 215589 694517
rect 215523 694452 215524 694516
rect 215588 694514 215589 694516
rect 215588 694454 215770 694514
rect 215588 694452 215589 694454
rect 215523 694451 215589 694452
rect 215710 694245 215770 694454
rect 222150 694381 222210 694723
rect 224355 694652 224421 694653
rect 224355 694588 224356 694652
rect 224420 694588 224421 694652
rect 224355 694587 224421 694588
rect 222147 694380 222213 694381
rect 222147 694316 222148 694380
rect 222212 694316 222213 694380
rect 222147 694315 222213 694316
rect 215707 694244 215773 694245
rect 215707 694180 215708 694244
rect 215772 694180 215773 694244
rect 215707 694179 215773 694180
rect 224358 694109 224418 694587
rect 226934 694381 226994 694723
rect 231902 694381 231962 694995
rect 236683 694788 236749 694789
rect 236683 694724 236684 694788
rect 236748 694724 236749 694788
rect 236683 694723 236749 694724
rect 226931 694380 226997 694381
rect 226931 694316 226932 694380
rect 226996 694316 226997 694380
rect 226931 694315 226997 694316
rect 231899 694380 231965 694381
rect 231899 694316 231900 694380
rect 231964 694316 231965 694380
rect 231899 694315 231965 694316
rect 232083 694380 232149 694381
rect 232083 694316 232084 694380
rect 232148 694316 232149 694380
rect 232083 694315 232149 694316
rect 235947 694380 236013 694381
rect 235947 694316 235948 694380
rect 236012 694316 236013 694380
rect 235947 694315 236013 694316
rect 120579 694108 120645 694109
rect 120579 694044 120580 694108
rect 120644 694044 120645 694108
rect 120579 694043 120645 694044
rect 130331 694108 130397 694109
rect 130331 694044 130332 694108
rect 130396 694044 130397 694108
rect 130331 694043 130397 694044
rect 137323 694108 137389 694109
rect 137323 694044 137324 694108
rect 137388 694044 137389 694108
rect 137323 694043 137389 694044
rect 138243 694108 138309 694109
rect 138243 694044 138244 694108
rect 138308 694044 138309 694108
rect 138243 694043 138309 694044
rect 146891 694108 146957 694109
rect 146891 694044 146892 694108
rect 146956 694044 146957 694108
rect 146891 694043 146957 694044
rect 152043 694108 152109 694109
rect 152043 694044 152044 694108
rect 152108 694044 152109 694108
rect 152043 694043 152109 694044
rect 159403 694108 159469 694109
rect 159403 694044 159404 694108
rect 159468 694044 159469 694108
rect 159403 694043 159469 694044
rect 166947 694108 167013 694109
rect 166947 694044 166948 694108
rect 167012 694044 167013 694108
rect 166947 694043 167013 694044
rect 176883 694108 176949 694109
rect 176883 694044 176884 694108
rect 176948 694044 176949 694108
rect 176883 694043 176949 694044
rect 185899 694108 185965 694109
rect 185899 694044 185900 694108
rect 185964 694044 185965 694108
rect 185899 694043 185965 694044
rect 186083 694108 186149 694109
rect 186083 694044 186084 694108
rect 186148 694044 186149 694108
rect 186083 694043 186149 694044
rect 186267 694108 186333 694109
rect 186267 694044 186268 694108
rect 186332 694044 186333 694108
rect 186267 694043 186333 694044
rect 186451 694108 186517 694109
rect 186451 694044 186452 694108
rect 186516 694044 186517 694108
rect 186451 694043 186517 694044
rect 205403 694108 205469 694109
rect 205403 694044 205404 694108
rect 205468 694106 205469 694108
rect 205955 694108 206021 694109
rect 205955 694106 205956 694108
rect 205468 694046 205956 694106
rect 205468 694044 205469 694046
rect 205403 694043 205469 694044
rect 205955 694044 205956 694046
rect 206020 694044 206021 694108
rect 205955 694043 206021 694044
rect 214971 694108 215037 694109
rect 214971 694044 214972 694108
rect 215036 694044 215037 694108
rect 214971 694043 215037 694044
rect 215339 694108 215405 694109
rect 215339 694044 215340 694108
rect 215404 694044 215405 694108
rect 215339 694043 215405 694044
rect 224355 694108 224421 694109
rect 224355 694044 224356 694108
rect 224420 694044 224421 694108
rect 224355 694043 224421 694044
rect 115798 693910 116042 693970
rect 185902 693970 185962 694043
rect 186454 693970 186514 694043
rect 185902 693910 186514 693970
rect 231899 693836 231965 693837
rect 231899 693772 231900 693836
rect 231964 693772 231965 693836
rect 231899 693771 231965 693772
rect 102731 693700 102797 693701
rect 102731 693636 102732 693700
rect 102796 693636 102797 693700
rect 102731 693635 102797 693636
rect 103283 693700 103349 693701
rect 103283 693636 103284 693700
rect 103348 693636 103349 693700
rect 103283 693635 103349 693636
rect 231902 692610 231962 693771
rect 232086 693701 232146 694315
rect 232635 693836 232701 693837
rect 232635 693772 232636 693836
rect 232700 693772 232701 693836
rect 232635 693771 232701 693772
rect 232083 693700 232149 693701
rect 232083 693636 232084 693700
rect 232148 693636 232149 693700
rect 232083 693635 232149 693636
rect 232638 692610 232698 693771
rect 235950 693701 236010 694315
rect 236686 694109 236746 694723
rect 236870 694245 236930 694995
rect 241099 694788 241165 694789
rect 241099 694724 241100 694788
rect 241164 694724 241165 694788
rect 241099 694723 241165 694724
rect 246067 694788 246133 694789
rect 246067 694724 246068 694788
rect 246132 694724 246133 694788
rect 246067 694723 246133 694724
rect 241102 694381 241162 694723
rect 243859 694652 243925 694653
rect 243859 694588 243860 694652
rect 243924 694588 243925 694652
rect 243859 694587 243925 694588
rect 241099 694380 241165 694381
rect 241099 694316 241100 694380
rect 241164 694316 241165 694380
rect 241099 694315 241165 694316
rect 236867 694244 236933 694245
rect 236867 694180 236868 694244
rect 236932 694180 236933 694244
rect 236867 694179 236933 694180
rect 243862 694109 243922 694587
rect 246070 694381 246130 694723
rect 251222 694381 251282 694995
rect 256003 694788 256069 694789
rect 256003 694724 256004 694788
rect 256068 694724 256069 694788
rect 256003 694723 256069 694724
rect 246067 694380 246133 694381
rect 246067 694316 246068 694380
rect 246132 694316 246133 694380
rect 246067 694315 246133 694316
rect 251219 694380 251285 694381
rect 251219 694316 251220 694380
rect 251284 694316 251285 694380
rect 251219 694315 251285 694316
rect 251403 694380 251469 694381
rect 251403 694316 251404 694380
rect 251468 694316 251469 694380
rect 251403 694315 251469 694316
rect 255267 694380 255333 694381
rect 255267 694316 255268 694380
rect 255332 694316 255333 694380
rect 255267 694315 255333 694316
rect 245699 694244 245765 694245
rect 245699 694180 245700 694244
rect 245764 694242 245765 694244
rect 246435 694244 246501 694245
rect 246435 694242 246436 694244
rect 245764 694182 246436 694242
rect 245764 694180 245765 694182
rect 245699 694179 245765 694180
rect 246435 694180 246436 694182
rect 246500 694180 246501 694244
rect 246435 694179 246501 694180
rect 236683 694108 236749 694109
rect 236683 694044 236684 694108
rect 236748 694044 236749 694108
rect 236683 694043 236749 694044
rect 243859 694108 243925 694109
rect 243859 694044 243860 694108
rect 243924 694044 243925 694108
rect 243859 694043 243925 694044
rect 251219 693836 251285 693837
rect 251219 693772 251220 693836
rect 251284 693772 251285 693836
rect 251219 693771 251285 693772
rect 235947 693700 236013 693701
rect 235947 693636 235948 693700
rect 236012 693636 236013 693700
rect 235947 693635 236013 693636
rect 231902 692550 232698 692610
rect 251222 692610 251282 693771
rect 251406 693701 251466 694315
rect 251955 693836 252021 693837
rect 251955 693772 251956 693836
rect 252020 693772 252021 693836
rect 251955 693771 252021 693772
rect 251403 693700 251469 693701
rect 251403 693636 251404 693700
rect 251468 693636 251469 693700
rect 251403 693635 251469 693636
rect 251958 692610 252018 693771
rect 255270 693701 255330 694315
rect 256006 694109 256066 694723
rect 256190 694245 256250 694995
rect 273115 694924 273181 694925
rect 273115 694860 273116 694924
rect 273180 694860 273181 694924
rect 273115 694859 273181 694860
rect 278819 694924 278885 694925
rect 278819 694860 278820 694924
rect 278884 694860 278885 694924
rect 278819 694859 278885 694860
rect 280107 694924 280173 694925
rect 280107 694860 280108 694924
rect 280172 694860 280173 694924
rect 280107 694859 280173 694860
rect 283235 694924 283301 694925
rect 283235 694860 283236 694924
rect 283300 694860 283301 694924
rect 283235 694859 283301 694860
rect 292803 694924 292869 694925
rect 292803 694860 292804 694924
rect 292868 694860 292869 694924
rect 292803 694859 292869 694860
rect 299059 694924 299125 694925
rect 299059 694860 299060 694924
rect 299124 694860 299125 694924
rect 299059 694859 299125 694860
rect 346347 694924 346413 694925
rect 346347 694860 346348 694924
rect 346412 694860 346413 694924
rect 346347 694859 346413 694860
rect 351315 694924 351381 694925
rect 351315 694860 351316 694924
rect 351380 694860 351381 694924
rect 351315 694859 351381 694860
rect 264283 694788 264349 694789
rect 264283 694724 264284 694788
rect 264348 694724 264349 694788
rect 264283 694723 264349 694724
rect 270355 694788 270421 694789
rect 270355 694724 270356 694788
rect 270420 694724 270421 694788
rect 270355 694723 270421 694724
rect 263179 694652 263245 694653
rect 263179 694588 263180 694652
rect 263244 694588 263245 694652
rect 263179 694587 263245 694588
rect 256187 694244 256253 694245
rect 256187 694180 256188 694244
rect 256252 694180 256253 694244
rect 256187 694179 256253 694180
rect 263182 694109 263242 694587
rect 264286 694245 264346 694723
rect 265571 694516 265637 694517
rect 265571 694452 265572 694516
rect 265636 694452 265637 694516
rect 265571 694451 265637 694452
rect 264283 694244 264349 694245
rect 264283 694180 264284 694244
rect 264348 694180 264349 694244
rect 264283 694179 264349 694180
rect 265574 694109 265634 694451
rect 270358 694245 270418 694723
rect 273118 694653 273178 694859
rect 273115 694652 273181 694653
rect 273115 694588 273116 694652
rect 273180 694588 273181 694652
rect 273115 694587 273181 694588
rect 270723 694380 270789 694381
rect 270723 694316 270724 694380
rect 270788 694316 270789 694380
rect 270723 694315 270789 694316
rect 270355 694244 270421 694245
rect 270355 694180 270356 694244
rect 270420 694180 270421 694244
rect 270726 694242 270786 694315
rect 278822 694245 278882 694859
rect 280110 694786 280170 694859
rect 279926 694726 280170 694786
rect 270355 694179 270421 694180
rect 270542 694182 270786 694242
rect 278819 694244 278885 694245
rect 270542 694109 270602 694182
rect 278819 694180 278820 694244
rect 278884 694180 278885 694244
rect 278819 694179 278885 694180
rect 279926 694109 279986 694726
rect 282683 694652 282749 694653
rect 282683 694588 282684 694652
rect 282748 694588 282749 694652
rect 282683 694587 282749 694588
rect 282686 694245 282746 694587
rect 283238 694381 283298 694859
rect 292806 694381 292866 694859
rect 299062 694514 299122 694859
rect 318747 694788 318813 694789
rect 318747 694724 318748 694788
rect 318812 694724 318813 694788
rect 318747 694723 318813 694724
rect 328315 694788 328381 694789
rect 328315 694724 328316 694788
rect 328380 694724 328381 694788
rect 328315 694723 328381 694724
rect 311939 694652 312005 694653
rect 311939 694588 311940 694652
rect 312004 694588 312005 694652
rect 311939 694587 312005 694588
rect 299243 694516 299309 694517
rect 299243 694514 299244 694516
rect 299062 694454 299244 694514
rect 299243 694452 299244 694454
rect 299308 694452 299309 694516
rect 299243 694451 299309 694452
rect 311571 694516 311637 694517
rect 311571 694452 311572 694516
rect 311636 694452 311637 694516
rect 311571 694451 311637 694452
rect 283051 694380 283117 694381
rect 283051 694316 283052 694380
rect 283116 694316 283117 694380
rect 283051 694315 283117 694316
rect 283235 694380 283301 694381
rect 283235 694316 283236 694380
rect 283300 694316 283301 694380
rect 283235 694315 283301 694316
rect 292803 694380 292869 694381
rect 292803 694316 292804 694380
rect 292868 694316 292869 694380
rect 292803 694315 292869 694316
rect 282683 694244 282749 694245
rect 282683 694180 282684 694244
rect 282748 694180 282749 694244
rect 282683 694179 282749 694180
rect 256003 694108 256069 694109
rect 256003 694044 256004 694108
rect 256068 694044 256069 694108
rect 256003 694043 256069 694044
rect 263179 694108 263245 694109
rect 263179 694044 263180 694108
rect 263244 694044 263245 694108
rect 263179 694043 263245 694044
rect 265571 694108 265637 694109
rect 265571 694044 265572 694108
rect 265636 694044 265637 694108
rect 265571 694043 265637 694044
rect 270539 694108 270605 694109
rect 270539 694044 270540 694108
rect 270604 694044 270605 694108
rect 270539 694043 270605 694044
rect 279923 694108 279989 694109
rect 279923 694044 279924 694108
rect 279988 694044 279989 694108
rect 283054 694106 283114 694315
rect 311574 694109 311634 694451
rect 311942 694109 312002 694587
rect 312123 694516 312189 694517
rect 312123 694452 312124 694516
rect 312188 694514 312189 694516
rect 312188 694454 312370 694514
rect 312188 694452 312189 694454
rect 312123 694451 312189 694452
rect 312310 694245 312370 694454
rect 318750 694381 318810 694723
rect 320955 694652 321021 694653
rect 320955 694588 320956 694652
rect 321020 694588 321021 694652
rect 320955 694587 321021 694588
rect 318747 694380 318813 694381
rect 318747 694316 318748 694380
rect 318812 694316 318813 694380
rect 318747 694315 318813 694316
rect 312307 694244 312373 694245
rect 312307 694180 312308 694244
rect 312372 694180 312373 694244
rect 312307 694179 312373 694180
rect 320958 694109 321018 694587
rect 328318 694381 328378 694723
rect 346350 694653 346410 694859
rect 350579 694788 350645 694789
rect 350579 694724 350580 694788
rect 350644 694724 350645 694788
rect 350579 694723 350645 694724
rect 332915 694652 332981 694653
rect 332915 694588 332916 694652
rect 332980 694588 332981 694652
rect 332915 694587 332981 694588
rect 338619 694652 338685 694653
rect 338619 694588 338620 694652
rect 338684 694588 338685 694652
rect 338619 694587 338685 694588
rect 340459 694652 340525 694653
rect 340459 694588 340460 694652
rect 340524 694588 340525 694652
rect 340459 694587 340525 694588
rect 346347 694652 346413 694653
rect 346347 694588 346348 694652
rect 346412 694588 346413 694652
rect 346347 694587 346413 694588
rect 328315 694380 328381 694381
rect 328315 694316 328316 694380
rect 328380 694316 328381 694380
rect 328315 694315 328381 694316
rect 332918 694109 332978 694587
rect 333099 694516 333165 694517
rect 333099 694452 333100 694516
rect 333164 694452 333165 694516
rect 333099 694451 333165 694452
rect 333102 694245 333162 694451
rect 338622 694381 338682 694587
rect 338619 694380 338685 694381
rect 338619 694316 338620 694380
rect 338684 694316 338685 694380
rect 338619 694315 338685 694316
rect 333099 694244 333165 694245
rect 333099 694180 333100 694244
rect 333164 694180 333165 694244
rect 333099 694179 333165 694180
rect 340462 694109 340522 694587
rect 341563 694516 341629 694517
rect 341563 694452 341564 694516
rect 341628 694452 341629 694516
rect 341563 694451 341629 694452
rect 341566 694245 341626 694451
rect 350395 694380 350461 694381
rect 350395 694316 350396 694380
rect 350460 694316 350461 694380
rect 350395 694315 350461 694316
rect 341563 694244 341629 694245
rect 341563 694180 341564 694244
rect 341628 694180 341629 694244
rect 341563 694179 341629 694180
rect 350398 694109 350458 694315
rect 350582 694245 350642 694723
rect 350763 694380 350829 694381
rect 350763 694316 350764 694380
rect 350828 694378 350829 694380
rect 351131 694380 351197 694381
rect 351131 694378 351132 694380
rect 350828 694318 351132 694378
rect 350828 694316 350829 694318
rect 350763 694315 350829 694316
rect 351131 694316 351132 694318
rect 351196 694316 351197 694380
rect 351131 694315 351197 694316
rect 351318 694245 351378 694859
rect 357390 694789 357450 694995
rect 357387 694788 357453 694789
rect 357387 694724 357388 694788
rect 357452 694724 357453 694788
rect 357387 694723 357453 694724
rect 359963 694652 360029 694653
rect 359963 694588 359964 694652
rect 360028 694588 360029 694652
rect 359963 694587 360029 694588
rect 359966 694245 360026 694587
rect 362174 694381 362234 694995
rect 370083 694924 370149 694925
rect 370083 694860 370084 694924
rect 370148 694860 370149 694924
rect 370083 694859 370149 694860
rect 376339 694924 376405 694925
rect 376339 694860 376340 694924
rect 376404 694860 376405 694924
rect 376339 694859 376405 694860
rect 389403 694924 389469 694925
rect 389403 694860 389404 694924
rect 389468 694860 389469 694924
rect 389403 694859 389469 694860
rect 395659 694924 395725 694925
rect 395659 694860 395660 694924
rect 395724 694860 395725 694924
rect 395659 694859 395725 694860
rect 370086 694381 370146 694859
rect 376342 694514 376402 694859
rect 376523 694516 376589 694517
rect 376523 694514 376524 694516
rect 376342 694454 376524 694514
rect 376523 694452 376524 694454
rect 376588 694452 376589 694516
rect 376523 694451 376589 694452
rect 389406 694381 389466 694859
rect 395662 694514 395722 694859
rect 434670 694789 434730 694995
rect 434667 694788 434733 694789
rect 434667 694724 434668 694788
rect 434732 694724 434733 694788
rect 434667 694723 434733 694724
rect 395843 694516 395909 694517
rect 395843 694514 395844 694516
rect 395662 694454 395844 694514
rect 395843 694452 395844 694454
rect 395908 694452 395909 694516
rect 427675 694516 427741 694517
rect 395843 694451 395909 694452
rect 417558 694454 417986 694514
rect 417558 694381 417618 694454
rect 362171 694380 362237 694381
rect 362171 694316 362172 694380
rect 362236 694316 362237 694380
rect 362171 694315 362237 694316
rect 370083 694380 370149 694381
rect 370083 694316 370084 694380
rect 370148 694316 370149 694380
rect 370083 694315 370149 694316
rect 389403 694380 389469 694381
rect 389403 694316 389404 694380
rect 389468 694316 389469 694380
rect 389403 694315 389469 694316
rect 417555 694380 417621 694381
rect 417555 694316 417556 694380
rect 417620 694316 417621 694380
rect 417555 694315 417621 694316
rect 417739 694380 417805 694381
rect 417739 694316 417740 694380
rect 417804 694316 417805 694380
rect 417926 694378 417986 694454
rect 427675 694452 427676 694516
rect 427740 694452 427741 694516
rect 427675 694451 427741 694452
rect 427859 694516 427925 694517
rect 427859 694452 427860 694516
rect 427924 694452 427925 694516
rect 427859 694451 427925 694452
rect 437243 694516 437309 694517
rect 437243 694452 437244 694516
rect 437308 694452 437309 694516
rect 437243 694451 437309 694452
rect 437427 694516 437493 694517
rect 437427 694452 437428 694516
rect 437492 694452 437493 694516
rect 437427 694451 437493 694452
rect 418475 694380 418541 694381
rect 418475 694378 418476 694380
rect 417926 694318 418476 694378
rect 417739 694315 417805 694316
rect 418475 694316 418476 694318
rect 418540 694316 418541 694380
rect 418475 694315 418541 694316
rect 350579 694244 350645 694245
rect 350579 694180 350580 694244
rect 350644 694180 350645 694244
rect 350579 694179 350645 694180
rect 351315 694244 351381 694245
rect 351315 694180 351316 694244
rect 351380 694180 351381 694244
rect 351315 694179 351381 694180
rect 359963 694244 360029 694245
rect 359963 694180 359964 694244
rect 360028 694180 360029 694244
rect 359963 694179 360029 694180
rect 410563 694244 410629 694245
rect 410563 694180 410564 694244
rect 410628 694180 410629 694244
rect 410563 694179 410629 694180
rect 414979 694244 415045 694245
rect 414979 694180 414980 694244
rect 415044 694180 415045 694244
rect 414979 694179 415045 694180
rect 283235 694108 283301 694109
rect 283235 694106 283236 694108
rect 283054 694046 283236 694106
rect 279923 694043 279989 694044
rect 283235 694044 283236 694046
rect 283300 694044 283301 694108
rect 283235 694043 283301 694044
rect 302003 694108 302069 694109
rect 302003 694044 302004 694108
rect 302068 694106 302069 694108
rect 302555 694108 302621 694109
rect 302555 694106 302556 694108
rect 302068 694046 302556 694106
rect 302068 694044 302069 694046
rect 302003 694043 302069 694044
rect 302555 694044 302556 694046
rect 302620 694044 302621 694108
rect 302555 694043 302621 694044
rect 311571 694108 311637 694109
rect 311571 694044 311572 694108
rect 311636 694044 311637 694108
rect 311571 694043 311637 694044
rect 311939 694108 312005 694109
rect 311939 694044 311940 694108
rect 312004 694044 312005 694108
rect 311939 694043 312005 694044
rect 320955 694108 321021 694109
rect 320955 694044 320956 694108
rect 321020 694044 321021 694108
rect 320955 694043 321021 694044
rect 332915 694108 332981 694109
rect 332915 694044 332916 694108
rect 332980 694044 332981 694108
rect 332915 694043 332981 694044
rect 340459 694108 340525 694109
rect 340459 694044 340460 694108
rect 340524 694044 340525 694108
rect 340459 694043 340525 694044
rect 350395 694108 350461 694109
rect 350395 694044 350396 694108
rect 350460 694044 350461 694108
rect 350395 694043 350461 694044
rect 379283 694108 379349 694109
rect 379283 694044 379284 694108
rect 379348 694106 379349 694108
rect 379835 694108 379901 694109
rect 379835 694106 379836 694108
rect 379348 694046 379836 694106
rect 379348 694044 379349 694046
rect 379283 694043 379349 694044
rect 379835 694044 379836 694046
rect 379900 694044 379901 694108
rect 379835 694043 379901 694044
rect 398603 694108 398669 694109
rect 398603 694044 398604 694108
rect 398668 694106 398669 694108
rect 399155 694108 399221 694109
rect 399155 694106 399156 694108
rect 398668 694046 399156 694106
rect 398668 694044 398669 694046
rect 398603 694043 398669 694044
rect 399155 694044 399156 694046
rect 399220 694044 399221 694108
rect 399155 694043 399221 694044
rect 410566 693973 410626 694179
rect 270539 693972 270605 693973
rect 270539 693908 270540 693972
rect 270604 693970 270605 693972
rect 270723 693972 270789 693973
rect 270723 693970 270724 693972
rect 270604 693910 270724 693970
rect 270604 693908 270605 693910
rect 270539 693907 270605 693908
rect 270723 693908 270724 693910
rect 270788 693908 270789 693972
rect 410563 693972 410629 693973
rect 270723 693907 270789 693908
rect 270910 693910 271338 693970
rect 270910 693701 270970 693910
rect 271278 693701 271338 693910
rect 410563 693908 410564 693972
rect 410628 693908 410629 693972
rect 414982 693970 415042 694179
rect 417742 694109 417802 694315
rect 427678 694109 427738 694451
rect 427862 694109 427922 694451
rect 437246 694109 437306 694451
rect 437430 694109 437490 694451
rect 439454 694381 439514 694995
rect 447182 694517 447242 698803
rect 450804 697952 451404 699008
rect 454404 698000 455004 707102
rect 458004 698000 458604 708982
rect 461604 698000 462204 710862
rect 479604 710478 480204 711440
rect 479604 710242 479786 710478
rect 480022 710242 480204 710478
rect 479604 710158 480204 710242
rect 479604 709922 479786 710158
rect 480022 709922 480204 710158
rect 476004 708598 476604 709560
rect 476004 708362 476186 708598
rect 476422 708362 476604 708598
rect 476004 708278 476604 708362
rect 476004 708042 476186 708278
rect 476422 708042 476604 708278
rect 472404 706718 473004 707680
rect 472404 706482 472586 706718
rect 472822 706482 473004 706718
rect 472404 706398 473004 706482
rect 472404 706162 472586 706398
rect 472822 706162 473004 706398
rect 468804 704838 469404 705800
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 701792 469404 704282
rect 468804 701728 468832 701792
rect 468896 701728 468912 701792
rect 468976 701728 468992 701792
rect 469056 701728 469072 701792
rect 469136 701728 469152 701792
rect 469216 701728 469232 701792
rect 469296 701728 469312 701792
rect 469376 701728 469404 701792
rect 468804 700704 469404 701728
rect 468804 700640 468832 700704
rect 468896 700640 468912 700704
rect 468976 700640 468992 700704
rect 469056 700640 469072 700704
rect 469136 700640 469152 700704
rect 469216 700640 469232 700704
rect 469296 700640 469312 700704
rect 469376 700640 469404 700704
rect 468804 699616 469404 700640
rect 468804 699552 468832 699616
rect 468896 699552 468912 699616
rect 468976 699552 468992 699616
rect 469056 699552 469072 699616
rect 469136 699552 469152 699616
rect 469216 699552 469232 699616
rect 469296 699552 469312 699616
rect 469376 699552 469404 699616
rect 468804 698528 469404 699552
rect 468804 698464 468832 698528
rect 468896 698464 468912 698528
rect 468976 698464 468992 698528
rect 469056 698464 469072 698528
rect 469136 698464 469152 698528
rect 469216 698464 469232 698528
rect 469296 698464 469312 698528
rect 469376 698464 469404 698528
rect 468804 697952 469404 698464
rect 472404 698000 473004 706162
rect 476004 698000 476604 708042
rect 479604 698000 480204 709922
rect 497604 711418 498204 711440
rect 497604 711182 497786 711418
rect 498022 711182 498204 711418
rect 497604 711098 498204 711182
rect 497604 710862 497786 711098
rect 498022 710862 498204 711098
rect 494004 709538 494604 709560
rect 494004 709302 494186 709538
rect 494422 709302 494604 709538
rect 494004 709218 494604 709302
rect 494004 708982 494186 709218
rect 494422 708982 494604 709218
rect 490404 707658 491004 707680
rect 490404 707422 490586 707658
rect 490822 707422 491004 707658
rect 490404 707338 491004 707422
rect 490404 707102 490586 707338
rect 490822 707102 491004 707338
rect 486804 705778 487404 705800
rect 486804 705542 486986 705778
rect 487222 705542 487404 705778
rect 486804 705458 487404 705542
rect 486804 705222 486986 705458
rect 487222 705222 487404 705458
rect 486804 701248 487404 705222
rect 486804 701184 486832 701248
rect 486896 701184 486912 701248
rect 486976 701184 486992 701248
rect 487056 701184 487072 701248
rect 487136 701184 487152 701248
rect 487216 701184 487232 701248
rect 487296 701184 487312 701248
rect 487376 701184 487404 701248
rect 486804 700160 487404 701184
rect 486804 700096 486832 700160
rect 486896 700096 486912 700160
rect 486976 700096 486992 700160
rect 487056 700096 487072 700160
rect 487136 700096 487152 700160
rect 487216 700096 487232 700160
rect 487296 700096 487312 700160
rect 487376 700096 487404 700160
rect 486804 699072 487404 700096
rect 486804 699008 486832 699072
rect 486896 699008 486912 699072
rect 486976 699008 486992 699072
rect 487056 699008 487072 699072
rect 487136 699008 487152 699072
rect 487216 699008 487232 699072
rect 487296 699008 487312 699072
rect 487376 699008 487404 699072
rect 486804 697952 487404 699008
rect 490404 698000 491004 707102
rect 494004 698000 494604 708982
rect 497604 698000 498204 710862
rect 515604 710478 516204 711440
rect 515604 710242 515786 710478
rect 516022 710242 516204 710478
rect 515604 710158 516204 710242
rect 515604 709922 515786 710158
rect 516022 709922 516204 710158
rect 512004 708598 512604 709560
rect 512004 708362 512186 708598
rect 512422 708362 512604 708598
rect 512004 708278 512604 708362
rect 512004 708042 512186 708278
rect 512422 708042 512604 708278
rect 508404 706718 509004 707680
rect 508404 706482 508586 706718
rect 508822 706482 509004 706718
rect 508404 706398 509004 706482
rect 508404 706162 508586 706398
rect 508822 706162 509004 706398
rect 504804 704838 505404 705800
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 701792 505404 704282
rect 504804 701728 504832 701792
rect 504896 701728 504912 701792
rect 504976 701728 504992 701792
rect 505056 701728 505072 701792
rect 505136 701728 505152 701792
rect 505216 701728 505232 701792
rect 505296 701728 505312 701792
rect 505376 701728 505404 701792
rect 504804 700704 505404 701728
rect 504804 700640 504832 700704
rect 504896 700640 504912 700704
rect 504976 700640 504992 700704
rect 505056 700640 505072 700704
rect 505136 700640 505152 700704
rect 505216 700640 505232 700704
rect 505296 700640 505312 700704
rect 505376 700640 505404 700704
rect 504804 699616 505404 700640
rect 504804 699552 504832 699616
rect 504896 699552 504912 699616
rect 504976 699552 504992 699616
rect 505056 699552 505072 699616
rect 505136 699552 505152 699616
rect 505216 699552 505232 699616
rect 505296 699552 505312 699616
rect 505376 699552 505404 699616
rect 504804 698528 505404 699552
rect 504804 698464 504832 698528
rect 504896 698464 504912 698528
rect 504976 698464 504992 698528
rect 505056 698464 505072 698528
rect 505136 698464 505152 698528
rect 505216 698464 505232 698528
rect 505296 698464 505312 698528
rect 505376 698464 505404 698528
rect 504804 697952 505404 698464
rect 508404 698000 509004 706162
rect 512004 698000 512604 708042
rect 515604 698000 516204 709922
rect 533604 711418 534204 711440
rect 533604 711182 533786 711418
rect 534022 711182 534204 711418
rect 533604 711098 534204 711182
rect 533604 710862 533786 711098
rect 534022 710862 534204 711098
rect 530004 709538 530604 709560
rect 530004 709302 530186 709538
rect 530422 709302 530604 709538
rect 530004 709218 530604 709302
rect 530004 708982 530186 709218
rect 530422 708982 530604 709218
rect 526404 707658 527004 707680
rect 526404 707422 526586 707658
rect 526822 707422 527004 707658
rect 526404 707338 527004 707422
rect 526404 707102 526586 707338
rect 526822 707102 527004 707338
rect 522804 705778 523404 705800
rect 522804 705542 522986 705778
rect 523222 705542 523404 705778
rect 522804 705458 523404 705542
rect 522804 705222 522986 705458
rect 523222 705222 523404 705458
rect 522804 701248 523404 705222
rect 522804 701184 522832 701248
rect 522896 701184 522912 701248
rect 522976 701184 522992 701248
rect 523056 701184 523072 701248
rect 523136 701184 523152 701248
rect 523216 701184 523232 701248
rect 523296 701184 523312 701248
rect 523376 701184 523404 701248
rect 522804 700160 523404 701184
rect 522804 700096 522832 700160
rect 522896 700096 522912 700160
rect 522976 700096 522992 700160
rect 523056 700096 523072 700160
rect 523136 700096 523152 700160
rect 523216 700096 523232 700160
rect 523296 700096 523312 700160
rect 523376 700096 523404 700160
rect 522804 699072 523404 700096
rect 522804 699008 522832 699072
rect 522896 699008 522912 699072
rect 522976 699008 522992 699072
rect 523056 699008 523072 699072
rect 523136 699008 523152 699072
rect 523216 699008 523232 699072
rect 523296 699008 523312 699072
rect 523376 699008 523404 699072
rect 522804 697952 523404 699008
rect 526404 698000 527004 707102
rect 530004 698000 530604 708982
rect 533604 698000 534204 710862
rect 551604 710478 552204 711440
rect 551604 710242 551786 710478
rect 552022 710242 552204 710478
rect 551604 710158 552204 710242
rect 551604 709922 551786 710158
rect 552022 709922 552204 710158
rect 548004 708598 548604 709560
rect 548004 708362 548186 708598
rect 548422 708362 548604 708598
rect 548004 708278 548604 708362
rect 548004 708042 548186 708278
rect 548422 708042 548604 708278
rect 544404 706718 545004 707680
rect 544404 706482 544586 706718
rect 544822 706482 545004 706718
rect 544404 706398 545004 706482
rect 544404 706162 544586 706398
rect 544822 706162 545004 706398
rect 540804 704838 541404 705800
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 701792 541404 704282
rect 540804 701728 540832 701792
rect 540896 701728 540912 701792
rect 540976 701728 540992 701792
rect 541056 701728 541072 701792
rect 541136 701728 541152 701792
rect 541216 701728 541232 701792
rect 541296 701728 541312 701792
rect 541376 701728 541404 701792
rect 540804 700704 541404 701728
rect 540804 700640 540832 700704
rect 540896 700640 540912 700704
rect 540976 700640 540992 700704
rect 541056 700640 541072 700704
rect 541136 700640 541152 700704
rect 541216 700640 541232 700704
rect 541296 700640 541312 700704
rect 541376 700640 541404 700704
rect 540804 699616 541404 700640
rect 540804 699552 540832 699616
rect 540896 699552 540912 699616
rect 540976 699552 540992 699616
rect 541056 699552 541072 699616
rect 541136 699552 541152 699616
rect 541216 699552 541232 699616
rect 541296 699552 541312 699616
rect 541376 699552 541404 699616
rect 540804 698528 541404 699552
rect 540804 698464 540832 698528
rect 540896 698464 540912 698528
rect 540976 698464 540992 698528
rect 541056 698464 541072 698528
rect 541136 698464 541152 698528
rect 541216 698464 541232 698528
rect 541296 698464 541312 698528
rect 541376 698464 541404 698528
rect 540804 697952 541404 698464
rect 544404 698000 545004 706162
rect 548004 698000 548604 708042
rect 551604 698000 552204 709922
rect 569604 711418 570204 711440
rect 569604 711182 569786 711418
rect 570022 711182 570204 711418
rect 569604 711098 570204 711182
rect 569604 710862 569786 711098
rect 570022 710862 570204 711098
rect 566004 709538 566604 709560
rect 566004 709302 566186 709538
rect 566422 709302 566604 709538
rect 566004 709218 566604 709302
rect 566004 708982 566186 709218
rect 566422 708982 566604 709218
rect 562404 707658 563004 707680
rect 562404 707422 562586 707658
rect 562822 707422 563004 707658
rect 562404 707338 563004 707422
rect 562404 707102 562586 707338
rect 562822 707102 563004 707338
rect 558804 705778 559404 705800
rect 558804 705542 558986 705778
rect 559222 705542 559404 705778
rect 558804 705458 559404 705542
rect 558804 705222 558986 705458
rect 559222 705222 559404 705458
rect 558804 701248 559404 705222
rect 558804 701184 558832 701248
rect 558896 701184 558912 701248
rect 558976 701184 558992 701248
rect 559056 701184 559072 701248
rect 559136 701184 559152 701248
rect 559216 701184 559232 701248
rect 559296 701184 559312 701248
rect 559376 701184 559404 701248
rect 558804 700160 559404 701184
rect 558804 700096 558832 700160
rect 558896 700096 558912 700160
rect 558976 700096 558992 700160
rect 559056 700096 559072 700160
rect 559136 700096 559152 700160
rect 559216 700096 559232 700160
rect 559296 700096 559312 700160
rect 559376 700096 559404 700160
rect 558804 699072 559404 700096
rect 558804 699008 558832 699072
rect 558896 699008 558912 699072
rect 558976 699008 558992 699072
rect 559056 699008 559072 699072
rect 559136 699008 559152 699072
rect 559216 699008 559232 699072
rect 559296 699008 559312 699072
rect 559376 699008 559404 699072
rect 558804 697952 559404 699008
rect 562404 698000 563004 707102
rect 566004 698000 566604 708982
rect 569604 698000 570204 710862
rect 591900 711418 592500 711440
rect 591900 711182 592082 711418
rect 592318 711182 592500 711418
rect 591900 711098 592500 711182
rect 591900 710862 592082 711098
rect 592318 710862 592500 711098
rect 590960 710478 591560 710500
rect 590960 710242 591142 710478
rect 591378 710242 591560 710478
rect 590960 710158 591560 710242
rect 590960 709922 591142 710158
rect 591378 709922 591560 710158
rect 590020 709538 590620 709560
rect 590020 709302 590202 709538
rect 590438 709302 590620 709538
rect 590020 709218 590620 709302
rect 590020 708982 590202 709218
rect 590438 708982 590620 709218
rect 589080 708598 589680 708620
rect 589080 708362 589262 708598
rect 589498 708362 589680 708598
rect 589080 708278 589680 708362
rect 589080 708042 589262 708278
rect 589498 708042 589680 708278
rect 580404 706718 581004 707680
rect 588140 707658 588740 707680
rect 588140 707422 588322 707658
rect 588558 707422 588740 707658
rect 588140 707338 588740 707422
rect 588140 707102 588322 707338
rect 588558 707102 588740 707338
rect 580404 706482 580586 706718
rect 580822 706482 581004 706718
rect 580404 706398 581004 706482
rect 580404 706162 580586 706398
rect 580822 706162 581004 706398
rect 576804 704838 577404 705800
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 701792 577404 704282
rect 576804 701728 576832 701792
rect 576896 701728 576912 701792
rect 576976 701728 576992 701792
rect 577056 701728 577072 701792
rect 577136 701728 577152 701792
rect 577216 701728 577232 701792
rect 577296 701728 577312 701792
rect 577376 701728 577404 701792
rect 576804 700704 577404 701728
rect 576804 700640 576832 700704
rect 576896 700640 576912 700704
rect 576976 700640 576992 700704
rect 577056 700640 577072 700704
rect 577136 700640 577152 700704
rect 577216 700640 577232 700704
rect 577296 700640 577312 700704
rect 577376 700640 577404 700704
rect 576804 699616 577404 700640
rect 576804 699552 576832 699616
rect 576896 699552 576912 699616
rect 576976 699552 576992 699616
rect 577056 699552 577072 699616
rect 577136 699552 577152 699616
rect 577216 699552 577232 699616
rect 577296 699552 577312 699616
rect 577376 699552 577404 699616
rect 576804 698528 577404 699552
rect 576804 698464 576832 698528
rect 576896 698464 576912 698528
rect 576976 698464 576992 698528
rect 577056 698464 577072 698528
rect 577136 698464 577152 698528
rect 577216 698464 577232 698528
rect 577296 698464 577312 698528
rect 577376 698464 577404 698528
rect 576804 697952 577404 698464
rect 521331 695332 521397 695333
rect 521331 695268 521332 695332
rect 521396 695268 521397 695332
rect 521331 695267 521397 695268
rect 500907 694924 500973 694925
rect 500907 694860 500908 694924
rect 500972 694860 500973 694924
rect 500907 694859 500973 694860
rect 505691 694924 505757 694925
rect 505691 694860 505692 694924
rect 505756 694860 505757 694924
rect 505691 694859 505757 694860
rect 500910 694653 500970 694859
rect 492811 694652 492877 694653
rect 492811 694588 492812 694652
rect 492876 694588 492877 694652
rect 492811 694587 492877 694588
rect 500907 694652 500973 694653
rect 500907 694588 500908 694652
rect 500972 694588 500973 694652
rect 500907 694587 500973 694588
rect 446995 694516 447061 694517
rect 446995 694452 446996 694516
rect 447060 694452 447061 694516
rect 446995 694451 447061 694452
rect 447179 694516 447245 694517
rect 447179 694452 447180 694516
rect 447244 694452 447245 694516
rect 447179 694451 447245 694452
rect 476067 694516 476133 694517
rect 476067 694452 476068 694516
rect 476132 694452 476133 694516
rect 476067 694451 476133 694452
rect 439451 694380 439517 694381
rect 439451 694316 439452 694380
rect 439516 694316 439517 694380
rect 439451 694315 439517 694316
rect 446998 694109 447058 694451
rect 451227 694380 451293 694381
rect 451227 694316 451228 694380
rect 451292 694316 451293 694380
rect 451227 694315 451293 694316
rect 475883 694380 475949 694381
rect 475883 694316 475884 694380
rect 475948 694316 475949 694380
rect 475883 694315 475949 694316
rect 417739 694108 417805 694109
rect 417739 694044 417740 694108
rect 417804 694044 417805 694108
rect 417739 694043 417805 694044
rect 427675 694108 427741 694109
rect 427675 694044 427676 694108
rect 427740 694044 427741 694108
rect 427675 694043 427741 694044
rect 427859 694108 427925 694109
rect 427859 694044 427860 694108
rect 427924 694044 427925 694108
rect 427859 694043 427925 694044
rect 437243 694108 437309 694109
rect 437243 694044 437244 694108
rect 437308 694044 437309 694108
rect 437243 694043 437309 694044
rect 437427 694108 437493 694109
rect 437427 694044 437428 694108
rect 437492 694044 437493 694108
rect 437427 694043 437493 694044
rect 446995 694108 447061 694109
rect 446995 694044 446996 694108
rect 447060 694044 447061 694108
rect 446995 694043 447061 694044
rect 415163 693972 415229 693973
rect 415163 693970 415164 693972
rect 414982 693910 415164 693970
rect 410563 693907 410629 693908
rect 415163 693908 415164 693910
rect 415228 693908 415229 693972
rect 451230 693970 451290 694315
rect 475886 694109 475946 694315
rect 476070 694245 476130 694451
rect 476067 694244 476133 694245
rect 476067 694180 476068 694244
rect 476132 694180 476133 694244
rect 476067 694179 476133 694180
rect 492627 694244 492693 694245
rect 492627 694180 492628 694244
rect 492692 694242 492693 694244
rect 492814 694242 492874 694587
rect 505694 694381 505754 694859
rect 505691 694380 505757 694381
rect 505691 694316 505692 694380
rect 505756 694316 505757 694380
rect 505691 694315 505757 694316
rect 492692 694182 492874 694242
rect 492692 694180 492693 694182
rect 492627 694179 492693 694180
rect 451411 694108 451477 694109
rect 451411 694044 451412 694108
rect 451476 694044 451477 694108
rect 451411 694043 451477 694044
rect 475883 694108 475949 694109
rect 475883 694044 475884 694108
rect 475948 694044 475949 694108
rect 475883 694043 475949 694044
rect 451414 693970 451474 694043
rect 451230 693910 451474 693970
rect 415163 693907 415229 693908
rect 521334 693701 521394 695267
rect 531267 694652 531333 694653
rect 531267 694588 531268 694652
rect 531332 694588 531333 694652
rect 531267 694587 531333 694588
rect 562918 694590 563162 694650
rect 521699 694516 521765 694517
rect 521699 694452 521700 694516
rect 521764 694452 521765 694516
rect 521699 694451 521765 694452
rect 521702 694245 521762 694451
rect 531270 694245 531330 694587
rect 562918 694381 562978 694590
rect 543595 694380 543661 694381
rect 543595 694316 543596 694380
rect 543660 694316 543661 694380
rect 543595 694315 543661 694316
rect 562915 694380 562981 694381
rect 562915 694316 562916 694380
rect 562980 694316 562981 694380
rect 562915 694315 562981 694316
rect 521699 694244 521765 694245
rect 521699 694180 521700 694244
rect 521764 694180 521765 694244
rect 521699 694179 521765 694180
rect 531267 694244 531333 694245
rect 531267 694180 531268 694244
rect 531332 694180 531333 694244
rect 531267 694179 531333 694180
rect 529243 694108 529309 694109
rect 529243 694044 529244 694108
rect 529308 694044 529309 694108
rect 529243 694043 529309 694044
rect 538811 694108 538877 694109
rect 538811 694044 538812 694108
rect 538876 694044 538877 694108
rect 543598 694106 543658 694315
rect 563102 694245 563162 694590
rect 568619 694380 568685 694381
rect 568619 694316 568620 694380
rect 568684 694316 568685 694380
rect 568619 694315 568685 694316
rect 568622 694245 568682 694315
rect 543779 694244 543845 694245
rect 543779 694180 543780 694244
rect 543844 694180 543845 694244
rect 543779 694179 543845 694180
rect 563099 694244 563165 694245
rect 563099 694180 563100 694244
rect 563164 694180 563165 694244
rect 563099 694179 563165 694180
rect 568619 694244 568685 694245
rect 568619 694180 568620 694244
rect 568684 694180 568685 694244
rect 568619 694179 568685 694180
rect 543782 694106 543842 694179
rect 543598 694046 543842 694106
rect 548563 694108 548629 694109
rect 538811 694043 538877 694044
rect 548563 694044 548564 694108
rect 548628 694044 548629 694108
rect 548563 694043 548629 694044
rect 529246 693701 529306 694043
rect 538814 693701 538874 694043
rect 548566 693701 548626 694043
rect 255267 693700 255333 693701
rect 255267 693636 255268 693700
rect 255332 693636 255333 693700
rect 255267 693635 255333 693636
rect 270907 693700 270973 693701
rect 270907 693636 270908 693700
rect 270972 693636 270973 693700
rect 270907 693635 270973 693636
rect 271275 693700 271341 693701
rect 271275 693636 271276 693700
rect 271340 693636 271341 693700
rect 271275 693635 271341 693636
rect 414427 693700 414493 693701
rect 414427 693636 414428 693700
rect 414492 693636 414493 693700
rect 414427 693635 414493 693636
rect 415163 693700 415229 693701
rect 415163 693636 415164 693700
rect 415228 693636 415229 693700
rect 415163 693635 415229 693636
rect 521331 693700 521397 693701
rect 521331 693636 521332 693700
rect 521396 693636 521397 693700
rect 521331 693635 521397 693636
rect 529243 693700 529309 693701
rect 529243 693636 529244 693700
rect 529308 693636 529309 693700
rect 529243 693635 529309 693636
rect 538811 693700 538877 693701
rect 538811 693636 538812 693700
rect 538876 693636 538877 693700
rect 538811 693635 538877 693636
rect 548563 693700 548629 693701
rect 548563 693636 548564 693700
rect 548628 693636 548629 693700
rect 548563 693635 548629 693636
rect 251222 692550 252018 692610
rect 414430 692610 414490 693635
rect 415166 692610 415226 693635
rect 414430 692550 415226 692610
rect 4404 689818 4586 690054
rect 4822 689818 5004 690054
rect 4404 689734 5004 689818
rect 4404 689498 4586 689734
rect 4822 689498 5004 689734
rect 4404 654054 5004 689498
rect 4404 653818 4586 654054
rect 4822 653818 5004 654054
rect 4404 653734 5004 653818
rect 4404 653498 4586 653734
rect 4822 653498 5004 653734
rect 4404 618054 5004 653498
rect 4404 617818 4586 618054
rect 4822 617818 5004 618054
rect 4404 617734 5004 617818
rect 4404 617498 4586 617734
rect 4822 617498 5004 617734
rect 4404 582054 5004 617498
rect 4404 581818 4586 582054
rect 4822 581818 5004 582054
rect 4404 581734 5004 581818
rect 4404 581498 4586 581734
rect 4822 581498 5004 581734
rect 4404 546054 5004 581498
rect 4404 545818 4586 546054
rect 4822 545818 5004 546054
rect 4404 545734 5004 545818
rect 4404 545498 4586 545734
rect 4822 545498 5004 545734
rect 4404 510054 5004 545498
rect 4404 509818 4586 510054
rect 4822 509818 5004 510054
rect 4404 509734 5004 509818
rect 4404 509498 4586 509734
rect 4822 509498 5004 509734
rect 4404 474054 5004 509498
rect 4404 473818 4586 474054
rect 4822 473818 5004 474054
rect 4404 473734 5004 473818
rect 4404 473498 4586 473734
rect 4822 473498 5004 473734
rect 4404 438054 5004 473498
rect 4404 437818 4586 438054
rect 4822 437818 5004 438054
rect 4404 437734 5004 437818
rect 4404 437498 4586 437734
rect 4822 437498 5004 437734
rect 4404 402054 5004 437498
rect 4404 401818 4586 402054
rect 4822 401818 5004 402054
rect 4404 401734 5004 401818
rect 4404 401498 4586 401734
rect 4822 401498 5004 401734
rect 4404 366054 5004 401498
rect 4404 365818 4586 366054
rect 4822 365818 5004 366054
rect 4404 365734 5004 365818
rect 4404 365498 4586 365734
rect 4822 365498 5004 365734
rect 4404 330054 5004 365498
rect 4404 329818 4586 330054
rect 4822 329818 5004 330054
rect 4404 329734 5004 329818
rect 4404 329498 4586 329734
rect 4822 329498 5004 329734
rect 4404 294054 5004 329498
rect 4404 293818 4586 294054
rect 4822 293818 5004 294054
rect 4404 293734 5004 293818
rect 4404 293498 4586 293734
rect 4822 293498 5004 293734
rect 4404 258054 5004 293498
rect 4404 257818 4586 258054
rect 4822 257818 5004 258054
rect 4404 257734 5004 257818
rect 4404 257498 4586 257734
rect 4822 257498 5004 257734
rect 4404 222054 5004 257498
rect 4404 221818 4586 222054
rect 4822 221818 5004 222054
rect 4404 221734 5004 221818
rect 4404 221498 4586 221734
rect 4822 221498 5004 221734
rect 4404 186054 5004 221498
rect 4404 185818 4586 186054
rect 4822 185818 5004 186054
rect 4404 185734 5004 185818
rect 4404 185498 4586 185734
rect 4822 185498 5004 185734
rect 4404 150054 5004 185498
rect 4404 149818 4586 150054
rect 4822 149818 5004 150054
rect 4404 149734 5004 149818
rect 4404 149498 4586 149734
rect 4822 149498 5004 149734
rect 4404 114054 5004 149498
rect 4404 113818 4586 114054
rect 4822 113818 5004 114054
rect 4404 113734 5004 113818
rect 4404 113498 4586 113734
rect 4822 113498 5004 113734
rect 4404 78054 5004 113498
rect 4404 77818 4586 78054
rect 4822 77818 5004 78054
rect 4404 77734 5004 77818
rect 4404 77498 4586 77734
rect 4822 77498 5004 77734
rect 4404 42054 5004 77498
rect 4404 41818 4586 42054
rect 4822 41818 5004 42054
rect 4404 41734 5004 41818
rect 4404 41498 4586 41734
rect 4822 41498 5004 41734
rect 4404 6054 5004 41498
rect 4404 5818 4586 6054
rect 4822 5818 5004 6054
rect 580404 690054 581004 706162
rect 587200 706718 587800 706740
rect 587200 706482 587382 706718
rect 587618 706482 587800 706718
rect 587200 706398 587800 706482
rect 587200 706162 587382 706398
rect 587618 706162 587800 706398
rect 586260 705778 586860 705800
rect 586260 705542 586442 705778
rect 586678 705542 586860 705778
rect 586260 705458 586860 705542
rect 586260 705222 586442 705458
rect 586678 705222 586860 705458
rect 580404 689818 580586 690054
rect 580822 689818 581004 690054
rect 580404 689734 581004 689818
rect 580404 689498 580586 689734
rect 580822 689498 581004 689734
rect 580404 654054 581004 689498
rect 580404 653818 580586 654054
rect 580822 653818 581004 654054
rect 580404 653734 581004 653818
rect 580404 653498 580586 653734
rect 580822 653498 581004 653734
rect 580404 618054 581004 653498
rect 580404 617818 580586 618054
rect 580822 617818 581004 618054
rect 580404 617734 581004 617818
rect 580404 617498 580586 617734
rect 580822 617498 581004 617734
rect 580404 582054 581004 617498
rect 580404 581818 580586 582054
rect 580822 581818 581004 582054
rect 580404 581734 581004 581818
rect 580404 581498 580586 581734
rect 580822 581498 581004 581734
rect 580404 546054 581004 581498
rect 580404 545818 580586 546054
rect 580822 545818 581004 546054
rect 580404 545734 581004 545818
rect 580404 545498 580586 545734
rect 580822 545498 581004 545734
rect 580404 510054 581004 545498
rect 580404 509818 580586 510054
rect 580822 509818 581004 510054
rect 580404 509734 581004 509818
rect 580404 509498 580586 509734
rect 580822 509498 581004 509734
rect 580404 474054 581004 509498
rect 580404 473818 580586 474054
rect 580822 473818 581004 474054
rect 580404 473734 581004 473818
rect 580404 473498 580586 473734
rect 580822 473498 581004 473734
rect 580404 438054 581004 473498
rect 580404 437818 580586 438054
rect 580822 437818 581004 438054
rect 580404 437734 581004 437818
rect 580404 437498 580586 437734
rect 580822 437498 581004 437734
rect 580404 402054 581004 437498
rect 580404 401818 580586 402054
rect 580822 401818 581004 402054
rect 580404 401734 581004 401818
rect 580404 401498 580586 401734
rect 580822 401498 581004 401734
rect 580404 366054 581004 401498
rect 580404 365818 580586 366054
rect 580822 365818 581004 366054
rect 580404 365734 581004 365818
rect 580404 365498 580586 365734
rect 580822 365498 581004 365734
rect 580404 330054 581004 365498
rect 580404 329818 580586 330054
rect 580822 329818 581004 330054
rect 580404 329734 581004 329818
rect 580404 329498 580586 329734
rect 580822 329498 581004 329734
rect 580404 294054 581004 329498
rect 580404 293818 580586 294054
rect 580822 293818 581004 294054
rect 580404 293734 581004 293818
rect 580404 293498 580586 293734
rect 580822 293498 581004 293734
rect 580404 258054 581004 293498
rect 580404 257818 580586 258054
rect 580822 257818 581004 258054
rect 580404 257734 581004 257818
rect 580404 257498 580586 257734
rect 580822 257498 581004 257734
rect 580404 222054 581004 257498
rect 580404 221818 580586 222054
rect 580822 221818 581004 222054
rect 580404 221734 581004 221818
rect 580404 221498 580586 221734
rect 580822 221498 581004 221734
rect 580404 186054 581004 221498
rect 580404 185818 580586 186054
rect 580822 185818 581004 186054
rect 580404 185734 581004 185818
rect 580404 185498 580586 185734
rect 580822 185498 581004 185734
rect 580404 150054 581004 185498
rect 580404 149818 580586 150054
rect 580822 149818 581004 150054
rect 580404 149734 581004 149818
rect 580404 149498 580586 149734
rect 580822 149498 581004 149734
rect 580404 114054 581004 149498
rect 580404 113818 580586 114054
rect 580822 113818 581004 114054
rect 580404 113734 581004 113818
rect 580404 113498 580586 113734
rect 580822 113498 581004 113734
rect 580404 78054 581004 113498
rect 580404 77818 580586 78054
rect 580822 77818 581004 78054
rect 580404 77734 581004 77818
rect 580404 77498 580586 77734
rect 580822 77498 581004 77734
rect 580404 42054 581004 77498
rect 580404 41818 580586 42054
rect 580822 41818 581004 42054
rect 580404 41734 581004 41818
rect 580404 41498 580586 41734
rect 580822 41498 581004 41734
rect 580404 6054 581004 41498
rect 18804 6016 19404 6048
rect 4404 5734 5004 5818
rect 4404 5498 4586 5734
rect 4822 5498 5004 5734
rect -3876 -2462 -3694 -2226
rect -3458 -2462 -3276 -2226
rect -3876 -2546 -3276 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 -3276 -2546
rect -3876 -2804 -3276 -2782
rect 4404 -2226 5004 5498
rect 4404 -2462 4586 -2226
rect 4822 -2462 5004 -2226
rect 4404 -2546 5004 -2462
rect 4404 -2782 4586 -2546
rect 4822 -2782 5004 -2546
rect -4816 -3402 -4634 -3166
rect -4398 -3402 -4216 -3166
rect -4816 -3486 -4216 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 -4216 -3486
rect -4816 -3744 -4216 -3722
rect 4404 -3744 5004 -2782
rect -5756 -4342 -5574 -4106
rect -5338 -4342 -5156 -4106
rect -5756 -4426 -5156 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 -5156 -4426
rect -5756 -4684 -5156 -4662
rect 8004 -4106 8604 6000
rect 8004 -4342 8186 -4106
rect 8422 -4342 8604 -4106
rect 8004 -4426 8604 -4342
rect 8004 -4662 8186 -4426
rect 8422 -4662 8604 -4426
rect -6696 -5282 -6514 -5046
rect -6278 -5282 -6096 -5046
rect -6696 -5366 -6096 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 -6096 -5366
rect -6696 -5624 -6096 -5602
rect 8004 -5624 8604 -4662
rect -7636 -6222 -7454 -5986
rect -7218 -6222 -7036 -5986
rect -7636 -6306 -7036 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 -7036 -6306
rect -7636 -6564 -7036 -6542
rect 11604 -5986 12204 6000
rect 18804 5952 18832 6016
rect 18896 5952 18912 6016
rect 18976 5952 18992 6016
rect 19056 5952 19072 6016
rect 19136 5952 19152 6016
rect 19216 5952 19232 6016
rect 19296 5952 19312 6016
rect 19376 5952 19404 6016
rect 18804 4928 19404 5952
rect 18804 4864 18832 4928
rect 18896 4864 18912 4928
rect 18976 4864 18992 4928
rect 19056 4864 19072 4928
rect 19136 4864 19152 4928
rect 19216 4864 19232 4928
rect 19296 4864 19312 4928
rect 19376 4864 19404 4928
rect 18804 3840 19404 4864
rect 18804 3776 18832 3840
rect 18896 3776 18912 3840
rect 18976 3776 18992 3840
rect 19056 3776 19072 3840
rect 19136 3776 19152 3840
rect 19216 3776 19232 3840
rect 19296 3776 19312 3840
rect 19376 3776 19404 3840
rect 18804 2752 19404 3776
rect 18804 2688 18832 2752
rect 18896 2688 18912 2752
rect 18976 2688 18992 2752
rect 19056 2688 19072 2752
rect 19136 2688 19152 2752
rect 19216 2688 19232 2752
rect 19296 2688 19312 2752
rect 19376 2688 19404 2752
rect 18804 -1286 19404 2688
rect 18804 -1522 18986 -1286
rect 19222 -1522 19404 -1286
rect 18804 -1606 19404 -1522
rect 18804 -1842 18986 -1606
rect 19222 -1842 19404 -1606
rect 18804 -1864 19404 -1842
rect 22404 -3166 23004 6000
rect 22404 -3402 22586 -3166
rect 22822 -3402 23004 -3166
rect 22404 -3486 23004 -3402
rect 22404 -3722 22586 -3486
rect 22822 -3722 23004 -3486
rect 22404 -3744 23004 -3722
rect 26004 -5046 26604 6000
rect 26004 -5282 26186 -5046
rect 26422 -5282 26604 -5046
rect 26004 -5366 26604 -5282
rect 26004 -5602 26186 -5366
rect 26422 -5602 26604 -5366
rect 26004 -5624 26604 -5602
rect 11604 -6222 11786 -5986
rect 12022 -6222 12204 -5986
rect 11604 -6306 12204 -6222
rect 11604 -6542 11786 -6306
rect 12022 -6542 12204 -6306
rect -8576 -7162 -8394 -6926
rect -8158 -7162 -7976 -6926
rect -8576 -7246 -7976 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 -7976 -7246
rect -8576 -7504 -7976 -7482
rect 11604 -7504 12204 -6542
rect 29604 -6926 30204 6000
rect 36804 5472 37404 6048
rect 54804 6016 55404 6048
rect 36804 5408 36832 5472
rect 36896 5408 36912 5472
rect 36976 5408 36992 5472
rect 37056 5408 37072 5472
rect 37136 5408 37152 5472
rect 37216 5408 37232 5472
rect 37296 5408 37312 5472
rect 37376 5408 37404 5472
rect 36804 4384 37404 5408
rect 36804 4320 36832 4384
rect 36896 4320 36912 4384
rect 36976 4320 36992 4384
rect 37056 4320 37072 4384
rect 37136 4320 37152 4384
rect 37216 4320 37232 4384
rect 37296 4320 37312 4384
rect 37376 4320 37404 4384
rect 36804 3296 37404 4320
rect 36804 3232 36832 3296
rect 36896 3232 36912 3296
rect 36976 3232 36992 3296
rect 37056 3232 37072 3296
rect 37136 3232 37152 3296
rect 37216 3232 37232 3296
rect 37296 3232 37312 3296
rect 37376 3232 37404 3296
rect 36804 2406 37404 3232
rect 36804 2208 36986 2406
rect 37222 2208 37404 2406
rect 36804 2144 36832 2208
rect 36896 2144 36912 2208
rect 36976 2170 36986 2208
rect 37222 2170 37232 2208
rect 36976 2144 36992 2170
rect 37056 2144 37072 2170
rect 37136 2144 37152 2170
rect 37216 2144 37232 2170
rect 37296 2144 37312 2208
rect 37376 2144 37404 2208
rect 36804 2086 37404 2144
rect 36804 1850 36986 2086
rect 37222 1850 37404 2086
rect 36804 -346 37404 1850
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1864 37404 -902
rect 40404 -2226 41004 6000
rect 40404 -2462 40586 -2226
rect 40822 -2462 41004 -2226
rect 40404 -2546 41004 -2462
rect 40404 -2782 40586 -2546
rect 40822 -2782 41004 -2546
rect 40404 -3744 41004 -2782
rect 44004 -4106 44604 6000
rect 44004 -4342 44186 -4106
rect 44422 -4342 44604 -4106
rect 44004 -4426 44604 -4342
rect 44004 -4662 44186 -4426
rect 44422 -4662 44604 -4426
rect 44004 -5624 44604 -4662
rect 29604 -7162 29786 -6926
rect 30022 -7162 30204 -6926
rect 29604 -7246 30204 -7162
rect 29604 -7482 29786 -7246
rect 30022 -7482 30204 -7246
rect 29604 -7504 30204 -7482
rect 47604 -5986 48204 6000
rect 54804 5952 54832 6016
rect 54896 5952 54912 6016
rect 54976 5952 54992 6016
rect 55056 5952 55072 6016
rect 55136 5952 55152 6016
rect 55216 5952 55232 6016
rect 55296 5952 55312 6016
rect 55376 5952 55404 6016
rect 54804 4928 55404 5952
rect 54804 4864 54832 4928
rect 54896 4864 54912 4928
rect 54976 4864 54992 4928
rect 55056 4864 55072 4928
rect 55136 4864 55152 4928
rect 55216 4864 55232 4928
rect 55296 4864 55312 4928
rect 55376 4864 55404 4928
rect 54804 3840 55404 4864
rect 54804 3776 54832 3840
rect 54896 3776 54912 3840
rect 54976 3776 54992 3840
rect 55056 3776 55072 3840
rect 55136 3776 55152 3840
rect 55216 3776 55232 3840
rect 55296 3776 55312 3840
rect 55376 3776 55404 3840
rect 54804 2752 55404 3776
rect 54804 2688 54832 2752
rect 54896 2688 54912 2752
rect 54976 2688 54992 2752
rect 55056 2688 55072 2752
rect 55136 2688 55152 2752
rect 55216 2688 55232 2752
rect 55296 2688 55312 2752
rect 55376 2688 55404 2752
rect 54804 -1286 55404 2688
rect 54804 -1522 54986 -1286
rect 55222 -1522 55404 -1286
rect 54804 -1606 55404 -1522
rect 54804 -1842 54986 -1606
rect 55222 -1842 55404 -1606
rect 54804 -1864 55404 -1842
rect 58404 -3166 59004 6000
rect 58404 -3402 58586 -3166
rect 58822 -3402 59004 -3166
rect 58404 -3486 59004 -3402
rect 58404 -3722 58586 -3486
rect 58822 -3722 59004 -3486
rect 58404 -3744 59004 -3722
rect 62004 -5046 62604 6000
rect 62004 -5282 62186 -5046
rect 62422 -5282 62604 -5046
rect 62004 -5366 62604 -5282
rect 62004 -5602 62186 -5366
rect 62422 -5602 62604 -5366
rect 62004 -5624 62604 -5602
rect 47604 -6222 47786 -5986
rect 48022 -6222 48204 -5986
rect 47604 -6306 48204 -6222
rect 47604 -6542 47786 -6306
rect 48022 -6542 48204 -6306
rect 47604 -7504 48204 -6542
rect 65604 -6926 66204 6000
rect 72804 5472 73404 6048
rect 90804 6016 91404 6048
rect 72804 5408 72832 5472
rect 72896 5408 72912 5472
rect 72976 5408 72992 5472
rect 73056 5408 73072 5472
rect 73136 5408 73152 5472
rect 73216 5408 73232 5472
rect 73296 5408 73312 5472
rect 73376 5408 73404 5472
rect 72804 4384 73404 5408
rect 72804 4320 72832 4384
rect 72896 4320 72912 4384
rect 72976 4320 72992 4384
rect 73056 4320 73072 4384
rect 73136 4320 73152 4384
rect 73216 4320 73232 4384
rect 73296 4320 73312 4384
rect 73376 4320 73404 4384
rect 72804 3296 73404 4320
rect 72804 3232 72832 3296
rect 72896 3232 72912 3296
rect 72976 3232 72992 3296
rect 73056 3232 73072 3296
rect 73136 3232 73152 3296
rect 73216 3232 73232 3296
rect 73296 3232 73312 3296
rect 73376 3232 73404 3296
rect 72804 2406 73404 3232
rect 72804 2208 72986 2406
rect 73222 2208 73404 2406
rect 72804 2144 72832 2208
rect 72896 2144 72912 2208
rect 72976 2170 72986 2208
rect 73222 2170 73232 2208
rect 72976 2144 72992 2170
rect 73056 2144 73072 2170
rect 73136 2144 73152 2170
rect 73216 2144 73232 2170
rect 73296 2144 73312 2208
rect 73376 2144 73404 2208
rect 72804 2086 73404 2144
rect 72804 1850 72986 2086
rect 73222 1850 73404 2086
rect 72804 -346 73404 1850
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1864 73404 -902
rect 76404 -2226 77004 6000
rect 76404 -2462 76586 -2226
rect 76822 -2462 77004 -2226
rect 76404 -2546 77004 -2462
rect 76404 -2782 76586 -2546
rect 76822 -2782 77004 -2546
rect 76404 -3744 77004 -2782
rect 80004 -4106 80604 6000
rect 80004 -4342 80186 -4106
rect 80422 -4342 80604 -4106
rect 80004 -4426 80604 -4342
rect 80004 -4662 80186 -4426
rect 80422 -4662 80604 -4426
rect 80004 -5624 80604 -4662
rect 65604 -7162 65786 -6926
rect 66022 -7162 66204 -6926
rect 65604 -7246 66204 -7162
rect 65604 -7482 65786 -7246
rect 66022 -7482 66204 -7246
rect 65604 -7504 66204 -7482
rect 83604 -5986 84204 6000
rect 90804 5952 90832 6016
rect 90896 5952 90912 6016
rect 90976 5952 90992 6016
rect 91056 5952 91072 6016
rect 91136 5952 91152 6016
rect 91216 5952 91232 6016
rect 91296 5952 91312 6016
rect 91376 5952 91404 6016
rect 90804 4928 91404 5952
rect 90804 4864 90832 4928
rect 90896 4864 90912 4928
rect 90976 4864 90992 4928
rect 91056 4864 91072 4928
rect 91136 4864 91152 4928
rect 91216 4864 91232 4928
rect 91296 4864 91312 4928
rect 91376 4864 91404 4928
rect 90804 3840 91404 4864
rect 90804 3776 90832 3840
rect 90896 3776 90912 3840
rect 90976 3776 90992 3840
rect 91056 3776 91072 3840
rect 91136 3776 91152 3840
rect 91216 3776 91232 3840
rect 91296 3776 91312 3840
rect 91376 3776 91404 3840
rect 90804 2752 91404 3776
rect 90804 2688 90832 2752
rect 90896 2688 90912 2752
rect 90976 2688 90992 2752
rect 91056 2688 91072 2752
rect 91136 2688 91152 2752
rect 91216 2688 91232 2752
rect 91296 2688 91312 2752
rect 91376 2688 91404 2752
rect 90804 -1286 91404 2688
rect 90804 -1522 90986 -1286
rect 91222 -1522 91404 -1286
rect 90804 -1606 91404 -1522
rect 90804 -1842 90986 -1606
rect 91222 -1842 91404 -1606
rect 90804 -1864 91404 -1842
rect 94404 -3166 95004 6000
rect 94404 -3402 94586 -3166
rect 94822 -3402 95004 -3166
rect 94404 -3486 95004 -3402
rect 94404 -3722 94586 -3486
rect 94822 -3722 95004 -3486
rect 94404 -3744 95004 -3722
rect 98004 -5046 98604 6000
rect 98004 -5282 98186 -5046
rect 98422 -5282 98604 -5046
rect 98004 -5366 98604 -5282
rect 98004 -5602 98186 -5366
rect 98422 -5602 98604 -5366
rect 98004 -5624 98604 -5602
rect 83604 -6222 83786 -5986
rect 84022 -6222 84204 -5986
rect 83604 -6306 84204 -6222
rect 83604 -6542 83786 -6306
rect 84022 -6542 84204 -6306
rect 83604 -7504 84204 -6542
rect 101604 -6926 102204 6000
rect 108804 5472 109404 6048
rect 126804 6016 127404 6048
rect 108804 5408 108832 5472
rect 108896 5408 108912 5472
rect 108976 5408 108992 5472
rect 109056 5408 109072 5472
rect 109136 5408 109152 5472
rect 109216 5408 109232 5472
rect 109296 5408 109312 5472
rect 109376 5408 109404 5472
rect 108804 4384 109404 5408
rect 108804 4320 108832 4384
rect 108896 4320 108912 4384
rect 108976 4320 108992 4384
rect 109056 4320 109072 4384
rect 109136 4320 109152 4384
rect 109216 4320 109232 4384
rect 109296 4320 109312 4384
rect 109376 4320 109404 4384
rect 108804 3296 109404 4320
rect 108804 3232 108832 3296
rect 108896 3232 108912 3296
rect 108976 3232 108992 3296
rect 109056 3232 109072 3296
rect 109136 3232 109152 3296
rect 109216 3232 109232 3296
rect 109296 3232 109312 3296
rect 109376 3232 109404 3296
rect 108804 2406 109404 3232
rect 108804 2208 108986 2406
rect 109222 2208 109404 2406
rect 108804 2144 108832 2208
rect 108896 2144 108912 2208
rect 108976 2170 108986 2208
rect 109222 2170 109232 2208
rect 108976 2144 108992 2170
rect 109056 2144 109072 2170
rect 109136 2144 109152 2170
rect 109216 2144 109232 2170
rect 109296 2144 109312 2208
rect 109376 2144 109404 2208
rect 108804 2086 109404 2144
rect 108804 1850 108986 2086
rect 109222 1850 109404 2086
rect 108804 -346 109404 1850
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1864 109404 -902
rect 112404 -2226 113004 6000
rect 112404 -2462 112586 -2226
rect 112822 -2462 113004 -2226
rect 112404 -2546 113004 -2462
rect 112404 -2782 112586 -2546
rect 112822 -2782 113004 -2546
rect 112404 -3744 113004 -2782
rect 116004 -4106 116604 6000
rect 116004 -4342 116186 -4106
rect 116422 -4342 116604 -4106
rect 116004 -4426 116604 -4342
rect 116004 -4662 116186 -4426
rect 116422 -4662 116604 -4426
rect 116004 -5624 116604 -4662
rect 101604 -7162 101786 -6926
rect 102022 -7162 102204 -6926
rect 101604 -7246 102204 -7162
rect 101604 -7482 101786 -7246
rect 102022 -7482 102204 -7246
rect 101604 -7504 102204 -7482
rect 119604 -5986 120204 6000
rect 126804 5952 126832 6016
rect 126896 5952 126912 6016
rect 126976 5952 126992 6016
rect 127056 5952 127072 6016
rect 127136 5952 127152 6016
rect 127216 5952 127232 6016
rect 127296 5952 127312 6016
rect 127376 5952 127404 6016
rect 126804 4928 127404 5952
rect 126804 4864 126832 4928
rect 126896 4864 126912 4928
rect 126976 4864 126992 4928
rect 127056 4864 127072 4928
rect 127136 4864 127152 4928
rect 127216 4864 127232 4928
rect 127296 4864 127312 4928
rect 127376 4864 127404 4928
rect 126804 3840 127404 4864
rect 126804 3776 126832 3840
rect 126896 3776 126912 3840
rect 126976 3776 126992 3840
rect 127056 3776 127072 3840
rect 127136 3776 127152 3840
rect 127216 3776 127232 3840
rect 127296 3776 127312 3840
rect 127376 3776 127404 3840
rect 126804 2752 127404 3776
rect 126804 2688 126832 2752
rect 126896 2688 126912 2752
rect 126976 2688 126992 2752
rect 127056 2688 127072 2752
rect 127136 2688 127152 2752
rect 127216 2688 127232 2752
rect 127296 2688 127312 2752
rect 127376 2688 127404 2752
rect 126804 -1286 127404 2688
rect 126804 -1522 126986 -1286
rect 127222 -1522 127404 -1286
rect 126804 -1606 127404 -1522
rect 126804 -1842 126986 -1606
rect 127222 -1842 127404 -1606
rect 126804 -1864 127404 -1842
rect 130404 -3166 131004 6000
rect 130404 -3402 130586 -3166
rect 130822 -3402 131004 -3166
rect 130404 -3486 131004 -3402
rect 130404 -3722 130586 -3486
rect 130822 -3722 131004 -3486
rect 130404 -3744 131004 -3722
rect 134004 -5046 134604 6000
rect 134004 -5282 134186 -5046
rect 134422 -5282 134604 -5046
rect 134004 -5366 134604 -5282
rect 134004 -5602 134186 -5366
rect 134422 -5602 134604 -5366
rect 134004 -5624 134604 -5602
rect 119604 -6222 119786 -5986
rect 120022 -6222 120204 -5986
rect 119604 -6306 120204 -6222
rect 119604 -6542 119786 -6306
rect 120022 -6542 120204 -6306
rect 119604 -7504 120204 -6542
rect 137604 -6926 138204 6000
rect 144804 5472 145404 6048
rect 162804 6016 163404 6048
rect 144804 5408 144832 5472
rect 144896 5408 144912 5472
rect 144976 5408 144992 5472
rect 145056 5408 145072 5472
rect 145136 5408 145152 5472
rect 145216 5408 145232 5472
rect 145296 5408 145312 5472
rect 145376 5408 145404 5472
rect 144804 4384 145404 5408
rect 144804 4320 144832 4384
rect 144896 4320 144912 4384
rect 144976 4320 144992 4384
rect 145056 4320 145072 4384
rect 145136 4320 145152 4384
rect 145216 4320 145232 4384
rect 145296 4320 145312 4384
rect 145376 4320 145404 4384
rect 144804 3296 145404 4320
rect 144804 3232 144832 3296
rect 144896 3232 144912 3296
rect 144976 3232 144992 3296
rect 145056 3232 145072 3296
rect 145136 3232 145152 3296
rect 145216 3232 145232 3296
rect 145296 3232 145312 3296
rect 145376 3232 145404 3296
rect 144804 2406 145404 3232
rect 144804 2208 144986 2406
rect 145222 2208 145404 2406
rect 144804 2144 144832 2208
rect 144896 2144 144912 2208
rect 144976 2170 144986 2208
rect 145222 2170 145232 2208
rect 144976 2144 144992 2170
rect 145056 2144 145072 2170
rect 145136 2144 145152 2170
rect 145216 2144 145232 2170
rect 145296 2144 145312 2208
rect 145376 2144 145404 2208
rect 144804 2086 145404 2144
rect 144804 1850 144986 2086
rect 145222 1850 145404 2086
rect 144804 -346 145404 1850
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1864 145404 -902
rect 148404 -2226 149004 6000
rect 148404 -2462 148586 -2226
rect 148822 -2462 149004 -2226
rect 148404 -2546 149004 -2462
rect 148404 -2782 148586 -2546
rect 148822 -2782 149004 -2546
rect 148404 -3744 149004 -2782
rect 152004 -4106 152604 6000
rect 152004 -4342 152186 -4106
rect 152422 -4342 152604 -4106
rect 152004 -4426 152604 -4342
rect 152004 -4662 152186 -4426
rect 152422 -4662 152604 -4426
rect 152004 -5624 152604 -4662
rect 137604 -7162 137786 -6926
rect 138022 -7162 138204 -6926
rect 137604 -7246 138204 -7162
rect 137604 -7482 137786 -7246
rect 138022 -7482 138204 -7246
rect 137604 -7504 138204 -7482
rect 155604 -5986 156204 6000
rect 162804 5952 162832 6016
rect 162896 5952 162912 6016
rect 162976 5952 162992 6016
rect 163056 5952 163072 6016
rect 163136 5952 163152 6016
rect 163216 5952 163232 6016
rect 163296 5952 163312 6016
rect 163376 5952 163404 6016
rect 162804 4928 163404 5952
rect 162804 4864 162832 4928
rect 162896 4864 162912 4928
rect 162976 4864 162992 4928
rect 163056 4864 163072 4928
rect 163136 4864 163152 4928
rect 163216 4864 163232 4928
rect 163296 4864 163312 4928
rect 163376 4864 163404 4928
rect 162804 3840 163404 4864
rect 162804 3776 162832 3840
rect 162896 3776 162912 3840
rect 162976 3776 162992 3840
rect 163056 3776 163072 3840
rect 163136 3776 163152 3840
rect 163216 3776 163232 3840
rect 163296 3776 163312 3840
rect 163376 3776 163404 3840
rect 162804 2752 163404 3776
rect 162804 2688 162832 2752
rect 162896 2688 162912 2752
rect 162976 2688 162992 2752
rect 163056 2688 163072 2752
rect 163136 2688 163152 2752
rect 163216 2688 163232 2752
rect 163296 2688 163312 2752
rect 163376 2688 163404 2752
rect 162804 -1286 163404 2688
rect 162804 -1522 162986 -1286
rect 163222 -1522 163404 -1286
rect 162804 -1606 163404 -1522
rect 162804 -1842 162986 -1606
rect 163222 -1842 163404 -1606
rect 162804 -1864 163404 -1842
rect 166404 -3166 167004 6000
rect 166404 -3402 166586 -3166
rect 166822 -3402 167004 -3166
rect 166404 -3486 167004 -3402
rect 166404 -3722 166586 -3486
rect 166822 -3722 167004 -3486
rect 166404 -3744 167004 -3722
rect 170004 -5046 170604 6000
rect 170004 -5282 170186 -5046
rect 170422 -5282 170604 -5046
rect 170004 -5366 170604 -5282
rect 170004 -5602 170186 -5366
rect 170422 -5602 170604 -5366
rect 170004 -5624 170604 -5602
rect 155604 -6222 155786 -5986
rect 156022 -6222 156204 -5986
rect 155604 -6306 156204 -6222
rect 155604 -6542 155786 -6306
rect 156022 -6542 156204 -6306
rect 155604 -7504 156204 -6542
rect 173604 -6926 174204 6000
rect 180804 5472 181404 6048
rect 198804 6016 199404 6048
rect 180804 5408 180832 5472
rect 180896 5408 180912 5472
rect 180976 5408 180992 5472
rect 181056 5408 181072 5472
rect 181136 5408 181152 5472
rect 181216 5408 181232 5472
rect 181296 5408 181312 5472
rect 181376 5408 181404 5472
rect 180804 4384 181404 5408
rect 180804 4320 180832 4384
rect 180896 4320 180912 4384
rect 180976 4320 180992 4384
rect 181056 4320 181072 4384
rect 181136 4320 181152 4384
rect 181216 4320 181232 4384
rect 181296 4320 181312 4384
rect 181376 4320 181404 4384
rect 180804 3296 181404 4320
rect 180804 3232 180832 3296
rect 180896 3232 180912 3296
rect 180976 3232 180992 3296
rect 181056 3232 181072 3296
rect 181136 3232 181152 3296
rect 181216 3232 181232 3296
rect 181296 3232 181312 3296
rect 181376 3232 181404 3296
rect 180804 2406 181404 3232
rect 180804 2208 180986 2406
rect 181222 2208 181404 2406
rect 180804 2144 180832 2208
rect 180896 2144 180912 2208
rect 180976 2170 180986 2208
rect 181222 2170 181232 2208
rect 180976 2144 180992 2170
rect 181056 2144 181072 2170
rect 181136 2144 181152 2170
rect 181216 2144 181232 2170
rect 181296 2144 181312 2208
rect 181376 2144 181404 2208
rect 180804 2086 181404 2144
rect 180804 1850 180986 2086
rect 181222 1850 181404 2086
rect 180804 -346 181404 1850
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1864 181404 -902
rect 184404 -2226 185004 6000
rect 184404 -2462 184586 -2226
rect 184822 -2462 185004 -2226
rect 184404 -2546 185004 -2462
rect 184404 -2782 184586 -2546
rect 184822 -2782 185004 -2546
rect 184404 -3744 185004 -2782
rect 188004 -4106 188604 6000
rect 188004 -4342 188186 -4106
rect 188422 -4342 188604 -4106
rect 188004 -4426 188604 -4342
rect 188004 -4662 188186 -4426
rect 188422 -4662 188604 -4426
rect 188004 -5624 188604 -4662
rect 173604 -7162 173786 -6926
rect 174022 -7162 174204 -6926
rect 173604 -7246 174204 -7162
rect 173604 -7482 173786 -7246
rect 174022 -7482 174204 -7246
rect 173604 -7504 174204 -7482
rect 191604 -5986 192204 6000
rect 198804 5952 198832 6016
rect 198896 5952 198912 6016
rect 198976 5952 198992 6016
rect 199056 5952 199072 6016
rect 199136 5952 199152 6016
rect 199216 5952 199232 6016
rect 199296 5952 199312 6016
rect 199376 5952 199404 6016
rect 198804 4928 199404 5952
rect 198804 4864 198832 4928
rect 198896 4864 198912 4928
rect 198976 4864 198992 4928
rect 199056 4864 199072 4928
rect 199136 4864 199152 4928
rect 199216 4864 199232 4928
rect 199296 4864 199312 4928
rect 199376 4864 199404 4928
rect 198804 3840 199404 4864
rect 198804 3776 198832 3840
rect 198896 3776 198912 3840
rect 198976 3776 198992 3840
rect 199056 3776 199072 3840
rect 199136 3776 199152 3840
rect 199216 3776 199232 3840
rect 199296 3776 199312 3840
rect 199376 3776 199404 3840
rect 198804 2752 199404 3776
rect 198804 2688 198832 2752
rect 198896 2688 198912 2752
rect 198976 2688 198992 2752
rect 199056 2688 199072 2752
rect 199136 2688 199152 2752
rect 199216 2688 199232 2752
rect 199296 2688 199312 2752
rect 199376 2688 199404 2752
rect 198804 -1286 199404 2688
rect 198804 -1522 198986 -1286
rect 199222 -1522 199404 -1286
rect 198804 -1606 199404 -1522
rect 198804 -1842 198986 -1606
rect 199222 -1842 199404 -1606
rect 198804 -1864 199404 -1842
rect 202404 -3166 203004 6000
rect 202404 -3402 202586 -3166
rect 202822 -3402 203004 -3166
rect 202404 -3486 203004 -3402
rect 202404 -3722 202586 -3486
rect 202822 -3722 203004 -3486
rect 202404 -3744 203004 -3722
rect 206004 -5046 206604 6000
rect 206004 -5282 206186 -5046
rect 206422 -5282 206604 -5046
rect 206004 -5366 206604 -5282
rect 206004 -5602 206186 -5366
rect 206422 -5602 206604 -5366
rect 206004 -5624 206604 -5602
rect 191604 -6222 191786 -5986
rect 192022 -6222 192204 -5986
rect 191604 -6306 192204 -6222
rect 191604 -6542 191786 -6306
rect 192022 -6542 192204 -6306
rect 191604 -7504 192204 -6542
rect 209604 -6926 210204 6000
rect 216804 5472 217404 6048
rect 234804 6016 235404 6048
rect 216804 5408 216832 5472
rect 216896 5408 216912 5472
rect 216976 5408 216992 5472
rect 217056 5408 217072 5472
rect 217136 5408 217152 5472
rect 217216 5408 217232 5472
rect 217296 5408 217312 5472
rect 217376 5408 217404 5472
rect 216804 4384 217404 5408
rect 216804 4320 216832 4384
rect 216896 4320 216912 4384
rect 216976 4320 216992 4384
rect 217056 4320 217072 4384
rect 217136 4320 217152 4384
rect 217216 4320 217232 4384
rect 217296 4320 217312 4384
rect 217376 4320 217404 4384
rect 216804 3296 217404 4320
rect 216804 3232 216832 3296
rect 216896 3232 216912 3296
rect 216976 3232 216992 3296
rect 217056 3232 217072 3296
rect 217136 3232 217152 3296
rect 217216 3232 217232 3296
rect 217296 3232 217312 3296
rect 217376 3232 217404 3296
rect 216804 2406 217404 3232
rect 216804 2208 216986 2406
rect 217222 2208 217404 2406
rect 216804 2144 216832 2208
rect 216896 2144 216912 2208
rect 216976 2170 216986 2208
rect 217222 2170 217232 2208
rect 216976 2144 216992 2170
rect 217056 2144 217072 2170
rect 217136 2144 217152 2170
rect 217216 2144 217232 2170
rect 217296 2144 217312 2208
rect 217376 2144 217404 2208
rect 216804 2086 217404 2144
rect 216804 1850 216986 2086
rect 217222 1850 217404 2086
rect 216804 -346 217404 1850
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1864 217404 -902
rect 220404 -2226 221004 6000
rect 220404 -2462 220586 -2226
rect 220822 -2462 221004 -2226
rect 220404 -2546 221004 -2462
rect 220404 -2782 220586 -2546
rect 220822 -2782 221004 -2546
rect 220404 -3744 221004 -2782
rect 224004 -4106 224604 6000
rect 224004 -4342 224186 -4106
rect 224422 -4342 224604 -4106
rect 224004 -4426 224604 -4342
rect 224004 -4662 224186 -4426
rect 224422 -4662 224604 -4426
rect 224004 -5624 224604 -4662
rect 209604 -7162 209786 -6926
rect 210022 -7162 210204 -6926
rect 209604 -7246 210204 -7162
rect 209604 -7482 209786 -7246
rect 210022 -7482 210204 -7246
rect 209604 -7504 210204 -7482
rect 227604 -5986 228204 6000
rect 234804 5952 234832 6016
rect 234896 5952 234912 6016
rect 234976 5952 234992 6016
rect 235056 5952 235072 6016
rect 235136 5952 235152 6016
rect 235216 5952 235232 6016
rect 235296 5952 235312 6016
rect 235376 5952 235404 6016
rect 234804 4928 235404 5952
rect 234804 4864 234832 4928
rect 234896 4864 234912 4928
rect 234976 4864 234992 4928
rect 235056 4864 235072 4928
rect 235136 4864 235152 4928
rect 235216 4864 235232 4928
rect 235296 4864 235312 4928
rect 235376 4864 235404 4928
rect 234804 3840 235404 4864
rect 234804 3776 234832 3840
rect 234896 3776 234912 3840
rect 234976 3776 234992 3840
rect 235056 3776 235072 3840
rect 235136 3776 235152 3840
rect 235216 3776 235232 3840
rect 235296 3776 235312 3840
rect 235376 3776 235404 3840
rect 234804 2752 235404 3776
rect 234804 2688 234832 2752
rect 234896 2688 234912 2752
rect 234976 2688 234992 2752
rect 235056 2688 235072 2752
rect 235136 2688 235152 2752
rect 235216 2688 235232 2752
rect 235296 2688 235312 2752
rect 235376 2688 235404 2752
rect 234804 -1286 235404 2688
rect 234804 -1522 234986 -1286
rect 235222 -1522 235404 -1286
rect 234804 -1606 235404 -1522
rect 234804 -1842 234986 -1606
rect 235222 -1842 235404 -1606
rect 234804 -1864 235404 -1842
rect 238404 -3166 239004 6000
rect 238404 -3402 238586 -3166
rect 238822 -3402 239004 -3166
rect 238404 -3486 239004 -3402
rect 238404 -3722 238586 -3486
rect 238822 -3722 239004 -3486
rect 238404 -3744 239004 -3722
rect 242004 -5046 242604 6000
rect 242004 -5282 242186 -5046
rect 242422 -5282 242604 -5046
rect 242004 -5366 242604 -5282
rect 242004 -5602 242186 -5366
rect 242422 -5602 242604 -5366
rect 242004 -5624 242604 -5602
rect 227604 -6222 227786 -5986
rect 228022 -6222 228204 -5986
rect 227604 -6306 228204 -6222
rect 227604 -6542 227786 -6306
rect 228022 -6542 228204 -6306
rect 227604 -7504 228204 -6542
rect 245604 -6926 246204 6000
rect 252804 5472 253404 6048
rect 270804 6016 271404 6048
rect 252804 5408 252832 5472
rect 252896 5408 252912 5472
rect 252976 5408 252992 5472
rect 253056 5408 253072 5472
rect 253136 5408 253152 5472
rect 253216 5408 253232 5472
rect 253296 5408 253312 5472
rect 253376 5408 253404 5472
rect 252804 4384 253404 5408
rect 252804 4320 252832 4384
rect 252896 4320 252912 4384
rect 252976 4320 252992 4384
rect 253056 4320 253072 4384
rect 253136 4320 253152 4384
rect 253216 4320 253232 4384
rect 253296 4320 253312 4384
rect 253376 4320 253404 4384
rect 252804 3296 253404 4320
rect 252804 3232 252832 3296
rect 252896 3232 252912 3296
rect 252976 3232 252992 3296
rect 253056 3232 253072 3296
rect 253136 3232 253152 3296
rect 253216 3232 253232 3296
rect 253296 3232 253312 3296
rect 253376 3232 253404 3296
rect 252804 2406 253404 3232
rect 252804 2208 252986 2406
rect 253222 2208 253404 2406
rect 252804 2144 252832 2208
rect 252896 2144 252912 2208
rect 252976 2170 252986 2208
rect 253222 2170 253232 2208
rect 252976 2144 252992 2170
rect 253056 2144 253072 2170
rect 253136 2144 253152 2170
rect 253216 2144 253232 2170
rect 253296 2144 253312 2208
rect 253376 2144 253404 2208
rect 252804 2086 253404 2144
rect 252804 1850 252986 2086
rect 253222 1850 253404 2086
rect 252804 -346 253404 1850
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1864 253404 -902
rect 256404 -2226 257004 6000
rect 256404 -2462 256586 -2226
rect 256822 -2462 257004 -2226
rect 256404 -2546 257004 -2462
rect 256404 -2782 256586 -2546
rect 256822 -2782 257004 -2546
rect 256404 -3744 257004 -2782
rect 260004 -4106 260604 6000
rect 260004 -4342 260186 -4106
rect 260422 -4342 260604 -4106
rect 260004 -4426 260604 -4342
rect 260004 -4662 260186 -4426
rect 260422 -4662 260604 -4426
rect 260004 -5624 260604 -4662
rect 245604 -7162 245786 -6926
rect 246022 -7162 246204 -6926
rect 245604 -7246 246204 -7162
rect 245604 -7482 245786 -7246
rect 246022 -7482 246204 -7246
rect 245604 -7504 246204 -7482
rect 263604 -5986 264204 6000
rect 270804 5952 270832 6016
rect 270896 5952 270912 6016
rect 270976 5952 270992 6016
rect 271056 5952 271072 6016
rect 271136 5952 271152 6016
rect 271216 5952 271232 6016
rect 271296 5952 271312 6016
rect 271376 5952 271404 6016
rect 270804 4928 271404 5952
rect 270804 4864 270832 4928
rect 270896 4864 270912 4928
rect 270976 4864 270992 4928
rect 271056 4864 271072 4928
rect 271136 4864 271152 4928
rect 271216 4864 271232 4928
rect 271296 4864 271312 4928
rect 271376 4864 271404 4928
rect 270804 3840 271404 4864
rect 270804 3776 270832 3840
rect 270896 3776 270912 3840
rect 270976 3776 270992 3840
rect 271056 3776 271072 3840
rect 271136 3776 271152 3840
rect 271216 3776 271232 3840
rect 271296 3776 271312 3840
rect 271376 3776 271404 3840
rect 270804 2752 271404 3776
rect 270804 2688 270832 2752
rect 270896 2688 270912 2752
rect 270976 2688 270992 2752
rect 271056 2688 271072 2752
rect 271136 2688 271152 2752
rect 271216 2688 271232 2752
rect 271296 2688 271312 2752
rect 271376 2688 271404 2752
rect 270804 -1286 271404 2688
rect 270804 -1522 270986 -1286
rect 271222 -1522 271404 -1286
rect 270804 -1606 271404 -1522
rect 270804 -1842 270986 -1606
rect 271222 -1842 271404 -1606
rect 270804 -1864 271404 -1842
rect 274404 -3166 275004 6000
rect 274404 -3402 274586 -3166
rect 274822 -3402 275004 -3166
rect 274404 -3486 275004 -3402
rect 274404 -3722 274586 -3486
rect 274822 -3722 275004 -3486
rect 274404 -3744 275004 -3722
rect 278004 -5046 278604 6000
rect 278004 -5282 278186 -5046
rect 278422 -5282 278604 -5046
rect 278004 -5366 278604 -5282
rect 278004 -5602 278186 -5366
rect 278422 -5602 278604 -5366
rect 278004 -5624 278604 -5602
rect 263604 -6222 263786 -5986
rect 264022 -6222 264204 -5986
rect 263604 -6306 264204 -6222
rect 263604 -6542 263786 -6306
rect 264022 -6542 264204 -6306
rect 263604 -7504 264204 -6542
rect 281604 -6926 282204 6000
rect 288804 5472 289404 6048
rect 306804 6016 307404 6048
rect 288804 5408 288832 5472
rect 288896 5408 288912 5472
rect 288976 5408 288992 5472
rect 289056 5408 289072 5472
rect 289136 5408 289152 5472
rect 289216 5408 289232 5472
rect 289296 5408 289312 5472
rect 289376 5408 289404 5472
rect 288804 4384 289404 5408
rect 288804 4320 288832 4384
rect 288896 4320 288912 4384
rect 288976 4320 288992 4384
rect 289056 4320 289072 4384
rect 289136 4320 289152 4384
rect 289216 4320 289232 4384
rect 289296 4320 289312 4384
rect 289376 4320 289404 4384
rect 288804 3296 289404 4320
rect 288804 3232 288832 3296
rect 288896 3232 288912 3296
rect 288976 3232 288992 3296
rect 289056 3232 289072 3296
rect 289136 3232 289152 3296
rect 289216 3232 289232 3296
rect 289296 3232 289312 3296
rect 289376 3232 289404 3296
rect 288804 2406 289404 3232
rect 288804 2208 288986 2406
rect 289222 2208 289404 2406
rect 288804 2144 288832 2208
rect 288896 2144 288912 2208
rect 288976 2170 288986 2208
rect 289222 2170 289232 2208
rect 288976 2144 288992 2170
rect 289056 2144 289072 2170
rect 289136 2144 289152 2170
rect 289216 2144 289232 2170
rect 289296 2144 289312 2208
rect 289376 2144 289404 2208
rect 288804 2086 289404 2144
rect 288804 1850 288986 2086
rect 289222 1850 289404 2086
rect 288804 -346 289404 1850
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1864 289404 -902
rect 292404 -2226 293004 6000
rect 292404 -2462 292586 -2226
rect 292822 -2462 293004 -2226
rect 292404 -2546 293004 -2462
rect 292404 -2782 292586 -2546
rect 292822 -2782 293004 -2546
rect 292404 -3744 293004 -2782
rect 296004 -4106 296604 6000
rect 296004 -4342 296186 -4106
rect 296422 -4342 296604 -4106
rect 296004 -4426 296604 -4342
rect 296004 -4662 296186 -4426
rect 296422 -4662 296604 -4426
rect 296004 -5624 296604 -4662
rect 281604 -7162 281786 -6926
rect 282022 -7162 282204 -6926
rect 281604 -7246 282204 -7162
rect 281604 -7482 281786 -7246
rect 282022 -7482 282204 -7246
rect 281604 -7504 282204 -7482
rect 299604 -5986 300204 6000
rect 306804 5952 306832 6016
rect 306896 5952 306912 6016
rect 306976 5952 306992 6016
rect 307056 5952 307072 6016
rect 307136 5952 307152 6016
rect 307216 5952 307232 6016
rect 307296 5952 307312 6016
rect 307376 5952 307404 6016
rect 306804 4928 307404 5952
rect 306804 4864 306832 4928
rect 306896 4864 306912 4928
rect 306976 4864 306992 4928
rect 307056 4864 307072 4928
rect 307136 4864 307152 4928
rect 307216 4864 307232 4928
rect 307296 4864 307312 4928
rect 307376 4864 307404 4928
rect 306804 3840 307404 4864
rect 306804 3776 306832 3840
rect 306896 3776 306912 3840
rect 306976 3776 306992 3840
rect 307056 3776 307072 3840
rect 307136 3776 307152 3840
rect 307216 3776 307232 3840
rect 307296 3776 307312 3840
rect 307376 3776 307404 3840
rect 306804 2752 307404 3776
rect 306804 2688 306832 2752
rect 306896 2688 306912 2752
rect 306976 2688 306992 2752
rect 307056 2688 307072 2752
rect 307136 2688 307152 2752
rect 307216 2688 307232 2752
rect 307296 2688 307312 2752
rect 307376 2688 307404 2752
rect 306804 -1286 307404 2688
rect 306804 -1522 306986 -1286
rect 307222 -1522 307404 -1286
rect 306804 -1606 307404 -1522
rect 306804 -1842 306986 -1606
rect 307222 -1842 307404 -1606
rect 306804 -1864 307404 -1842
rect 310404 -3166 311004 6000
rect 310404 -3402 310586 -3166
rect 310822 -3402 311004 -3166
rect 310404 -3486 311004 -3402
rect 310404 -3722 310586 -3486
rect 310822 -3722 311004 -3486
rect 310404 -3744 311004 -3722
rect 314004 -5046 314604 6000
rect 314004 -5282 314186 -5046
rect 314422 -5282 314604 -5046
rect 314004 -5366 314604 -5282
rect 314004 -5602 314186 -5366
rect 314422 -5602 314604 -5366
rect 314004 -5624 314604 -5602
rect 299604 -6222 299786 -5986
rect 300022 -6222 300204 -5986
rect 299604 -6306 300204 -6222
rect 299604 -6542 299786 -6306
rect 300022 -6542 300204 -6306
rect 299604 -7504 300204 -6542
rect 317604 -6926 318204 6000
rect 324804 5472 325404 6048
rect 342804 6016 343404 6048
rect 324804 5408 324832 5472
rect 324896 5408 324912 5472
rect 324976 5408 324992 5472
rect 325056 5408 325072 5472
rect 325136 5408 325152 5472
rect 325216 5408 325232 5472
rect 325296 5408 325312 5472
rect 325376 5408 325404 5472
rect 324804 4384 325404 5408
rect 324804 4320 324832 4384
rect 324896 4320 324912 4384
rect 324976 4320 324992 4384
rect 325056 4320 325072 4384
rect 325136 4320 325152 4384
rect 325216 4320 325232 4384
rect 325296 4320 325312 4384
rect 325376 4320 325404 4384
rect 324804 3296 325404 4320
rect 324804 3232 324832 3296
rect 324896 3232 324912 3296
rect 324976 3232 324992 3296
rect 325056 3232 325072 3296
rect 325136 3232 325152 3296
rect 325216 3232 325232 3296
rect 325296 3232 325312 3296
rect 325376 3232 325404 3296
rect 324804 2406 325404 3232
rect 324804 2208 324986 2406
rect 325222 2208 325404 2406
rect 324804 2144 324832 2208
rect 324896 2144 324912 2208
rect 324976 2170 324986 2208
rect 325222 2170 325232 2208
rect 324976 2144 324992 2170
rect 325056 2144 325072 2170
rect 325136 2144 325152 2170
rect 325216 2144 325232 2170
rect 325296 2144 325312 2208
rect 325376 2144 325404 2208
rect 324804 2086 325404 2144
rect 324804 1850 324986 2086
rect 325222 1850 325404 2086
rect 324804 -346 325404 1850
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1864 325404 -902
rect 328404 -2226 329004 6000
rect 328404 -2462 328586 -2226
rect 328822 -2462 329004 -2226
rect 328404 -2546 329004 -2462
rect 328404 -2782 328586 -2546
rect 328822 -2782 329004 -2546
rect 328404 -3744 329004 -2782
rect 332004 -4106 332604 6000
rect 332004 -4342 332186 -4106
rect 332422 -4342 332604 -4106
rect 332004 -4426 332604 -4342
rect 332004 -4662 332186 -4426
rect 332422 -4662 332604 -4426
rect 332004 -5624 332604 -4662
rect 317604 -7162 317786 -6926
rect 318022 -7162 318204 -6926
rect 317604 -7246 318204 -7162
rect 317604 -7482 317786 -7246
rect 318022 -7482 318204 -7246
rect 317604 -7504 318204 -7482
rect 335604 -5986 336204 6000
rect 342804 5952 342832 6016
rect 342896 5952 342912 6016
rect 342976 5952 342992 6016
rect 343056 5952 343072 6016
rect 343136 5952 343152 6016
rect 343216 5952 343232 6016
rect 343296 5952 343312 6016
rect 343376 5952 343404 6016
rect 342804 4928 343404 5952
rect 342804 4864 342832 4928
rect 342896 4864 342912 4928
rect 342976 4864 342992 4928
rect 343056 4864 343072 4928
rect 343136 4864 343152 4928
rect 343216 4864 343232 4928
rect 343296 4864 343312 4928
rect 343376 4864 343404 4928
rect 342804 3840 343404 4864
rect 342804 3776 342832 3840
rect 342896 3776 342912 3840
rect 342976 3776 342992 3840
rect 343056 3776 343072 3840
rect 343136 3776 343152 3840
rect 343216 3776 343232 3840
rect 343296 3776 343312 3840
rect 343376 3776 343404 3840
rect 342804 2752 343404 3776
rect 342804 2688 342832 2752
rect 342896 2688 342912 2752
rect 342976 2688 342992 2752
rect 343056 2688 343072 2752
rect 343136 2688 343152 2752
rect 343216 2688 343232 2752
rect 343296 2688 343312 2752
rect 343376 2688 343404 2752
rect 342804 -1286 343404 2688
rect 342804 -1522 342986 -1286
rect 343222 -1522 343404 -1286
rect 342804 -1606 343404 -1522
rect 342804 -1842 342986 -1606
rect 343222 -1842 343404 -1606
rect 342804 -1864 343404 -1842
rect 346404 -3166 347004 6000
rect 346404 -3402 346586 -3166
rect 346822 -3402 347004 -3166
rect 346404 -3486 347004 -3402
rect 346404 -3722 346586 -3486
rect 346822 -3722 347004 -3486
rect 346404 -3744 347004 -3722
rect 350004 -5046 350604 6000
rect 350004 -5282 350186 -5046
rect 350422 -5282 350604 -5046
rect 350004 -5366 350604 -5282
rect 350004 -5602 350186 -5366
rect 350422 -5602 350604 -5366
rect 350004 -5624 350604 -5602
rect 335604 -6222 335786 -5986
rect 336022 -6222 336204 -5986
rect 335604 -6306 336204 -6222
rect 335604 -6542 335786 -6306
rect 336022 -6542 336204 -6306
rect 335604 -7504 336204 -6542
rect 353604 -6926 354204 6000
rect 360804 5472 361404 6048
rect 378804 6016 379404 6048
rect 360804 5408 360832 5472
rect 360896 5408 360912 5472
rect 360976 5408 360992 5472
rect 361056 5408 361072 5472
rect 361136 5408 361152 5472
rect 361216 5408 361232 5472
rect 361296 5408 361312 5472
rect 361376 5408 361404 5472
rect 360804 4384 361404 5408
rect 360804 4320 360832 4384
rect 360896 4320 360912 4384
rect 360976 4320 360992 4384
rect 361056 4320 361072 4384
rect 361136 4320 361152 4384
rect 361216 4320 361232 4384
rect 361296 4320 361312 4384
rect 361376 4320 361404 4384
rect 360804 3296 361404 4320
rect 360804 3232 360832 3296
rect 360896 3232 360912 3296
rect 360976 3232 360992 3296
rect 361056 3232 361072 3296
rect 361136 3232 361152 3296
rect 361216 3232 361232 3296
rect 361296 3232 361312 3296
rect 361376 3232 361404 3296
rect 360804 2406 361404 3232
rect 360804 2208 360986 2406
rect 361222 2208 361404 2406
rect 360804 2144 360832 2208
rect 360896 2144 360912 2208
rect 360976 2170 360986 2208
rect 361222 2170 361232 2208
rect 360976 2144 360992 2170
rect 361056 2144 361072 2170
rect 361136 2144 361152 2170
rect 361216 2144 361232 2170
rect 361296 2144 361312 2208
rect 361376 2144 361404 2208
rect 360804 2086 361404 2144
rect 360804 1850 360986 2086
rect 361222 1850 361404 2086
rect 360804 -346 361404 1850
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1864 361404 -902
rect 364404 -2226 365004 6000
rect 364404 -2462 364586 -2226
rect 364822 -2462 365004 -2226
rect 364404 -2546 365004 -2462
rect 364404 -2782 364586 -2546
rect 364822 -2782 365004 -2546
rect 364404 -3744 365004 -2782
rect 368004 -4106 368604 6000
rect 368004 -4342 368186 -4106
rect 368422 -4342 368604 -4106
rect 368004 -4426 368604 -4342
rect 368004 -4662 368186 -4426
rect 368422 -4662 368604 -4426
rect 368004 -5624 368604 -4662
rect 353604 -7162 353786 -6926
rect 354022 -7162 354204 -6926
rect 353604 -7246 354204 -7162
rect 353604 -7482 353786 -7246
rect 354022 -7482 354204 -7246
rect 353604 -7504 354204 -7482
rect 371604 -5986 372204 6000
rect 378804 5952 378832 6016
rect 378896 5952 378912 6016
rect 378976 5952 378992 6016
rect 379056 5952 379072 6016
rect 379136 5952 379152 6016
rect 379216 5952 379232 6016
rect 379296 5952 379312 6016
rect 379376 5952 379404 6016
rect 378804 4928 379404 5952
rect 378804 4864 378832 4928
rect 378896 4864 378912 4928
rect 378976 4864 378992 4928
rect 379056 4864 379072 4928
rect 379136 4864 379152 4928
rect 379216 4864 379232 4928
rect 379296 4864 379312 4928
rect 379376 4864 379404 4928
rect 378804 3840 379404 4864
rect 378804 3776 378832 3840
rect 378896 3776 378912 3840
rect 378976 3776 378992 3840
rect 379056 3776 379072 3840
rect 379136 3776 379152 3840
rect 379216 3776 379232 3840
rect 379296 3776 379312 3840
rect 379376 3776 379404 3840
rect 378804 2752 379404 3776
rect 378804 2688 378832 2752
rect 378896 2688 378912 2752
rect 378976 2688 378992 2752
rect 379056 2688 379072 2752
rect 379136 2688 379152 2752
rect 379216 2688 379232 2752
rect 379296 2688 379312 2752
rect 379376 2688 379404 2752
rect 378804 -1286 379404 2688
rect 378804 -1522 378986 -1286
rect 379222 -1522 379404 -1286
rect 378804 -1606 379404 -1522
rect 378804 -1842 378986 -1606
rect 379222 -1842 379404 -1606
rect 378804 -1864 379404 -1842
rect 382404 -3166 383004 6000
rect 382404 -3402 382586 -3166
rect 382822 -3402 383004 -3166
rect 382404 -3486 383004 -3402
rect 382404 -3722 382586 -3486
rect 382822 -3722 383004 -3486
rect 382404 -3744 383004 -3722
rect 386004 -5046 386604 6000
rect 386004 -5282 386186 -5046
rect 386422 -5282 386604 -5046
rect 386004 -5366 386604 -5282
rect 386004 -5602 386186 -5366
rect 386422 -5602 386604 -5366
rect 386004 -5624 386604 -5602
rect 371604 -6222 371786 -5986
rect 372022 -6222 372204 -5986
rect 371604 -6306 372204 -6222
rect 371604 -6542 371786 -6306
rect 372022 -6542 372204 -6306
rect 371604 -7504 372204 -6542
rect 389604 -6926 390204 6000
rect 396804 5472 397404 6048
rect 414804 6016 415404 6048
rect 396804 5408 396832 5472
rect 396896 5408 396912 5472
rect 396976 5408 396992 5472
rect 397056 5408 397072 5472
rect 397136 5408 397152 5472
rect 397216 5408 397232 5472
rect 397296 5408 397312 5472
rect 397376 5408 397404 5472
rect 396804 4384 397404 5408
rect 396804 4320 396832 4384
rect 396896 4320 396912 4384
rect 396976 4320 396992 4384
rect 397056 4320 397072 4384
rect 397136 4320 397152 4384
rect 397216 4320 397232 4384
rect 397296 4320 397312 4384
rect 397376 4320 397404 4384
rect 396804 3296 397404 4320
rect 396804 3232 396832 3296
rect 396896 3232 396912 3296
rect 396976 3232 396992 3296
rect 397056 3232 397072 3296
rect 397136 3232 397152 3296
rect 397216 3232 397232 3296
rect 397296 3232 397312 3296
rect 397376 3232 397404 3296
rect 396804 2406 397404 3232
rect 396804 2208 396986 2406
rect 397222 2208 397404 2406
rect 396804 2144 396832 2208
rect 396896 2144 396912 2208
rect 396976 2170 396986 2208
rect 397222 2170 397232 2208
rect 396976 2144 396992 2170
rect 397056 2144 397072 2170
rect 397136 2144 397152 2170
rect 397216 2144 397232 2170
rect 397296 2144 397312 2208
rect 397376 2144 397404 2208
rect 396804 2086 397404 2144
rect 396804 1850 396986 2086
rect 397222 1850 397404 2086
rect 396804 -346 397404 1850
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1864 397404 -902
rect 400404 -2226 401004 6000
rect 400404 -2462 400586 -2226
rect 400822 -2462 401004 -2226
rect 400404 -2546 401004 -2462
rect 400404 -2782 400586 -2546
rect 400822 -2782 401004 -2546
rect 400404 -3744 401004 -2782
rect 404004 -4106 404604 6000
rect 404004 -4342 404186 -4106
rect 404422 -4342 404604 -4106
rect 404004 -4426 404604 -4342
rect 404004 -4662 404186 -4426
rect 404422 -4662 404604 -4426
rect 404004 -5624 404604 -4662
rect 389604 -7162 389786 -6926
rect 390022 -7162 390204 -6926
rect 389604 -7246 390204 -7162
rect 389604 -7482 389786 -7246
rect 390022 -7482 390204 -7246
rect 389604 -7504 390204 -7482
rect 407604 -5986 408204 6000
rect 414804 5952 414832 6016
rect 414896 5952 414912 6016
rect 414976 5952 414992 6016
rect 415056 5952 415072 6016
rect 415136 5952 415152 6016
rect 415216 5952 415232 6016
rect 415296 5952 415312 6016
rect 415376 5952 415404 6016
rect 414804 4928 415404 5952
rect 414804 4864 414832 4928
rect 414896 4864 414912 4928
rect 414976 4864 414992 4928
rect 415056 4864 415072 4928
rect 415136 4864 415152 4928
rect 415216 4864 415232 4928
rect 415296 4864 415312 4928
rect 415376 4864 415404 4928
rect 414804 3840 415404 4864
rect 414804 3776 414832 3840
rect 414896 3776 414912 3840
rect 414976 3776 414992 3840
rect 415056 3776 415072 3840
rect 415136 3776 415152 3840
rect 415216 3776 415232 3840
rect 415296 3776 415312 3840
rect 415376 3776 415404 3840
rect 414804 2752 415404 3776
rect 414804 2688 414832 2752
rect 414896 2688 414912 2752
rect 414976 2688 414992 2752
rect 415056 2688 415072 2752
rect 415136 2688 415152 2752
rect 415216 2688 415232 2752
rect 415296 2688 415312 2752
rect 415376 2688 415404 2752
rect 414804 -1286 415404 2688
rect 414804 -1522 414986 -1286
rect 415222 -1522 415404 -1286
rect 414804 -1606 415404 -1522
rect 414804 -1842 414986 -1606
rect 415222 -1842 415404 -1606
rect 414804 -1864 415404 -1842
rect 418404 -3166 419004 6000
rect 418404 -3402 418586 -3166
rect 418822 -3402 419004 -3166
rect 418404 -3486 419004 -3402
rect 418404 -3722 418586 -3486
rect 418822 -3722 419004 -3486
rect 418404 -3744 419004 -3722
rect 422004 -5046 422604 6000
rect 422004 -5282 422186 -5046
rect 422422 -5282 422604 -5046
rect 422004 -5366 422604 -5282
rect 422004 -5602 422186 -5366
rect 422422 -5602 422604 -5366
rect 422004 -5624 422604 -5602
rect 407604 -6222 407786 -5986
rect 408022 -6222 408204 -5986
rect 407604 -6306 408204 -6222
rect 407604 -6542 407786 -6306
rect 408022 -6542 408204 -6306
rect 407604 -7504 408204 -6542
rect 425604 -6926 426204 6000
rect 432804 5472 433404 6048
rect 450804 6016 451404 6048
rect 432804 5408 432832 5472
rect 432896 5408 432912 5472
rect 432976 5408 432992 5472
rect 433056 5408 433072 5472
rect 433136 5408 433152 5472
rect 433216 5408 433232 5472
rect 433296 5408 433312 5472
rect 433376 5408 433404 5472
rect 432804 4384 433404 5408
rect 432804 4320 432832 4384
rect 432896 4320 432912 4384
rect 432976 4320 432992 4384
rect 433056 4320 433072 4384
rect 433136 4320 433152 4384
rect 433216 4320 433232 4384
rect 433296 4320 433312 4384
rect 433376 4320 433404 4384
rect 432804 3296 433404 4320
rect 432804 3232 432832 3296
rect 432896 3232 432912 3296
rect 432976 3232 432992 3296
rect 433056 3232 433072 3296
rect 433136 3232 433152 3296
rect 433216 3232 433232 3296
rect 433296 3232 433312 3296
rect 433376 3232 433404 3296
rect 432804 2406 433404 3232
rect 432804 2208 432986 2406
rect 433222 2208 433404 2406
rect 432804 2144 432832 2208
rect 432896 2144 432912 2208
rect 432976 2170 432986 2208
rect 433222 2170 433232 2208
rect 432976 2144 432992 2170
rect 433056 2144 433072 2170
rect 433136 2144 433152 2170
rect 433216 2144 433232 2170
rect 433296 2144 433312 2208
rect 433376 2144 433404 2208
rect 432804 2086 433404 2144
rect 432804 1850 432986 2086
rect 433222 1850 433404 2086
rect 432804 -346 433404 1850
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1864 433404 -902
rect 436404 -2226 437004 6000
rect 436404 -2462 436586 -2226
rect 436822 -2462 437004 -2226
rect 436404 -2546 437004 -2462
rect 436404 -2782 436586 -2546
rect 436822 -2782 437004 -2546
rect 436404 -3744 437004 -2782
rect 440004 -4106 440604 6000
rect 440004 -4342 440186 -4106
rect 440422 -4342 440604 -4106
rect 440004 -4426 440604 -4342
rect 440004 -4662 440186 -4426
rect 440422 -4662 440604 -4426
rect 440004 -5624 440604 -4662
rect 425604 -7162 425786 -6926
rect 426022 -7162 426204 -6926
rect 425604 -7246 426204 -7162
rect 425604 -7482 425786 -7246
rect 426022 -7482 426204 -7246
rect 425604 -7504 426204 -7482
rect 443604 -5986 444204 6000
rect 450804 5952 450832 6016
rect 450896 5952 450912 6016
rect 450976 5952 450992 6016
rect 451056 5952 451072 6016
rect 451136 5952 451152 6016
rect 451216 5952 451232 6016
rect 451296 5952 451312 6016
rect 451376 5952 451404 6016
rect 450804 4928 451404 5952
rect 450804 4864 450832 4928
rect 450896 4864 450912 4928
rect 450976 4864 450992 4928
rect 451056 4864 451072 4928
rect 451136 4864 451152 4928
rect 451216 4864 451232 4928
rect 451296 4864 451312 4928
rect 451376 4864 451404 4928
rect 450804 3840 451404 4864
rect 450804 3776 450832 3840
rect 450896 3776 450912 3840
rect 450976 3776 450992 3840
rect 451056 3776 451072 3840
rect 451136 3776 451152 3840
rect 451216 3776 451232 3840
rect 451296 3776 451312 3840
rect 451376 3776 451404 3840
rect 450804 2752 451404 3776
rect 450804 2688 450832 2752
rect 450896 2688 450912 2752
rect 450976 2688 450992 2752
rect 451056 2688 451072 2752
rect 451136 2688 451152 2752
rect 451216 2688 451232 2752
rect 451296 2688 451312 2752
rect 451376 2688 451404 2752
rect 450804 -1286 451404 2688
rect 450804 -1522 450986 -1286
rect 451222 -1522 451404 -1286
rect 450804 -1606 451404 -1522
rect 450804 -1842 450986 -1606
rect 451222 -1842 451404 -1606
rect 450804 -1864 451404 -1842
rect 454404 -3166 455004 6000
rect 454404 -3402 454586 -3166
rect 454822 -3402 455004 -3166
rect 454404 -3486 455004 -3402
rect 454404 -3722 454586 -3486
rect 454822 -3722 455004 -3486
rect 454404 -3744 455004 -3722
rect 458004 -5046 458604 6000
rect 458004 -5282 458186 -5046
rect 458422 -5282 458604 -5046
rect 458004 -5366 458604 -5282
rect 458004 -5602 458186 -5366
rect 458422 -5602 458604 -5366
rect 458004 -5624 458604 -5602
rect 443604 -6222 443786 -5986
rect 444022 -6222 444204 -5986
rect 443604 -6306 444204 -6222
rect 443604 -6542 443786 -6306
rect 444022 -6542 444204 -6306
rect 443604 -7504 444204 -6542
rect 461604 -6926 462204 6000
rect 468804 5472 469404 6048
rect 486804 6016 487404 6048
rect 468804 5408 468832 5472
rect 468896 5408 468912 5472
rect 468976 5408 468992 5472
rect 469056 5408 469072 5472
rect 469136 5408 469152 5472
rect 469216 5408 469232 5472
rect 469296 5408 469312 5472
rect 469376 5408 469404 5472
rect 468804 4384 469404 5408
rect 468804 4320 468832 4384
rect 468896 4320 468912 4384
rect 468976 4320 468992 4384
rect 469056 4320 469072 4384
rect 469136 4320 469152 4384
rect 469216 4320 469232 4384
rect 469296 4320 469312 4384
rect 469376 4320 469404 4384
rect 468804 3296 469404 4320
rect 468804 3232 468832 3296
rect 468896 3232 468912 3296
rect 468976 3232 468992 3296
rect 469056 3232 469072 3296
rect 469136 3232 469152 3296
rect 469216 3232 469232 3296
rect 469296 3232 469312 3296
rect 469376 3232 469404 3296
rect 468804 2406 469404 3232
rect 468804 2208 468986 2406
rect 469222 2208 469404 2406
rect 468804 2144 468832 2208
rect 468896 2144 468912 2208
rect 468976 2170 468986 2208
rect 469222 2170 469232 2208
rect 468976 2144 468992 2170
rect 469056 2144 469072 2170
rect 469136 2144 469152 2170
rect 469216 2144 469232 2170
rect 469296 2144 469312 2208
rect 469376 2144 469404 2208
rect 468804 2086 469404 2144
rect 468804 1850 468986 2086
rect 469222 1850 469404 2086
rect 468804 -346 469404 1850
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1864 469404 -902
rect 472404 -2226 473004 6000
rect 472404 -2462 472586 -2226
rect 472822 -2462 473004 -2226
rect 472404 -2546 473004 -2462
rect 472404 -2782 472586 -2546
rect 472822 -2782 473004 -2546
rect 472404 -3744 473004 -2782
rect 476004 -4106 476604 6000
rect 476004 -4342 476186 -4106
rect 476422 -4342 476604 -4106
rect 476004 -4426 476604 -4342
rect 476004 -4662 476186 -4426
rect 476422 -4662 476604 -4426
rect 476004 -5624 476604 -4662
rect 461604 -7162 461786 -6926
rect 462022 -7162 462204 -6926
rect 461604 -7246 462204 -7162
rect 461604 -7482 461786 -7246
rect 462022 -7482 462204 -7246
rect 461604 -7504 462204 -7482
rect 479604 -5986 480204 6000
rect 486804 5952 486832 6016
rect 486896 5952 486912 6016
rect 486976 5952 486992 6016
rect 487056 5952 487072 6016
rect 487136 5952 487152 6016
rect 487216 5952 487232 6016
rect 487296 5952 487312 6016
rect 487376 5952 487404 6016
rect 486804 4928 487404 5952
rect 486804 4864 486832 4928
rect 486896 4864 486912 4928
rect 486976 4864 486992 4928
rect 487056 4864 487072 4928
rect 487136 4864 487152 4928
rect 487216 4864 487232 4928
rect 487296 4864 487312 4928
rect 487376 4864 487404 4928
rect 486804 3840 487404 4864
rect 486804 3776 486832 3840
rect 486896 3776 486912 3840
rect 486976 3776 486992 3840
rect 487056 3776 487072 3840
rect 487136 3776 487152 3840
rect 487216 3776 487232 3840
rect 487296 3776 487312 3840
rect 487376 3776 487404 3840
rect 486804 2752 487404 3776
rect 486804 2688 486832 2752
rect 486896 2688 486912 2752
rect 486976 2688 486992 2752
rect 487056 2688 487072 2752
rect 487136 2688 487152 2752
rect 487216 2688 487232 2752
rect 487296 2688 487312 2752
rect 487376 2688 487404 2752
rect 486804 -1286 487404 2688
rect 486804 -1522 486986 -1286
rect 487222 -1522 487404 -1286
rect 486804 -1606 487404 -1522
rect 486804 -1842 486986 -1606
rect 487222 -1842 487404 -1606
rect 486804 -1864 487404 -1842
rect 490404 -3166 491004 6000
rect 490404 -3402 490586 -3166
rect 490822 -3402 491004 -3166
rect 490404 -3486 491004 -3402
rect 490404 -3722 490586 -3486
rect 490822 -3722 491004 -3486
rect 490404 -3744 491004 -3722
rect 494004 -5046 494604 6000
rect 494004 -5282 494186 -5046
rect 494422 -5282 494604 -5046
rect 494004 -5366 494604 -5282
rect 494004 -5602 494186 -5366
rect 494422 -5602 494604 -5366
rect 494004 -5624 494604 -5602
rect 479604 -6222 479786 -5986
rect 480022 -6222 480204 -5986
rect 479604 -6306 480204 -6222
rect 479604 -6542 479786 -6306
rect 480022 -6542 480204 -6306
rect 479604 -7504 480204 -6542
rect 497604 -6926 498204 6000
rect 504804 5472 505404 6048
rect 522804 6016 523404 6048
rect 504804 5408 504832 5472
rect 504896 5408 504912 5472
rect 504976 5408 504992 5472
rect 505056 5408 505072 5472
rect 505136 5408 505152 5472
rect 505216 5408 505232 5472
rect 505296 5408 505312 5472
rect 505376 5408 505404 5472
rect 504804 4384 505404 5408
rect 504804 4320 504832 4384
rect 504896 4320 504912 4384
rect 504976 4320 504992 4384
rect 505056 4320 505072 4384
rect 505136 4320 505152 4384
rect 505216 4320 505232 4384
rect 505296 4320 505312 4384
rect 505376 4320 505404 4384
rect 504804 3296 505404 4320
rect 504804 3232 504832 3296
rect 504896 3232 504912 3296
rect 504976 3232 504992 3296
rect 505056 3232 505072 3296
rect 505136 3232 505152 3296
rect 505216 3232 505232 3296
rect 505296 3232 505312 3296
rect 505376 3232 505404 3296
rect 504804 2406 505404 3232
rect 504804 2208 504986 2406
rect 505222 2208 505404 2406
rect 504804 2144 504832 2208
rect 504896 2144 504912 2208
rect 504976 2170 504986 2208
rect 505222 2170 505232 2208
rect 504976 2144 504992 2170
rect 505056 2144 505072 2170
rect 505136 2144 505152 2170
rect 505216 2144 505232 2170
rect 505296 2144 505312 2208
rect 505376 2144 505404 2208
rect 504804 2086 505404 2144
rect 504804 1850 504986 2086
rect 505222 1850 505404 2086
rect 504804 -346 505404 1850
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1864 505404 -902
rect 508404 -2226 509004 6000
rect 508404 -2462 508586 -2226
rect 508822 -2462 509004 -2226
rect 508404 -2546 509004 -2462
rect 508404 -2782 508586 -2546
rect 508822 -2782 509004 -2546
rect 508404 -3744 509004 -2782
rect 512004 -4106 512604 6000
rect 512004 -4342 512186 -4106
rect 512422 -4342 512604 -4106
rect 512004 -4426 512604 -4342
rect 512004 -4662 512186 -4426
rect 512422 -4662 512604 -4426
rect 512004 -5624 512604 -4662
rect 497604 -7162 497786 -6926
rect 498022 -7162 498204 -6926
rect 497604 -7246 498204 -7162
rect 497604 -7482 497786 -7246
rect 498022 -7482 498204 -7246
rect 497604 -7504 498204 -7482
rect 515604 -5986 516204 6000
rect 522804 5952 522832 6016
rect 522896 5952 522912 6016
rect 522976 5952 522992 6016
rect 523056 5952 523072 6016
rect 523136 5952 523152 6016
rect 523216 5952 523232 6016
rect 523296 5952 523312 6016
rect 523376 5952 523404 6016
rect 522804 4928 523404 5952
rect 522804 4864 522832 4928
rect 522896 4864 522912 4928
rect 522976 4864 522992 4928
rect 523056 4864 523072 4928
rect 523136 4864 523152 4928
rect 523216 4864 523232 4928
rect 523296 4864 523312 4928
rect 523376 4864 523404 4928
rect 522804 3840 523404 4864
rect 522804 3776 522832 3840
rect 522896 3776 522912 3840
rect 522976 3776 522992 3840
rect 523056 3776 523072 3840
rect 523136 3776 523152 3840
rect 523216 3776 523232 3840
rect 523296 3776 523312 3840
rect 523376 3776 523404 3840
rect 522804 2752 523404 3776
rect 522804 2688 522832 2752
rect 522896 2688 522912 2752
rect 522976 2688 522992 2752
rect 523056 2688 523072 2752
rect 523136 2688 523152 2752
rect 523216 2688 523232 2752
rect 523296 2688 523312 2752
rect 523376 2688 523404 2752
rect 522804 -1286 523404 2688
rect 522804 -1522 522986 -1286
rect 523222 -1522 523404 -1286
rect 522804 -1606 523404 -1522
rect 522804 -1842 522986 -1606
rect 523222 -1842 523404 -1606
rect 522804 -1864 523404 -1842
rect 526404 -3166 527004 6000
rect 526404 -3402 526586 -3166
rect 526822 -3402 527004 -3166
rect 526404 -3486 527004 -3402
rect 526404 -3722 526586 -3486
rect 526822 -3722 527004 -3486
rect 526404 -3744 527004 -3722
rect 530004 -5046 530604 6000
rect 530004 -5282 530186 -5046
rect 530422 -5282 530604 -5046
rect 530004 -5366 530604 -5282
rect 530004 -5602 530186 -5366
rect 530422 -5602 530604 -5366
rect 530004 -5624 530604 -5602
rect 515604 -6222 515786 -5986
rect 516022 -6222 516204 -5986
rect 515604 -6306 516204 -6222
rect 515604 -6542 515786 -6306
rect 516022 -6542 516204 -6306
rect 515604 -7504 516204 -6542
rect 533604 -6926 534204 6000
rect 540804 5472 541404 6048
rect 558804 6016 559404 6048
rect 540804 5408 540832 5472
rect 540896 5408 540912 5472
rect 540976 5408 540992 5472
rect 541056 5408 541072 5472
rect 541136 5408 541152 5472
rect 541216 5408 541232 5472
rect 541296 5408 541312 5472
rect 541376 5408 541404 5472
rect 540804 4384 541404 5408
rect 540804 4320 540832 4384
rect 540896 4320 540912 4384
rect 540976 4320 540992 4384
rect 541056 4320 541072 4384
rect 541136 4320 541152 4384
rect 541216 4320 541232 4384
rect 541296 4320 541312 4384
rect 541376 4320 541404 4384
rect 540804 3296 541404 4320
rect 540804 3232 540832 3296
rect 540896 3232 540912 3296
rect 540976 3232 540992 3296
rect 541056 3232 541072 3296
rect 541136 3232 541152 3296
rect 541216 3232 541232 3296
rect 541296 3232 541312 3296
rect 541376 3232 541404 3296
rect 540804 2406 541404 3232
rect 540804 2208 540986 2406
rect 541222 2208 541404 2406
rect 540804 2144 540832 2208
rect 540896 2144 540912 2208
rect 540976 2170 540986 2208
rect 541222 2170 541232 2208
rect 540976 2144 540992 2170
rect 541056 2144 541072 2170
rect 541136 2144 541152 2170
rect 541216 2144 541232 2170
rect 541296 2144 541312 2208
rect 541376 2144 541404 2208
rect 540804 2086 541404 2144
rect 540804 1850 540986 2086
rect 541222 1850 541404 2086
rect 540804 -346 541404 1850
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1864 541404 -902
rect 544404 -2226 545004 6000
rect 544404 -2462 544586 -2226
rect 544822 -2462 545004 -2226
rect 544404 -2546 545004 -2462
rect 544404 -2782 544586 -2546
rect 544822 -2782 545004 -2546
rect 544404 -3744 545004 -2782
rect 548004 -4106 548604 6000
rect 548004 -4342 548186 -4106
rect 548422 -4342 548604 -4106
rect 548004 -4426 548604 -4342
rect 548004 -4662 548186 -4426
rect 548422 -4662 548604 -4426
rect 548004 -5624 548604 -4662
rect 533604 -7162 533786 -6926
rect 534022 -7162 534204 -6926
rect 533604 -7246 534204 -7162
rect 533604 -7482 533786 -7246
rect 534022 -7482 534204 -7246
rect 533604 -7504 534204 -7482
rect 551604 -5986 552204 6000
rect 558804 5952 558832 6016
rect 558896 5952 558912 6016
rect 558976 5952 558992 6016
rect 559056 5952 559072 6016
rect 559136 5952 559152 6016
rect 559216 5952 559232 6016
rect 559296 5952 559312 6016
rect 559376 5952 559404 6016
rect 558804 4928 559404 5952
rect 558804 4864 558832 4928
rect 558896 4864 558912 4928
rect 558976 4864 558992 4928
rect 559056 4864 559072 4928
rect 559136 4864 559152 4928
rect 559216 4864 559232 4928
rect 559296 4864 559312 4928
rect 559376 4864 559404 4928
rect 558804 3840 559404 4864
rect 558804 3776 558832 3840
rect 558896 3776 558912 3840
rect 558976 3776 558992 3840
rect 559056 3776 559072 3840
rect 559136 3776 559152 3840
rect 559216 3776 559232 3840
rect 559296 3776 559312 3840
rect 559376 3776 559404 3840
rect 558804 2752 559404 3776
rect 558804 2688 558832 2752
rect 558896 2688 558912 2752
rect 558976 2688 558992 2752
rect 559056 2688 559072 2752
rect 559136 2688 559152 2752
rect 559216 2688 559232 2752
rect 559296 2688 559312 2752
rect 559376 2688 559404 2752
rect 558804 -1286 559404 2688
rect 558804 -1522 558986 -1286
rect 559222 -1522 559404 -1286
rect 558804 -1606 559404 -1522
rect 558804 -1842 558986 -1606
rect 559222 -1842 559404 -1606
rect 558804 -1864 559404 -1842
rect 562404 -3166 563004 6000
rect 562404 -3402 562586 -3166
rect 562822 -3402 563004 -3166
rect 562404 -3486 563004 -3402
rect 562404 -3722 562586 -3486
rect 562822 -3722 563004 -3486
rect 562404 -3744 563004 -3722
rect 566004 -5046 566604 6000
rect 566004 -5282 566186 -5046
rect 566422 -5282 566604 -5046
rect 566004 -5366 566604 -5282
rect 566004 -5602 566186 -5366
rect 566422 -5602 566604 -5366
rect 566004 -5624 566604 -5602
rect 551604 -6222 551786 -5986
rect 552022 -6222 552204 -5986
rect 551604 -6306 552204 -6222
rect 551604 -6542 551786 -6306
rect 552022 -6542 552204 -6306
rect 551604 -7504 552204 -6542
rect 569604 -6926 570204 6000
rect 576804 5472 577404 6048
rect 576804 5408 576832 5472
rect 576896 5408 576912 5472
rect 576976 5408 576992 5472
rect 577056 5408 577072 5472
rect 577136 5408 577152 5472
rect 577216 5408 577232 5472
rect 577296 5408 577312 5472
rect 577376 5408 577404 5472
rect 576804 4384 577404 5408
rect 576804 4320 576832 4384
rect 576896 4320 576912 4384
rect 576976 4320 576992 4384
rect 577056 4320 577072 4384
rect 577136 4320 577152 4384
rect 577216 4320 577232 4384
rect 577296 4320 577312 4384
rect 577376 4320 577404 4384
rect 576804 3296 577404 4320
rect 576804 3232 576832 3296
rect 576896 3232 576912 3296
rect 576976 3232 576992 3296
rect 577056 3232 577072 3296
rect 577136 3232 577152 3296
rect 577216 3232 577232 3296
rect 577296 3232 577312 3296
rect 577376 3232 577404 3296
rect 576804 2406 577404 3232
rect 576804 2208 576986 2406
rect 577222 2208 577404 2406
rect 576804 2144 576832 2208
rect 576896 2144 576912 2208
rect 576976 2170 576986 2208
rect 577222 2170 577232 2208
rect 576976 2144 576992 2170
rect 577056 2144 577072 2170
rect 577136 2144 577152 2170
rect 577216 2144 577232 2170
rect 577296 2144 577312 2208
rect 577376 2144 577404 2208
rect 576804 2086 577404 2144
rect 576804 1850 576986 2086
rect 577222 1850 577404 2086
rect 576804 -346 577404 1850
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1864 577404 -902
rect 580404 5818 580586 6054
rect 580822 5818 581004 6054
rect 580404 5734 581004 5818
rect 580404 5498 580586 5734
rect 580822 5498 581004 5734
rect 580404 -2226 581004 5498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686406 585920 704282
rect 585320 686170 585502 686406
rect 585738 686170 585920 686406
rect 585320 686086 585920 686170
rect 585320 685850 585502 686086
rect 585738 685850 585920 686086
rect 585320 650406 585920 685850
rect 585320 650170 585502 650406
rect 585738 650170 585920 650406
rect 585320 650086 585920 650170
rect 585320 649850 585502 650086
rect 585738 649850 585920 650086
rect 585320 614406 585920 649850
rect 585320 614170 585502 614406
rect 585738 614170 585920 614406
rect 585320 614086 585920 614170
rect 585320 613850 585502 614086
rect 585738 613850 585920 614086
rect 585320 578406 585920 613850
rect 585320 578170 585502 578406
rect 585738 578170 585920 578406
rect 585320 578086 585920 578170
rect 585320 577850 585502 578086
rect 585738 577850 585920 578086
rect 585320 542406 585920 577850
rect 585320 542170 585502 542406
rect 585738 542170 585920 542406
rect 585320 542086 585920 542170
rect 585320 541850 585502 542086
rect 585738 541850 585920 542086
rect 585320 506406 585920 541850
rect 585320 506170 585502 506406
rect 585738 506170 585920 506406
rect 585320 506086 585920 506170
rect 585320 505850 585502 506086
rect 585738 505850 585920 506086
rect 585320 470406 585920 505850
rect 585320 470170 585502 470406
rect 585738 470170 585920 470406
rect 585320 470086 585920 470170
rect 585320 469850 585502 470086
rect 585738 469850 585920 470086
rect 585320 434406 585920 469850
rect 585320 434170 585502 434406
rect 585738 434170 585920 434406
rect 585320 434086 585920 434170
rect 585320 433850 585502 434086
rect 585738 433850 585920 434086
rect 585320 398406 585920 433850
rect 585320 398170 585502 398406
rect 585738 398170 585920 398406
rect 585320 398086 585920 398170
rect 585320 397850 585502 398086
rect 585738 397850 585920 398086
rect 585320 362406 585920 397850
rect 585320 362170 585502 362406
rect 585738 362170 585920 362406
rect 585320 362086 585920 362170
rect 585320 361850 585502 362086
rect 585738 361850 585920 362086
rect 585320 326406 585920 361850
rect 585320 326170 585502 326406
rect 585738 326170 585920 326406
rect 585320 326086 585920 326170
rect 585320 325850 585502 326086
rect 585738 325850 585920 326086
rect 585320 290406 585920 325850
rect 585320 290170 585502 290406
rect 585738 290170 585920 290406
rect 585320 290086 585920 290170
rect 585320 289850 585502 290086
rect 585738 289850 585920 290086
rect 585320 254406 585920 289850
rect 585320 254170 585502 254406
rect 585738 254170 585920 254406
rect 585320 254086 585920 254170
rect 585320 253850 585502 254086
rect 585738 253850 585920 254086
rect 585320 218406 585920 253850
rect 585320 218170 585502 218406
rect 585738 218170 585920 218406
rect 585320 218086 585920 218170
rect 585320 217850 585502 218086
rect 585738 217850 585920 218086
rect 585320 182406 585920 217850
rect 585320 182170 585502 182406
rect 585738 182170 585920 182406
rect 585320 182086 585920 182170
rect 585320 181850 585502 182086
rect 585738 181850 585920 182086
rect 585320 146406 585920 181850
rect 585320 146170 585502 146406
rect 585738 146170 585920 146406
rect 585320 146086 585920 146170
rect 585320 145850 585502 146086
rect 585738 145850 585920 146086
rect 585320 110406 585920 145850
rect 585320 110170 585502 110406
rect 585738 110170 585920 110406
rect 585320 110086 585920 110170
rect 585320 109850 585502 110086
rect 585738 109850 585920 110086
rect 585320 74406 585920 109850
rect 585320 74170 585502 74406
rect 585738 74170 585920 74406
rect 585320 74086 585920 74170
rect 585320 73850 585502 74086
rect 585738 73850 585920 74086
rect 585320 38406 585920 73850
rect 585320 38170 585502 38406
rect 585738 38170 585920 38406
rect 585320 38086 585920 38170
rect 585320 37850 585502 38086
rect 585738 37850 585920 38086
rect 585320 2406 585920 37850
rect 585320 2170 585502 2406
rect 585738 2170 585920 2406
rect 585320 2086 585920 2170
rect 585320 1850 585502 2086
rect 585738 1850 585920 2086
rect 585320 -346 585920 1850
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586260 668406 586860 705222
rect 586260 668170 586442 668406
rect 586678 668170 586860 668406
rect 586260 668086 586860 668170
rect 586260 667850 586442 668086
rect 586678 667850 586860 668086
rect 586260 632406 586860 667850
rect 586260 632170 586442 632406
rect 586678 632170 586860 632406
rect 586260 632086 586860 632170
rect 586260 631850 586442 632086
rect 586678 631850 586860 632086
rect 586260 596406 586860 631850
rect 586260 596170 586442 596406
rect 586678 596170 586860 596406
rect 586260 596086 586860 596170
rect 586260 595850 586442 596086
rect 586678 595850 586860 596086
rect 586260 560406 586860 595850
rect 586260 560170 586442 560406
rect 586678 560170 586860 560406
rect 586260 560086 586860 560170
rect 586260 559850 586442 560086
rect 586678 559850 586860 560086
rect 586260 524406 586860 559850
rect 586260 524170 586442 524406
rect 586678 524170 586860 524406
rect 586260 524086 586860 524170
rect 586260 523850 586442 524086
rect 586678 523850 586860 524086
rect 586260 488406 586860 523850
rect 586260 488170 586442 488406
rect 586678 488170 586860 488406
rect 586260 488086 586860 488170
rect 586260 487850 586442 488086
rect 586678 487850 586860 488086
rect 586260 452406 586860 487850
rect 586260 452170 586442 452406
rect 586678 452170 586860 452406
rect 586260 452086 586860 452170
rect 586260 451850 586442 452086
rect 586678 451850 586860 452086
rect 586260 416406 586860 451850
rect 586260 416170 586442 416406
rect 586678 416170 586860 416406
rect 586260 416086 586860 416170
rect 586260 415850 586442 416086
rect 586678 415850 586860 416086
rect 586260 380406 586860 415850
rect 586260 380170 586442 380406
rect 586678 380170 586860 380406
rect 586260 380086 586860 380170
rect 586260 379850 586442 380086
rect 586678 379850 586860 380086
rect 586260 344406 586860 379850
rect 586260 344170 586442 344406
rect 586678 344170 586860 344406
rect 586260 344086 586860 344170
rect 586260 343850 586442 344086
rect 586678 343850 586860 344086
rect 586260 308406 586860 343850
rect 586260 308170 586442 308406
rect 586678 308170 586860 308406
rect 586260 308086 586860 308170
rect 586260 307850 586442 308086
rect 586678 307850 586860 308086
rect 586260 272406 586860 307850
rect 586260 272170 586442 272406
rect 586678 272170 586860 272406
rect 586260 272086 586860 272170
rect 586260 271850 586442 272086
rect 586678 271850 586860 272086
rect 586260 236406 586860 271850
rect 586260 236170 586442 236406
rect 586678 236170 586860 236406
rect 586260 236086 586860 236170
rect 586260 235850 586442 236086
rect 586678 235850 586860 236086
rect 586260 200406 586860 235850
rect 586260 200170 586442 200406
rect 586678 200170 586860 200406
rect 586260 200086 586860 200170
rect 586260 199850 586442 200086
rect 586678 199850 586860 200086
rect 586260 164406 586860 199850
rect 586260 164170 586442 164406
rect 586678 164170 586860 164406
rect 586260 164086 586860 164170
rect 586260 163850 586442 164086
rect 586678 163850 586860 164086
rect 586260 128406 586860 163850
rect 586260 128170 586442 128406
rect 586678 128170 586860 128406
rect 586260 128086 586860 128170
rect 586260 127850 586442 128086
rect 586678 127850 586860 128086
rect 586260 92406 586860 127850
rect 586260 92170 586442 92406
rect 586678 92170 586860 92406
rect 586260 92086 586860 92170
rect 586260 91850 586442 92086
rect 586678 91850 586860 92086
rect 586260 56406 586860 91850
rect 586260 56170 586442 56406
rect 586678 56170 586860 56406
rect 586260 56086 586860 56170
rect 586260 55850 586442 56086
rect 586678 55850 586860 56086
rect 586260 20406 586860 55850
rect 586260 20170 586442 20406
rect 586678 20170 586860 20406
rect 586260 20086 586860 20170
rect 586260 19850 586442 20086
rect 586678 19850 586860 20086
rect 586260 -1286 586860 19850
rect 586260 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect 586260 -1606 586860 -1522
rect 586260 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect 586260 -1864 586860 -1842
rect 587200 690054 587800 706162
rect 587200 689818 587382 690054
rect 587618 689818 587800 690054
rect 587200 689734 587800 689818
rect 587200 689498 587382 689734
rect 587618 689498 587800 689734
rect 587200 654054 587800 689498
rect 587200 653818 587382 654054
rect 587618 653818 587800 654054
rect 587200 653734 587800 653818
rect 587200 653498 587382 653734
rect 587618 653498 587800 653734
rect 587200 618054 587800 653498
rect 587200 617818 587382 618054
rect 587618 617818 587800 618054
rect 587200 617734 587800 617818
rect 587200 617498 587382 617734
rect 587618 617498 587800 617734
rect 587200 582054 587800 617498
rect 587200 581818 587382 582054
rect 587618 581818 587800 582054
rect 587200 581734 587800 581818
rect 587200 581498 587382 581734
rect 587618 581498 587800 581734
rect 587200 546054 587800 581498
rect 587200 545818 587382 546054
rect 587618 545818 587800 546054
rect 587200 545734 587800 545818
rect 587200 545498 587382 545734
rect 587618 545498 587800 545734
rect 587200 510054 587800 545498
rect 587200 509818 587382 510054
rect 587618 509818 587800 510054
rect 587200 509734 587800 509818
rect 587200 509498 587382 509734
rect 587618 509498 587800 509734
rect 587200 474054 587800 509498
rect 587200 473818 587382 474054
rect 587618 473818 587800 474054
rect 587200 473734 587800 473818
rect 587200 473498 587382 473734
rect 587618 473498 587800 473734
rect 587200 438054 587800 473498
rect 587200 437818 587382 438054
rect 587618 437818 587800 438054
rect 587200 437734 587800 437818
rect 587200 437498 587382 437734
rect 587618 437498 587800 437734
rect 587200 402054 587800 437498
rect 587200 401818 587382 402054
rect 587618 401818 587800 402054
rect 587200 401734 587800 401818
rect 587200 401498 587382 401734
rect 587618 401498 587800 401734
rect 587200 366054 587800 401498
rect 587200 365818 587382 366054
rect 587618 365818 587800 366054
rect 587200 365734 587800 365818
rect 587200 365498 587382 365734
rect 587618 365498 587800 365734
rect 587200 330054 587800 365498
rect 587200 329818 587382 330054
rect 587618 329818 587800 330054
rect 587200 329734 587800 329818
rect 587200 329498 587382 329734
rect 587618 329498 587800 329734
rect 587200 294054 587800 329498
rect 587200 293818 587382 294054
rect 587618 293818 587800 294054
rect 587200 293734 587800 293818
rect 587200 293498 587382 293734
rect 587618 293498 587800 293734
rect 587200 258054 587800 293498
rect 587200 257818 587382 258054
rect 587618 257818 587800 258054
rect 587200 257734 587800 257818
rect 587200 257498 587382 257734
rect 587618 257498 587800 257734
rect 587200 222054 587800 257498
rect 587200 221818 587382 222054
rect 587618 221818 587800 222054
rect 587200 221734 587800 221818
rect 587200 221498 587382 221734
rect 587618 221498 587800 221734
rect 587200 186054 587800 221498
rect 587200 185818 587382 186054
rect 587618 185818 587800 186054
rect 587200 185734 587800 185818
rect 587200 185498 587382 185734
rect 587618 185498 587800 185734
rect 587200 150054 587800 185498
rect 587200 149818 587382 150054
rect 587618 149818 587800 150054
rect 587200 149734 587800 149818
rect 587200 149498 587382 149734
rect 587618 149498 587800 149734
rect 587200 114054 587800 149498
rect 587200 113818 587382 114054
rect 587618 113818 587800 114054
rect 587200 113734 587800 113818
rect 587200 113498 587382 113734
rect 587618 113498 587800 113734
rect 587200 78054 587800 113498
rect 587200 77818 587382 78054
rect 587618 77818 587800 78054
rect 587200 77734 587800 77818
rect 587200 77498 587382 77734
rect 587618 77498 587800 77734
rect 587200 42054 587800 77498
rect 587200 41818 587382 42054
rect 587618 41818 587800 42054
rect 587200 41734 587800 41818
rect 587200 41498 587382 41734
rect 587618 41498 587800 41734
rect 587200 6054 587800 41498
rect 587200 5818 587382 6054
rect 587618 5818 587800 6054
rect 587200 5734 587800 5818
rect 587200 5498 587382 5734
rect 587618 5498 587800 5734
rect 580404 -2462 580586 -2226
rect 580822 -2462 581004 -2226
rect 580404 -2546 581004 -2462
rect 580404 -2782 580586 -2546
rect 580822 -2782 581004 -2546
rect 580404 -3744 581004 -2782
rect 587200 -2226 587800 5498
rect 587200 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect 587200 -2546 587800 -2462
rect 587200 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect 587200 -2804 587800 -2782
rect 588140 672054 588740 707102
rect 588140 671818 588322 672054
rect 588558 671818 588740 672054
rect 588140 671734 588740 671818
rect 588140 671498 588322 671734
rect 588558 671498 588740 671734
rect 588140 636054 588740 671498
rect 588140 635818 588322 636054
rect 588558 635818 588740 636054
rect 588140 635734 588740 635818
rect 588140 635498 588322 635734
rect 588558 635498 588740 635734
rect 588140 600054 588740 635498
rect 588140 599818 588322 600054
rect 588558 599818 588740 600054
rect 588140 599734 588740 599818
rect 588140 599498 588322 599734
rect 588558 599498 588740 599734
rect 588140 564054 588740 599498
rect 588140 563818 588322 564054
rect 588558 563818 588740 564054
rect 588140 563734 588740 563818
rect 588140 563498 588322 563734
rect 588558 563498 588740 563734
rect 588140 528054 588740 563498
rect 588140 527818 588322 528054
rect 588558 527818 588740 528054
rect 588140 527734 588740 527818
rect 588140 527498 588322 527734
rect 588558 527498 588740 527734
rect 588140 492054 588740 527498
rect 588140 491818 588322 492054
rect 588558 491818 588740 492054
rect 588140 491734 588740 491818
rect 588140 491498 588322 491734
rect 588558 491498 588740 491734
rect 588140 456054 588740 491498
rect 588140 455818 588322 456054
rect 588558 455818 588740 456054
rect 588140 455734 588740 455818
rect 588140 455498 588322 455734
rect 588558 455498 588740 455734
rect 588140 420054 588740 455498
rect 588140 419818 588322 420054
rect 588558 419818 588740 420054
rect 588140 419734 588740 419818
rect 588140 419498 588322 419734
rect 588558 419498 588740 419734
rect 588140 384054 588740 419498
rect 588140 383818 588322 384054
rect 588558 383818 588740 384054
rect 588140 383734 588740 383818
rect 588140 383498 588322 383734
rect 588558 383498 588740 383734
rect 588140 348054 588740 383498
rect 588140 347818 588322 348054
rect 588558 347818 588740 348054
rect 588140 347734 588740 347818
rect 588140 347498 588322 347734
rect 588558 347498 588740 347734
rect 588140 312054 588740 347498
rect 588140 311818 588322 312054
rect 588558 311818 588740 312054
rect 588140 311734 588740 311818
rect 588140 311498 588322 311734
rect 588558 311498 588740 311734
rect 588140 276054 588740 311498
rect 588140 275818 588322 276054
rect 588558 275818 588740 276054
rect 588140 275734 588740 275818
rect 588140 275498 588322 275734
rect 588558 275498 588740 275734
rect 588140 240054 588740 275498
rect 588140 239818 588322 240054
rect 588558 239818 588740 240054
rect 588140 239734 588740 239818
rect 588140 239498 588322 239734
rect 588558 239498 588740 239734
rect 588140 204054 588740 239498
rect 588140 203818 588322 204054
rect 588558 203818 588740 204054
rect 588140 203734 588740 203818
rect 588140 203498 588322 203734
rect 588558 203498 588740 203734
rect 588140 168054 588740 203498
rect 588140 167818 588322 168054
rect 588558 167818 588740 168054
rect 588140 167734 588740 167818
rect 588140 167498 588322 167734
rect 588558 167498 588740 167734
rect 588140 132054 588740 167498
rect 588140 131818 588322 132054
rect 588558 131818 588740 132054
rect 588140 131734 588740 131818
rect 588140 131498 588322 131734
rect 588558 131498 588740 131734
rect 588140 96054 588740 131498
rect 588140 95818 588322 96054
rect 588558 95818 588740 96054
rect 588140 95734 588740 95818
rect 588140 95498 588322 95734
rect 588558 95498 588740 95734
rect 588140 60054 588740 95498
rect 588140 59818 588322 60054
rect 588558 59818 588740 60054
rect 588140 59734 588740 59818
rect 588140 59498 588322 59734
rect 588558 59498 588740 59734
rect 588140 24054 588740 59498
rect 588140 23818 588322 24054
rect 588558 23818 588740 24054
rect 588140 23734 588740 23818
rect 588140 23498 588322 23734
rect 588558 23498 588740 23734
rect 588140 -3166 588740 23498
rect 588140 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect 588140 -3486 588740 -3402
rect 588140 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect 588140 -3744 588740 -3722
rect 589080 693654 589680 708042
rect 589080 693418 589262 693654
rect 589498 693418 589680 693654
rect 589080 693334 589680 693418
rect 589080 693098 589262 693334
rect 589498 693098 589680 693334
rect 589080 657654 589680 693098
rect 589080 657418 589262 657654
rect 589498 657418 589680 657654
rect 589080 657334 589680 657418
rect 589080 657098 589262 657334
rect 589498 657098 589680 657334
rect 589080 621654 589680 657098
rect 589080 621418 589262 621654
rect 589498 621418 589680 621654
rect 589080 621334 589680 621418
rect 589080 621098 589262 621334
rect 589498 621098 589680 621334
rect 589080 585654 589680 621098
rect 589080 585418 589262 585654
rect 589498 585418 589680 585654
rect 589080 585334 589680 585418
rect 589080 585098 589262 585334
rect 589498 585098 589680 585334
rect 589080 549654 589680 585098
rect 589080 549418 589262 549654
rect 589498 549418 589680 549654
rect 589080 549334 589680 549418
rect 589080 549098 589262 549334
rect 589498 549098 589680 549334
rect 589080 513654 589680 549098
rect 589080 513418 589262 513654
rect 589498 513418 589680 513654
rect 589080 513334 589680 513418
rect 589080 513098 589262 513334
rect 589498 513098 589680 513334
rect 589080 477654 589680 513098
rect 589080 477418 589262 477654
rect 589498 477418 589680 477654
rect 589080 477334 589680 477418
rect 589080 477098 589262 477334
rect 589498 477098 589680 477334
rect 589080 441654 589680 477098
rect 589080 441418 589262 441654
rect 589498 441418 589680 441654
rect 589080 441334 589680 441418
rect 589080 441098 589262 441334
rect 589498 441098 589680 441334
rect 589080 405654 589680 441098
rect 589080 405418 589262 405654
rect 589498 405418 589680 405654
rect 589080 405334 589680 405418
rect 589080 405098 589262 405334
rect 589498 405098 589680 405334
rect 589080 369654 589680 405098
rect 589080 369418 589262 369654
rect 589498 369418 589680 369654
rect 589080 369334 589680 369418
rect 589080 369098 589262 369334
rect 589498 369098 589680 369334
rect 589080 333654 589680 369098
rect 589080 333418 589262 333654
rect 589498 333418 589680 333654
rect 589080 333334 589680 333418
rect 589080 333098 589262 333334
rect 589498 333098 589680 333334
rect 589080 297654 589680 333098
rect 589080 297418 589262 297654
rect 589498 297418 589680 297654
rect 589080 297334 589680 297418
rect 589080 297098 589262 297334
rect 589498 297098 589680 297334
rect 589080 261654 589680 297098
rect 589080 261418 589262 261654
rect 589498 261418 589680 261654
rect 589080 261334 589680 261418
rect 589080 261098 589262 261334
rect 589498 261098 589680 261334
rect 589080 225654 589680 261098
rect 589080 225418 589262 225654
rect 589498 225418 589680 225654
rect 589080 225334 589680 225418
rect 589080 225098 589262 225334
rect 589498 225098 589680 225334
rect 589080 189654 589680 225098
rect 589080 189418 589262 189654
rect 589498 189418 589680 189654
rect 589080 189334 589680 189418
rect 589080 189098 589262 189334
rect 589498 189098 589680 189334
rect 589080 153654 589680 189098
rect 589080 153418 589262 153654
rect 589498 153418 589680 153654
rect 589080 153334 589680 153418
rect 589080 153098 589262 153334
rect 589498 153098 589680 153334
rect 589080 117654 589680 153098
rect 589080 117418 589262 117654
rect 589498 117418 589680 117654
rect 589080 117334 589680 117418
rect 589080 117098 589262 117334
rect 589498 117098 589680 117334
rect 589080 81654 589680 117098
rect 589080 81418 589262 81654
rect 589498 81418 589680 81654
rect 589080 81334 589680 81418
rect 589080 81098 589262 81334
rect 589498 81098 589680 81334
rect 589080 45654 589680 81098
rect 589080 45418 589262 45654
rect 589498 45418 589680 45654
rect 589080 45334 589680 45418
rect 589080 45098 589262 45334
rect 589498 45098 589680 45334
rect 589080 9654 589680 45098
rect 589080 9418 589262 9654
rect 589498 9418 589680 9654
rect 589080 9334 589680 9418
rect 589080 9098 589262 9334
rect 589498 9098 589680 9334
rect 589080 -4106 589680 9098
rect 589080 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect 589080 -4426 589680 -4342
rect 589080 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect 589080 -4684 589680 -4662
rect 590020 675654 590620 708982
rect 590020 675418 590202 675654
rect 590438 675418 590620 675654
rect 590020 675334 590620 675418
rect 590020 675098 590202 675334
rect 590438 675098 590620 675334
rect 590020 639654 590620 675098
rect 590020 639418 590202 639654
rect 590438 639418 590620 639654
rect 590020 639334 590620 639418
rect 590020 639098 590202 639334
rect 590438 639098 590620 639334
rect 590020 603654 590620 639098
rect 590020 603418 590202 603654
rect 590438 603418 590620 603654
rect 590020 603334 590620 603418
rect 590020 603098 590202 603334
rect 590438 603098 590620 603334
rect 590020 567654 590620 603098
rect 590020 567418 590202 567654
rect 590438 567418 590620 567654
rect 590020 567334 590620 567418
rect 590020 567098 590202 567334
rect 590438 567098 590620 567334
rect 590020 531654 590620 567098
rect 590020 531418 590202 531654
rect 590438 531418 590620 531654
rect 590020 531334 590620 531418
rect 590020 531098 590202 531334
rect 590438 531098 590620 531334
rect 590020 495654 590620 531098
rect 590020 495418 590202 495654
rect 590438 495418 590620 495654
rect 590020 495334 590620 495418
rect 590020 495098 590202 495334
rect 590438 495098 590620 495334
rect 590020 459654 590620 495098
rect 590020 459418 590202 459654
rect 590438 459418 590620 459654
rect 590020 459334 590620 459418
rect 590020 459098 590202 459334
rect 590438 459098 590620 459334
rect 590020 423654 590620 459098
rect 590020 423418 590202 423654
rect 590438 423418 590620 423654
rect 590020 423334 590620 423418
rect 590020 423098 590202 423334
rect 590438 423098 590620 423334
rect 590020 387654 590620 423098
rect 590020 387418 590202 387654
rect 590438 387418 590620 387654
rect 590020 387334 590620 387418
rect 590020 387098 590202 387334
rect 590438 387098 590620 387334
rect 590020 351654 590620 387098
rect 590020 351418 590202 351654
rect 590438 351418 590620 351654
rect 590020 351334 590620 351418
rect 590020 351098 590202 351334
rect 590438 351098 590620 351334
rect 590020 315654 590620 351098
rect 590020 315418 590202 315654
rect 590438 315418 590620 315654
rect 590020 315334 590620 315418
rect 590020 315098 590202 315334
rect 590438 315098 590620 315334
rect 590020 279654 590620 315098
rect 590020 279418 590202 279654
rect 590438 279418 590620 279654
rect 590020 279334 590620 279418
rect 590020 279098 590202 279334
rect 590438 279098 590620 279334
rect 590020 243654 590620 279098
rect 590020 243418 590202 243654
rect 590438 243418 590620 243654
rect 590020 243334 590620 243418
rect 590020 243098 590202 243334
rect 590438 243098 590620 243334
rect 590020 207654 590620 243098
rect 590020 207418 590202 207654
rect 590438 207418 590620 207654
rect 590020 207334 590620 207418
rect 590020 207098 590202 207334
rect 590438 207098 590620 207334
rect 590020 171654 590620 207098
rect 590020 171418 590202 171654
rect 590438 171418 590620 171654
rect 590020 171334 590620 171418
rect 590020 171098 590202 171334
rect 590438 171098 590620 171334
rect 590020 135654 590620 171098
rect 590020 135418 590202 135654
rect 590438 135418 590620 135654
rect 590020 135334 590620 135418
rect 590020 135098 590202 135334
rect 590438 135098 590620 135334
rect 590020 99654 590620 135098
rect 590020 99418 590202 99654
rect 590438 99418 590620 99654
rect 590020 99334 590620 99418
rect 590020 99098 590202 99334
rect 590438 99098 590620 99334
rect 590020 63654 590620 99098
rect 590020 63418 590202 63654
rect 590438 63418 590620 63654
rect 590020 63334 590620 63418
rect 590020 63098 590202 63334
rect 590438 63098 590620 63334
rect 590020 27654 590620 63098
rect 590020 27418 590202 27654
rect 590438 27418 590620 27654
rect 590020 27334 590620 27418
rect 590020 27098 590202 27334
rect 590438 27098 590620 27334
rect 590020 -5046 590620 27098
rect 590020 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect 590020 -5366 590620 -5282
rect 590020 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect 590020 -5624 590620 -5602
rect 590960 697254 591560 709922
rect 590960 697018 591142 697254
rect 591378 697018 591560 697254
rect 590960 696934 591560 697018
rect 590960 696698 591142 696934
rect 591378 696698 591560 696934
rect 590960 661254 591560 696698
rect 590960 661018 591142 661254
rect 591378 661018 591560 661254
rect 590960 660934 591560 661018
rect 590960 660698 591142 660934
rect 591378 660698 591560 660934
rect 590960 625254 591560 660698
rect 590960 625018 591142 625254
rect 591378 625018 591560 625254
rect 590960 624934 591560 625018
rect 590960 624698 591142 624934
rect 591378 624698 591560 624934
rect 590960 589254 591560 624698
rect 590960 589018 591142 589254
rect 591378 589018 591560 589254
rect 590960 588934 591560 589018
rect 590960 588698 591142 588934
rect 591378 588698 591560 588934
rect 590960 553254 591560 588698
rect 590960 553018 591142 553254
rect 591378 553018 591560 553254
rect 590960 552934 591560 553018
rect 590960 552698 591142 552934
rect 591378 552698 591560 552934
rect 590960 517254 591560 552698
rect 590960 517018 591142 517254
rect 591378 517018 591560 517254
rect 590960 516934 591560 517018
rect 590960 516698 591142 516934
rect 591378 516698 591560 516934
rect 590960 481254 591560 516698
rect 590960 481018 591142 481254
rect 591378 481018 591560 481254
rect 590960 480934 591560 481018
rect 590960 480698 591142 480934
rect 591378 480698 591560 480934
rect 590960 445254 591560 480698
rect 590960 445018 591142 445254
rect 591378 445018 591560 445254
rect 590960 444934 591560 445018
rect 590960 444698 591142 444934
rect 591378 444698 591560 444934
rect 590960 409254 591560 444698
rect 590960 409018 591142 409254
rect 591378 409018 591560 409254
rect 590960 408934 591560 409018
rect 590960 408698 591142 408934
rect 591378 408698 591560 408934
rect 590960 373254 591560 408698
rect 590960 373018 591142 373254
rect 591378 373018 591560 373254
rect 590960 372934 591560 373018
rect 590960 372698 591142 372934
rect 591378 372698 591560 372934
rect 590960 337254 591560 372698
rect 590960 337018 591142 337254
rect 591378 337018 591560 337254
rect 590960 336934 591560 337018
rect 590960 336698 591142 336934
rect 591378 336698 591560 336934
rect 590960 301254 591560 336698
rect 590960 301018 591142 301254
rect 591378 301018 591560 301254
rect 590960 300934 591560 301018
rect 590960 300698 591142 300934
rect 591378 300698 591560 300934
rect 590960 265254 591560 300698
rect 590960 265018 591142 265254
rect 591378 265018 591560 265254
rect 590960 264934 591560 265018
rect 590960 264698 591142 264934
rect 591378 264698 591560 264934
rect 590960 229254 591560 264698
rect 590960 229018 591142 229254
rect 591378 229018 591560 229254
rect 590960 228934 591560 229018
rect 590960 228698 591142 228934
rect 591378 228698 591560 228934
rect 590960 193254 591560 228698
rect 590960 193018 591142 193254
rect 591378 193018 591560 193254
rect 590960 192934 591560 193018
rect 590960 192698 591142 192934
rect 591378 192698 591560 192934
rect 590960 157254 591560 192698
rect 590960 157018 591142 157254
rect 591378 157018 591560 157254
rect 590960 156934 591560 157018
rect 590960 156698 591142 156934
rect 591378 156698 591560 156934
rect 590960 121254 591560 156698
rect 590960 121018 591142 121254
rect 591378 121018 591560 121254
rect 590960 120934 591560 121018
rect 590960 120698 591142 120934
rect 591378 120698 591560 120934
rect 590960 85254 591560 120698
rect 590960 85018 591142 85254
rect 591378 85018 591560 85254
rect 590960 84934 591560 85018
rect 590960 84698 591142 84934
rect 591378 84698 591560 84934
rect 590960 49254 591560 84698
rect 590960 49018 591142 49254
rect 591378 49018 591560 49254
rect 590960 48934 591560 49018
rect 590960 48698 591142 48934
rect 591378 48698 591560 48934
rect 590960 13254 591560 48698
rect 590960 13018 591142 13254
rect 591378 13018 591560 13254
rect 590960 12934 591560 13018
rect 590960 12698 591142 12934
rect 591378 12698 591560 12934
rect 590960 -5986 591560 12698
rect 590960 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect 590960 -6306 591560 -6222
rect 590960 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect 590960 -6564 591560 -6542
rect 591900 679254 592500 710862
rect 591900 679018 592082 679254
rect 592318 679018 592500 679254
rect 591900 678934 592500 679018
rect 591900 678698 592082 678934
rect 592318 678698 592500 678934
rect 591900 643254 592500 678698
rect 591900 643018 592082 643254
rect 592318 643018 592500 643254
rect 591900 642934 592500 643018
rect 591900 642698 592082 642934
rect 592318 642698 592500 642934
rect 591900 607254 592500 642698
rect 591900 607018 592082 607254
rect 592318 607018 592500 607254
rect 591900 606934 592500 607018
rect 591900 606698 592082 606934
rect 592318 606698 592500 606934
rect 591900 571254 592500 606698
rect 591900 571018 592082 571254
rect 592318 571018 592500 571254
rect 591900 570934 592500 571018
rect 591900 570698 592082 570934
rect 592318 570698 592500 570934
rect 591900 535254 592500 570698
rect 591900 535018 592082 535254
rect 592318 535018 592500 535254
rect 591900 534934 592500 535018
rect 591900 534698 592082 534934
rect 592318 534698 592500 534934
rect 591900 499254 592500 534698
rect 591900 499018 592082 499254
rect 592318 499018 592500 499254
rect 591900 498934 592500 499018
rect 591900 498698 592082 498934
rect 592318 498698 592500 498934
rect 591900 463254 592500 498698
rect 591900 463018 592082 463254
rect 592318 463018 592500 463254
rect 591900 462934 592500 463018
rect 591900 462698 592082 462934
rect 592318 462698 592500 462934
rect 591900 427254 592500 462698
rect 591900 427018 592082 427254
rect 592318 427018 592500 427254
rect 591900 426934 592500 427018
rect 591900 426698 592082 426934
rect 592318 426698 592500 426934
rect 591900 391254 592500 426698
rect 591900 391018 592082 391254
rect 592318 391018 592500 391254
rect 591900 390934 592500 391018
rect 591900 390698 592082 390934
rect 592318 390698 592500 390934
rect 591900 355254 592500 390698
rect 591900 355018 592082 355254
rect 592318 355018 592500 355254
rect 591900 354934 592500 355018
rect 591900 354698 592082 354934
rect 592318 354698 592500 354934
rect 591900 319254 592500 354698
rect 591900 319018 592082 319254
rect 592318 319018 592500 319254
rect 591900 318934 592500 319018
rect 591900 318698 592082 318934
rect 592318 318698 592500 318934
rect 591900 283254 592500 318698
rect 591900 283018 592082 283254
rect 592318 283018 592500 283254
rect 591900 282934 592500 283018
rect 591900 282698 592082 282934
rect 592318 282698 592500 282934
rect 591900 247254 592500 282698
rect 591900 247018 592082 247254
rect 592318 247018 592500 247254
rect 591900 246934 592500 247018
rect 591900 246698 592082 246934
rect 592318 246698 592500 246934
rect 591900 211254 592500 246698
rect 591900 211018 592082 211254
rect 592318 211018 592500 211254
rect 591900 210934 592500 211018
rect 591900 210698 592082 210934
rect 592318 210698 592500 210934
rect 591900 175254 592500 210698
rect 591900 175018 592082 175254
rect 592318 175018 592500 175254
rect 591900 174934 592500 175018
rect 591900 174698 592082 174934
rect 592318 174698 592500 174934
rect 591900 139254 592500 174698
rect 591900 139018 592082 139254
rect 592318 139018 592500 139254
rect 591900 138934 592500 139018
rect 591900 138698 592082 138934
rect 592318 138698 592500 138934
rect 591900 103254 592500 138698
rect 591900 103018 592082 103254
rect 592318 103018 592500 103254
rect 591900 102934 592500 103018
rect 591900 102698 592082 102934
rect 592318 102698 592500 102934
rect 591900 67254 592500 102698
rect 591900 67018 592082 67254
rect 592318 67018 592500 67254
rect 591900 66934 592500 67018
rect 591900 66698 592082 66934
rect 592318 66698 592500 66934
rect 591900 31254 592500 66698
rect 591900 31018 592082 31254
rect 592318 31018 592500 31254
rect 591900 30934 592500 31018
rect 591900 30698 592082 30934
rect 592318 30698 592500 30934
rect 569604 -7162 569786 -6926
rect 570022 -7162 570204 -6926
rect 569604 -7246 570204 -7162
rect 569604 -7482 569786 -7246
rect 570022 -7482 570204 -7246
rect 569604 -7504 570204 -7482
rect 591900 -6926 592500 30698
rect 591900 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect 591900 -7246 592500 -7162
rect 591900 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect 591900 -7504 592500 -7482
<< via4 >>
rect -8394 711182 -8158 711418
rect -8394 710862 -8158 711098
rect -8394 679018 -8158 679254
rect -8394 678698 -8158 678934
rect -8394 643018 -8158 643254
rect -8394 642698 -8158 642934
rect -8394 607018 -8158 607254
rect -8394 606698 -8158 606934
rect -8394 571018 -8158 571254
rect -8394 570698 -8158 570934
rect -8394 535018 -8158 535254
rect -8394 534698 -8158 534934
rect -8394 499018 -8158 499254
rect -8394 498698 -8158 498934
rect -8394 463018 -8158 463254
rect -8394 462698 -8158 462934
rect -8394 427018 -8158 427254
rect -8394 426698 -8158 426934
rect -8394 391018 -8158 391254
rect -8394 390698 -8158 390934
rect -8394 355018 -8158 355254
rect -8394 354698 -8158 354934
rect -8394 319018 -8158 319254
rect -8394 318698 -8158 318934
rect -8394 283018 -8158 283254
rect -8394 282698 -8158 282934
rect -8394 247018 -8158 247254
rect -8394 246698 -8158 246934
rect -8394 211018 -8158 211254
rect -8394 210698 -8158 210934
rect -8394 175018 -8158 175254
rect -8394 174698 -8158 174934
rect -8394 139018 -8158 139254
rect -8394 138698 -8158 138934
rect -8394 103018 -8158 103254
rect -8394 102698 -8158 102934
rect -8394 67018 -8158 67254
rect -8394 66698 -8158 66934
rect -8394 31018 -8158 31254
rect -8394 30698 -8158 30934
rect -7454 710242 -7218 710478
rect -7454 709922 -7218 710158
rect 11786 710242 12022 710478
rect 11786 709922 12022 710158
rect -7454 697018 -7218 697254
rect -7454 696698 -7218 696934
rect -7454 661018 -7218 661254
rect -7454 660698 -7218 660934
rect -7454 625018 -7218 625254
rect -7454 624698 -7218 624934
rect -7454 589018 -7218 589254
rect -7454 588698 -7218 588934
rect -7454 553018 -7218 553254
rect -7454 552698 -7218 552934
rect -7454 517018 -7218 517254
rect -7454 516698 -7218 516934
rect -7454 481018 -7218 481254
rect -7454 480698 -7218 480934
rect -7454 445018 -7218 445254
rect -7454 444698 -7218 444934
rect -7454 409018 -7218 409254
rect -7454 408698 -7218 408934
rect -7454 373018 -7218 373254
rect -7454 372698 -7218 372934
rect -7454 337018 -7218 337254
rect -7454 336698 -7218 336934
rect -7454 301018 -7218 301254
rect -7454 300698 -7218 300934
rect -7454 265018 -7218 265254
rect -7454 264698 -7218 264934
rect -7454 229018 -7218 229254
rect -7454 228698 -7218 228934
rect -7454 193018 -7218 193254
rect -7454 192698 -7218 192934
rect -7454 157018 -7218 157254
rect -7454 156698 -7218 156934
rect -7454 121018 -7218 121254
rect -7454 120698 -7218 120934
rect -7454 85018 -7218 85254
rect -7454 84698 -7218 84934
rect -7454 49018 -7218 49254
rect -7454 48698 -7218 48934
rect -7454 13018 -7218 13254
rect -7454 12698 -7218 12934
rect -6514 709302 -6278 709538
rect -6514 708982 -6278 709218
rect -6514 675418 -6278 675654
rect -6514 675098 -6278 675334
rect -6514 639418 -6278 639654
rect -6514 639098 -6278 639334
rect -6514 603418 -6278 603654
rect -6514 603098 -6278 603334
rect -6514 567418 -6278 567654
rect -6514 567098 -6278 567334
rect -6514 531418 -6278 531654
rect -6514 531098 -6278 531334
rect -6514 495418 -6278 495654
rect -6514 495098 -6278 495334
rect -6514 459418 -6278 459654
rect -6514 459098 -6278 459334
rect -6514 423418 -6278 423654
rect -6514 423098 -6278 423334
rect -6514 387418 -6278 387654
rect -6514 387098 -6278 387334
rect -6514 351418 -6278 351654
rect -6514 351098 -6278 351334
rect -6514 315418 -6278 315654
rect -6514 315098 -6278 315334
rect -6514 279418 -6278 279654
rect -6514 279098 -6278 279334
rect -6514 243418 -6278 243654
rect -6514 243098 -6278 243334
rect -6514 207418 -6278 207654
rect -6514 207098 -6278 207334
rect -6514 171418 -6278 171654
rect -6514 171098 -6278 171334
rect -6514 135418 -6278 135654
rect -6514 135098 -6278 135334
rect -6514 99418 -6278 99654
rect -6514 99098 -6278 99334
rect -6514 63418 -6278 63654
rect -6514 63098 -6278 63334
rect -6514 27418 -6278 27654
rect -6514 27098 -6278 27334
rect -5574 708362 -5338 708598
rect -5574 708042 -5338 708278
rect 8186 708362 8422 708598
rect 8186 708042 8422 708278
rect -5574 693418 -5338 693654
rect -5574 693098 -5338 693334
rect -5574 657418 -5338 657654
rect -5574 657098 -5338 657334
rect -5574 621418 -5338 621654
rect -5574 621098 -5338 621334
rect -5574 585418 -5338 585654
rect -5574 585098 -5338 585334
rect -5574 549418 -5338 549654
rect -5574 549098 -5338 549334
rect -5574 513418 -5338 513654
rect -5574 513098 -5338 513334
rect -5574 477418 -5338 477654
rect -5574 477098 -5338 477334
rect -5574 441418 -5338 441654
rect -5574 441098 -5338 441334
rect -5574 405418 -5338 405654
rect -5574 405098 -5338 405334
rect -5574 369418 -5338 369654
rect -5574 369098 -5338 369334
rect -5574 333418 -5338 333654
rect -5574 333098 -5338 333334
rect -5574 297418 -5338 297654
rect -5574 297098 -5338 297334
rect -5574 261418 -5338 261654
rect -5574 261098 -5338 261334
rect -5574 225418 -5338 225654
rect -5574 225098 -5338 225334
rect -5574 189418 -5338 189654
rect -5574 189098 -5338 189334
rect -5574 153418 -5338 153654
rect -5574 153098 -5338 153334
rect -5574 117418 -5338 117654
rect -5574 117098 -5338 117334
rect -5574 81418 -5338 81654
rect -5574 81098 -5338 81334
rect -5574 45418 -5338 45654
rect -5574 45098 -5338 45334
rect -5574 9418 -5338 9654
rect -5574 9098 -5338 9334
rect -4634 707422 -4398 707658
rect -4634 707102 -4398 707338
rect -4634 671818 -4398 672054
rect -4634 671498 -4398 671734
rect -4634 635818 -4398 636054
rect -4634 635498 -4398 635734
rect -4634 599818 -4398 600054
rect -4634 599498 -4398 599734
rect -4634 563818 -4398 564054
rect -4634 563498 -4398 563734
rect -4634 527818 -4398 528054
rect -4634 527498 -4398 527734
rect -4634 491818 -4398 492054
rect -4634 491498 -4398 491734
rect -4634 455818 -4398 456054
rect -4634 455498 -4398 455734
rect -4634 419818 -4398 420054
rect -4634 419498 -4398 419734
rect -4634 383818 -4398 384054
rect -4634 383498 -4398 383734
rect -4634 347818 -4398 348054
rect -4634 347498 -4398 347734
rect -4634 311818 -4398 312054
rect -4634 311498 -4398 311734
rect -4634 275818 -4398 276054
rect -4634 275498 -4398 275734
rect -4634 239818 -4398 240054
rect -4634 239498 -4398 239734
rect -4634 203818 -4398 204054
rect -4634 203498 -4398 203734
rect -4634 167818 -4398 168054
rect -4634 167498 -4398 167734
rect -4634 131818 -4398 132054
rect -4634 131498 -4398 131734
rect -4634 95818 -4398 96054
rect -4634 95498 -4398 95734
rect -4634 59818 -4398 60054
rect -4634 59498 -4398 59734
rect -4634 23818 -4398 24054
rect -4634 23498 -4398 23734
rect -3694 706482 -3458 706718
rect -3694 706162 -3458 706398
rect 4586 706482 4822 706718
rect 4586 706162 4822 706398
rect -3694 689818 -3458 690054
rect -3694 689498 -3458 689734
rect -3694 653818 -3458 654054
rect -3694 653498 -3458 653734
rect -3694 617818 -3458 618054
rect -3694 617498 -3458 617734
rect -3694 581818 -3458 582054
rect -3694 581498 -3458 581734
rect -3694 545818 -3458 546054
rect -3694 545498 -3458 545734
rect -3694 509818 -3458 510054
rect -3694 509498 -3458 509734
rect -3694 473818 -3458 474054
rect -3694 473498 -3458 473734
rect -3694 437818 -3458 438054
rect -3694 437498 -3458 437734
rect -3694 401818 -3458 402054
rect -3694 401498 -3458 401734
rect -3694 365818 -3458 366054
rect -3694 365498 -3458 365734
rect -3694 329818 -3458 330054
rect -3694 329498 -3458 329734
rect -3694 293818 -3458 294054
rect -3694 293498 -3458 293734
rect -3694 257818 -3458 258054
rect -3694 257498 -3458 257734
rect -3694 221818 -3458 222054
rect -3694 221498 -3458 221734
rect -3694 185818 -3458 186054
rect -3694 185498 -3458 185734
rect -3694 149818 -3458 150054
rect -3694 149498 -3458 149734
rect -3694 113818 -3458 114054
rect -3694 113498 -3458 113734
rect -3694 77818 -3458 78054
rect -3694 77498 -3458 77734
rect -3694 41818 -3458 42054
rect -3694 41498 -3458 41734
rect -3694 5818 -3458 6054
rect -3694 5498 -3458 5734
rect -2754 705542 -2518 705778
rect -2754 705222 -2518 705458
rect -2754 668170 -2518 668406
rect -2754 667850 -2518 668086
rect -2754 632170 -2518 632406
rect -2754 631850 -2518 632086
rect -2754 596170 -2518 596406
rect -2754 595850 -2518 596086
rect -2754 560170 -2518 560406
rect -2754 559850 -2518 560086
rect -2754 524170 -2518 524406
rect -2754 523850 -2518 524086
rect -2754 488170 -2518 488406
rect -2754 487850 -2518 488086
rect -2754 452170 -2518 452406
rect -2754 451850 -2518 452086
rect -2754 416170 -2518 416406
rect -2754 415850 -2518 416086
rect -2754 380170 -2518 380406
rect -2754 379850 -2518 380086
rect -2754 344170 -2518 344406
rect -2754 343850 -2518 344086
rect -2754 308170 -2518 308406
rect -2754 307850 -2518 308086
rect -2754 272170 -2518 272406
rect -2754 271850 -2518 272086
rect -2754 236170 -2518 236406
rect -2754 235850 -2518 236086
rect -2754 200170 -2518 200406
rect -2754 199850 -2518 200086
rect -2754 164170 -2518 164406
rect -2754 163850 -2518 164086
rect -2754 128170 -2518 128406
rect -2754 127850 -2518 128086
rect -2754 92170 -2518 92406
rect -2754 91850 -2518 92086
rect -2754 56170 -2518 56406
rect -2754 55850 -2518 56086
rect -2754 20170 -2518 20406
rect -2754 19850 -2518 20086
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686170 -1578 686406
rect -1814 685850 -1578 686086
rect -1814 650170 -1578 650406
rect -1814 649850 -1578 650086
rect -1814 614170 -1578 614406
rect -1814 613850 -1578 614086
rect -1814 578170 -1578 578406
rect -1814 577850 -1578 578086
rect -1814 542170 -1578 542406
rect -1814 541850 -1578 542086
rect -1814 506170 -1578 506406
rect -1814 505850 -1578 506086
rect -1814 470170 -1578 470406
rect -1814 469850 -1578 470086
rect -1814 434170 -1578 434406
rect -1814 433850 -1578 434086
rect -1814 398170 -1578 398406
rect -1814 397850 -1578 398086
rect -1814 362170 -1578 362406
rect -1814 361850 -1578 362086
rect -1814 326170 -1578 326406
rect -1814 325850 -1578 326086
rect -1814 290170 -1578 290406
rect -1814 289850 -1578 290086
rect -1814 254170 -1578 254406
rect -1814 253850 -1578 254086
rect -1814 218170 -1578 218406
rect -1814 217850 -1578 218086
rect -1814 182170 -1578 182406
rect -1814 181850 -1578 182086
rect -1814 146170 -1578 146406
rect -1814 145850 -1578 146086
rect -1814 110170 -1578 110406
rect -1814 109850 -1578 110086
rect -1814 74170 -1578 74406
rect -1814 73850 -1578 74086
rect -1814 38170 -1578 38406
rect -1814 37850 -1578 38086
rect -1814 2170 -1578 2406
rect -1814 1850 -1578 2086
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686170 1222 686406
rect 986 685850 1222 686086
rect 986 650170 1222 650406
rect 986 649850 1222 650086
rect 986 614170 1222 614406
rect 986 613850 1222 614086
rect 986 578170 1222 578406
rect 986 577850 1222 578086
rect 986 542170 1222 542406
rect 986 541850 1222 542086
rect 986 506170 1222 506406
rect 986 505850 1222 506086
rect 986 470170 1222 470406
rect 986 469850 1222 470086
rect 986 434170 1222 434406
rect 986 433850 1222 434086
rect 986 398170 1222 398406
rect 986 397850 1222 398086
rect 986 362170 1222 362406
rect 986 361850 1222 362086
rect 986 326170 1222 326406
rect 986 325850 1222 326086
rect 986 290170 1222 290406
rect 986 289850 1222 290086
rect 986 254170 1222 254406
rect 986 253850 1222 254086
rect 986 218170 1222 218406
rect 986 217850 1222 218086
rect 986 182170 1222 182406
rect 986 181850 1222 182086
rect 986 146170 1222 146406
rect 986 145850 1222 146086
rect 986 110170 1222 110406
rect 986 109850 1222 110086
rect 986 74170 1222 74406
rect 986 73850 1222 74086
rect 986 38170 1222 38406
rect 986 37850 1222 38086
rect 986 2170 1222 2406
rect 986 1850 1222 2086
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2754 -1522 -2518 -1286
rect -2754 -1842 -2518 -1606
rect 29786 711182 30022 711418
rect 29786 710862 30022 711098
rect 26186 709302 26422 709538
rect 26186 708982 26422 709218
rect 22586 707422 22822 707658
rect 22586 707102 22822 707338
rect 18986 705542 19222 705778
rect 18986 705222 19222 705458
rect 47786 710242 48022 710478
rect 47786 709922 48022 710158
rect 44186 708362 44422 708598
rect 44186 708042 44422 708278
rect 40586 706482 40822 706718
rect 40586 706162 40822 706398
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 65786 711182 66022 711418
rect 65786 710862 66022 711098
rect 62186 709302 62422 709538
rect 62186 708982 62422 709218
rect 58586 707422 58822 707658
rect 58586 707102 58822 707338
rect 54986 705542 55222 705778
rect 54986 705222 55222 705458
rect 83786 710242 84022 710478
rect 83786 709922 84022 710158
rect 80186 708362 80422 708598
rect 80186 708042 80422 708278
rect 76586 706482 76822 706718
rect 76586 706162 76822 706398
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 101786 711182 102022 711418
rect 101786 710862 102022 711098
rect 98186 709302 98422 709538
rect 98186 708982 98422 709218
rect 94586 707422 94822 707658
rect 94586 707102 94822 707338
rect 90986 705542 91222 705778
rect 90986 705222 91222 705458
rect 119786 710242 120022 710478
rect 119786 709922 120022 710158
rect 116186 708362 116422 708598
rect 116186 708042 116422 708278
rect 112586 706482 112822 706718
rect 112586 706162 112822 706398
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 137786 711182 138022 711418
rect 137786 710862 138022 711098
rect 134186 709302 134422 709538
rect 134186 708982 134422 709218
rect 130586 707422 130822 707658
rect 130586 707102 130822 707338
rect 126986 705542 127222 705778
rect 126986 705222 127222 705458
rect 155786 710242 156022 710478
rect 155786 709922 156022 710158
rect 152186 708362 152422 708598
rect 152186 708042 152422 708278
rect 148586 706482 148822 706718
rect 148586 706162 148822 706398
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 173786 711182 174022 711418
rect 173786 710862 174022 711098
rect 170186 709302 170422 709538
rect 170186 708982 170422 709218
rect 166586 707422 166822 707658
rect 166586 707102 166822 707338
rect 162986 705542 163222 705778
rect 162986 705222 163222 705458
rect 191786 710242 192022 710478
rect 191786 709922 192022 710158
rect 188186 708362 188422 708598
rect 188186 708042 188422 708278
rect 184586 706482 184822 706718
rect 184586 706162 184822 706398
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 209786 711182 210022 711418
rect 209786 710862 210022 711098
rect 206186 709302 206422 709538
rect 206186 708982 206422 709218
rect 202586 707422 202822 707658
rect 202586 707102 202822 707338
rect 198986 705542 199222 705778
rect 198986 705222 199222 705458
rect 227786 710242 228022 710478
rect 227786 709922 228022 710158
rect 224186 708362 224422 708598
rect 224186 708042 224422 708278
rect 220586 706482 220822 706718
rect 220586 706162 220822 706398
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 245786 711182 246022 711418
rect 245786 710862 246022 711098
rect 242186 709302 242422 709538
rect 242186 708982 242422 709218
rect 238586 707422 238822 707658
rect 238586 707102 238822 707338
rect 234986 705542 235222 705778
rect 234986 705222 235222 705458
rect 263786 710242 264022 710478
rect 263786 709922 264022 710158
rect 260186 708362 260422 708598
rect 260186 708042 260422 708278
rect 256586 706482 256822 706718
rect 256586 706162 256822 706398
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 281786 711182 282022 711418
rect 281786 710862 282022 711098
rect 278186 709302 278422 709538
rect 278186 708982 278422 709218
rect 274586 707422 274822 707658
rect 274586 707102 274822 707338
rect 270986 705542 271222 705778
rect 270986 705222 271222 705458
rect 299786 710242 300022 710478
rect 299786 709922 300022 710158
rect 296186 708362 296422 708598
rect 296186 708042 296422 708278
rect 292586 706482 292822 706718
rect 292586 706162 292822 706398
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 317786 711182 318022 711418
rect 317786 710862 318022 711098
rect 314186 709302 314422 709538
rect 314186 708982 314422 709218
rect 310586 707422 310822 707658
rect 310586 707102 310822 707338
rect 306986 705542 307222 705778
rect 306986 705222 307222 705458
rect 335786 710242 336022 710478
rect 335786 709922 336022 710158
rect 332186 708362 332422 708598
rect 332186 708042 332422 708278
rect 328586 706482 328822 706718
rect 328586 706162 328822 706398
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 353786 711182 354022 711418
rect 353786 710862 354022 711098
rect 350186 709302 350422 709538
rect 350186 708982 350422 709218
rect 346586 707422 346822 707658
rect 346586 707102 346822 707338
rect 342986 705542 343222 705778
rect 342986 705222 343222 705458
rect 371786 710242 372022 710478
rect 371786 709922 372022 710158
rect 368186 708362 368422 708598
rect 368186 708042 368422 708278
rect 364586 706482 364822 706718
rect 364586 706162 364822 706398
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 389786 711182 390022 711418
rect 389786 710862 390022 711098
rect 386186 709302 386422 709538
rect 386186 708982 386422 709218
rect 382586 707422 382822 707658
rect 382586 707102 382822 707338
rect 378986 705542 379222 705778
rect 378986 705222 379222 705458
rect 407786 710242 408022 710478
rect 407786 709922 408022 710158
rect 404186 708362 404422 708598
rect 404186 708042 404422 708278
rect 400586 706482 400822 706718
rect 400586 706162 400822 706398
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 425786 711182 426022 711418
rect 425786 710862 426022 711098
rect 422186 709302 422422 709538
rect 422186 708982 422422 709218
rect 418586 707422 418822 707658
rect 418586 707102 418822 707338
rect 414986 705542 415222 705778
rect 414986 705222 415222 705458
rect 443786 710242 444022 710478
rect 443786 709922 444022 710158
rect 440186 708362 440422 708598
rect 440186 708042 440422 708278
rect 436586 706482 436822 706718
rect 436586 706162 436822 706398
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 461786 711182 462022 711418
rect 461786 710862 462022 711098
rect 458186 709302 458422 709538
rect 458186 708982 458422 709218
rect 454586 707422 454822 707658
rect 454586 707102 454822 707338
rect 450986 705542 451222 705778
rect 450986 705222 451222 705458
rect 18926 692462 19162 692698
rect 27022 692462 27258 692698
rect 76886 692462 77122 692698
rect 85166 692462 85402 692698
rect 479786 710242 480022 710478
rect 479786 709922 480022 710158
rect 476186 708362 476422 708598
rect 476186 708042 476422 708278
rect 472586 706482 472822 706718
rect 472586 706162 472822 706398
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 497786 711182 498022 711418
rect 497786 710862 498022 711098
rect 494186 709302 494422 709538
rect 494186 708982 494422 709218
rect 490586 707422 490822 707658
rect 490586 707102 490822 707338
rect 486986 705542 487222 705778
rect 486986 705222 487222 705458
rect 515786 710242 516022 710478
rect 515786 709922 516022 710158
rect 512186 708362 512422 708598
rect 512186 708042 512422 708278
rect 508586 706482 508822 706718
rect 508586 706162 508822 706398
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 533786 711182 534022 711418
rect 533786 710862 534022 711098
rect 530186 709302 530422 709538
rect 530186 708982 530422 709218
rect 526586 707422 526822 707658
rect 526586 707102 526822 707338
rect 522986 705542 523222 705778
rect 522986 705222 523222 705458
rect 551786 710242 552022 710478
rect 551786 709922 552022 710158
rect 548186 708362 548422 708598
rect 548186 708042 548422 708278
rect 544586 706482 544822 706718
rect 544586 706162 544822 706398
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 569786 711182 570022 711418
rect 569786 710862 570022 711098
rect 566186 709302 566422 709538
rect 566186 708982 566422 709218
rect 562586 707422 562822 707658
rect 562586 707102 562822 707338
rect 558986 705542 559222 705778
rect 558986 705222 559222 705458
rect 592082 711182 592318 711418
rect 592082 710862 592318 711098
rect 591142 710242 591378 710478
rect 591142 709922 591378 710158
rect 590202 709302 590438 709538
rect 590202 708982 590438 709218
rect 589262 708362 589498 708598
rect 589262 708042 589498 708278
rect 588322 707422 588558 707658
rect 588322 707102 588558 707338
rect 580586 706482 580822 706718
rect 580586 706162 580822 706398
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 4586 689818 4822 690054
rect 4586 689498 4822 689734
rect 4586 653818 4822 654054
rect 4586 653498 4822 653734
rect 4586 617818 4822 618054
rect 4586 617498 4822 617734
rect 4586 581818 4822 582054
rect 4586 581498 4822 581734
rect 4586 545818 4822 546054
rect 4586 545498 4822 545734
rect 4586 509818 4822 510054
rect 4586 509498 4822 509734
rect 4586 473818 4822 474054
rect 4586 473498 4822 473734
rect 4586 437818 4822 438054
rect 4586 437498 4822 437734
rect 4586 401818 4822 402054
rect 4586 401498 4822 401734
rect 4586 365818 4822 366054
rect 4586 365498 4822 365734
rect 4586 329818 4822 330054
rect 4586 329498 4822 329734
rect 4586 293818 4822 294054
rect 4586 293498 4822 293734
rect 4586 257818 4822 258054
rect 4586 257498 4822 257734
rect 4586 221818 4822 222054
rect 4586 221498 4822 221734
rect 4586 185818 4822 186054
rect 4586 185498 4822 185734
rect 4586 149818 4822 150054
rect 4586 149498 4822 149734
rect 4586 113818 4822 114054
rect 4586 113498 4822 113734
rect 4586 77818 4822 78054
rect 4586 77498 4822 77734
rect 4586 41818 4822 42054
rect 4586 41498 4822 41734
rect 4586 5818 4822 6054
rect 587382 706482 587618 706718
rect 587382 706162 587618 706398
rect 586442 705542 586678 705778
rect 586442 705222 586678 705458
rect 580586 689818 580822 690054
rect 580586 689498 580822 689734
rect 580586 653818 580822 654054
rect 580586 653498 580822 653734
rect 580586 617818 580822 618054
rect 580586 617498 580822 617734
rect 580586 581818 580822 582054
rect 580586 581498 580822 581734
rect 580586 545818 580822 546054
rect 580586 545498 580822 545734
rect 580586 509818 580822 510054
rect 580586 509498 580822 509734
rect 580586 473818 580822 474054
rect 580586 473498 580822 473734
rect 580586 437818 580822 438054
rect 580586 437498 580822 437734
rect 580586 401818 580822 402054
rect 580586 401498 580822 401734
rect 580586 365818 580822 366054
rect 580586 365498 580822 365734
rect 580586 329818 580822 330054
rect 580586 329498 580822 329734
rect 580586 293818 580822 294054
rect 580586 293498 580822 293734
rect 580586 257818 580822 258054
rect 580586 257498 580822 257734
rect 580586 221818 580822 222054
rect 580586 221498 580822 221734
rect 580586 185818 580822 186054
rect 580586 185498 580822 185734
rect 580586 149818 580822 150054
rect 580586 149498 580822 149734
rect 580586 113818 580822 114054
rect 580586 113498 580822 113734
rect 580586 77818 580822 78054
rect 580586 77498 580822 77734
rect 580586 41818 580822 42054
rect 580586 41498 580822 41734
rect 4586 5498 4822 5734
rect -3694 -2462 -3458 -2226
rect -3694 -2782 -3458 -2546
rect 4586 -2462 4822 -2226
rect 4586 -2782 4822 -2546
rect -4634 -3402 -4398 -3166
rect -4634 -3722 -4398 -3486
rect -5574 -4342 -5338 -4106
rect -5574 -4662 -5338 -4426
rect 8186 -4342 8422 -4106
rect 8186 -4662 8422 -4426
rect -6514 -5282 -6278 -5046
rect -6514 -5602 -6278 -5366
rect -7454 -6222 -7218 -5986
rect -7454 -6542 -7218 -6306
rect 18986 -1522 19222 -1286
rect 18986 -1842 19222 -1606
rect 22586 -3402 22822 -3166
rect 22586 -3722 22822 -3486
rect 26186 -5282 26422 -5046
rect 26186 -5602 26422 -5366
rect 11786 -6222 12022 -5986
rect 11786 -6542 12022 -6306
rect -8394 -7162 -8158 -6926
rect -8394 -7482 -8158 -7246
rect 36986 2208 37222 2406
rect 36986 2170 36992 2208
rect 36992 2170 37056 2208
rect 37056 2170 37072 2208
rect 37072 2170 37136 2208
rect 37136 2170 37152 2208
rect 37152 2170 37216 2208
rect 37216 2170 37222 2208
rect 36986 1850 37222 2086
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 40586 -2462 40822 -2226
rect 40586 -2782 40822 -2546
rect 44186 -4342 44422 -4106
rect 44186 -4662 44422 -4426
rect 29786 -7162 30022 -6926
rect 29786 -7482 30022 -7246
rect 54986 -1522 55222 -1286
rect 54986 -1842 55222 -1606
rect 58586 -3402 58822 -3166
rect 58586 -3722 58822 -3486
rect 62186 -5282 62422 -5046
rect 62186 -5602 62422 -5366
rect 47786 -6222 48022 -5986
rect 47786 -6542 48022 -6306
rect 72986 2208 73222 2406
rect 72986 2170 72992 2208
rect 72992 2170 73056 2208
rect 73056 2170 73072 2208
rect 73072 2170 73136 2208
rect 73136 2170 73152 2208
rect 73152 2170 73216 2208
rect 73216 2170 73222 2208
rect 72986 1850 73222 2086
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76586 -2462 76822 -2226
rect 76586 -2782 76822 -2546
rect 80186 -4342 80422 -4106
rect 80186 -4662 80422 -4426
rect 65786 -7162 66022 -6926
rect 65786 -7482 66022 -7246
rect 90986 -1522 91222 -1286
rect 90986 -1842 91222 -1606
rect 94586 -3402 94822 -3166
rect 94586 -3722 94822 -3486
rect 98186 -5282 98422 -5046
rect 98186 -5602 98422 -5366
rect 83786 -6222 84022 -5986
rect 83786 -6542 84022 -6306
rect 108986 2208 109222 2406
rect 108986 2170 108992 2208
rect 108992 2170 109056 2208
rect 109056 2170 109072 2208
rect 109072 2170 109136 2208
rect 109136 2170 109152 2208
rect 109152 2170 109216 2208
rect 109216 2170 109222 2208
rect 108986 1850 109222 2086
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112586 -2462 112822 -2226
rect 112586 -2782 112822 -2546
rect 116186 -4342 116422 -4106
rect 116186 -4662 116422 -4426
rect 101786 -7162 102022 -6926
rect 101786 -7482 102022 -7246
rect 126986 -1522 127222 -1286
rect 126986 -1842 127222 -1606
rect 130586 -3402 130822 -3166
rect 130586 -3722 130822 -3486
rect 134186 -5282 134422 -5046
rect 134186 -5602 134422 -5366
rect 119786 -6222 120022 -5986
rect 119786 -6542 120022 -6306
rect 144986 2208 145222 2406
rect 144986 2170 144992 2208
rect 144992 2170 145056 2208
rect 145056 2170 145072 2208
rect 145072 2170 145136 2208
rect 145136 2170 145152 2208
rect 145152 2170 145216 2208
rect 145216 2170 145222 2208
rect 144986 1850 145222 2086
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148586 -2462 148822 -2226
rect 148586 -2782 148822 -2546
rect 152186 -4342 152422 -4106
rect 152186 -4662 152422 -4426
rect 137786 -7162 138022 -6926
rect 137786 -7482 138022 -7246
rect 162986 -1522 163222 -1286
rect 162986 -1842 163222 -1606
rect 166586 -3402 166822 -3166
rect 166586 -3722 166822 -3486
rect 170186 -5282 170422 -5046
rect 170186 -5602 170422 -5366
rect 155786 -6222 156022 -5986
rect 155786 -6542 156022 -6306
rect 180986 2208 181222 2406
rect 180986 2170 180992 2208
rect 180992 2170 181056 2208
rect 181056 2170 181072 2208
rect 181072 2170 181136 2208
rect 181136 2170 181152 2208
rect 181152 2170 181216 2208
rect 181216 2170 181222 2208
rect 180986 1850 181222 2086
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 -2462 184822 -2226
rect 184586 -2782 184822 -2546
rect 188186 -4342 188422 -4106
rect 188186 -4662 188422 -4426
rect 173786 -7162 174022 -6926
rect 173786 -7482 174022 -7246
rect 198986 -1522 199222 -1286
rect 198986 -1842 199222 -1606
rect 202586 -3402 202822 -3166
rect 202586 -3722 202822 -3486
rect 206186 -5282 206422 -5046
rect 206186 -5602 206422 -5366
rect 191786 -6222 192022 -5986
rect 191786 -6542 192022 -6306
rect 216986 2208 217222 2406
rect 216986 2170 216992 2208
rect 216992 2170 217056 2208
rect 217056 2170 217072 2208
rect 217072 2170 217136 2208
rect 217136 2170 217152 2208
rect 217152 2170 217216 2208
rect 217216 2170 217222 2208
rect 216986 1850 217222 2086
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 -2462 220822 -2226
rect 220586 -2782 220822 -2546
rect 224186 -4342 224422 -4106
rect 224186 -4662 224422 -4426
rect 209786 -7162 210022 -6926
rect 209786 -7482 210022 -7246
rect 234986 -1522 235222 -1286
rect 234986 -1842 235222 -1606
rect 238586 -3402 238822 -3166
rect 238586 -3722 238822 -3486
rect 242186 -5282 242422 -5046
rect 242186 -5602 242422 -5366
rect 227786 -6222 228022 -5986
rect 227786 -6542 228022 -6306
rect 252986 2208 253222 2406
rect 252986 2170 252992 2208
rect 252992 2170 253056 2208
rect 253056 2170 253072 2208
rect 253072 2170 253136 2208
rect 253136 2170 253152 2208
rect 253152 2170 253216 2208
rect 253216 2170 253222 2208
rect 252986 1850 253222 2086
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256586 -2462 256822 -2226
rect 256586 -2782 256822 -2546
rect 260186 -4342 260422 -4106
rect 260186 -4662 260422 -4426
rect 245786 -7162 246022 -6926
rect 245786 -7482 246022 -7246
rect 270986 -1522 271222 -1286
rect 270986 -1842 271222 -1606
rect 274586 -3402 274822 -3166
rect 274586 -3722 274822 -3486
rect 278186 -5282 278422 -5046
rect 278186 -5602 278422 -5366
rect 263786 -6222 264022 -5986
rect 263786 -6542 264022 -6306
rect 288986 2208 289222 2406
rect 288986 2170 288992 2208
rect 288992 2170 289056 2208
rect 289056 2170 289072 2208
rect 289072 2170 289136 2208
rect 289136 2170 289152 2208
rect 289152 2170 289216 2208
rect 289216 2170 289222 2208
rect 288986 1850 289222 2086
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 -2462 292822 -2226
rect 292586 -2782 292822 -2546
rect 296186 -4342 296422 -4106
rect 296186 -4662 296422 -4426
rect 281786 -7162 282022 -6926
rect 281786 -7482 282022 -7246
rect 306986 -1522 307222 -1286
rect 306986 -1842 307222 -1606
rect 310586 -3402 310822 -3166
rect 310586 -3722 310822 -3486
rect 314186 -5282 314422 -5046
rect 314186 -5602 314422 -5366
rect 299786 -6222 300022 -5986
rect 299786 -6542 300022 -6306
rect 324986 2208 325222 2406
rect 324986 2170 324992 2208
rect 324992 2170 325056 2208
rect 325056 2170 325072 2208
rect 325072 2170 325136 2208
rect 325136 2170 325152 2208
rect 325152 2170 325216 2208
rect 325216 2170 325222 2208
rect 324986 1850 325222 2086
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328586 -2462 328822 -2226
rect 328586 -2782 328822 -2546
rect 332186 -4342 332422 -4106
rect 332186 -4662 332422 -4426
rect 317786 -7162 318022 -6926
rect 317786 -7482 318022 -7246
rect 342986 -1522 343222 -1286
rect 342986 -1842 343222 -1606
rect 346586 -3402 346822 -3166
rect 346586 -3722 346822 -3486
rect 350186 -5282 350422 -5046
rect 350186 -5602 350422 -5366
rect 335786 -6222 336022 -5986
rect 335786 -6542 336022 -6306
rect 360986 2208 361222 2406
rect 360986 2170 360992 2208
rect 360992 2170 361056 2208
rect 361056 2170 361072 2208
rect 361072 2170 361136 2208
rect 361136 2170 361152 2208
rect 361152 2170 361216 2208
rect 361216 2170 361222 2208
rect 360986 1850 361222 2086
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 -2462 364822 -2226
rect 364586 -2782 364822 -2546
rect 368186 -4342 368422 -4106
rect 368186 -4662 368422 -4426
rect 353786 -7162 354022 -6926
rect 353786 -7482 354022 -7246
rect 378986 -1522 379222 -1286
rect 378986 -1842 379222 -1606
rect 382586 -3402 382822 -3166
rect 382586 -3722 382822 -3486
rect 386186 -5282 386422 -5046
rect 386186 -5602 386422 -5366
rect 371786 -6222 372022 -5986
rect 371786 -6542 372022 -6306
rect 396986 2208 397222 2406
rect 396986 2170 396992 2208
rect 396992 2170 397056 2208
rect 397056 2170 397072 2208
rect 397072 2170 397136 2208
rect 397136 2170 397152 2208
rect 397152 2170 397216 2208
rect 397216 2170 397222 2208
rect 396986 1850 397222 2086
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400586 -2462 400822 -2226
rect 400586 -2782 400822 -2546
rect 404186 -4342 404422 -4106
rect 404186 -4662 404422 -4426
rect 389786 -7162 390022 -6926
rect 389786 -7482 390022 -7246
rect 414986 -1522 415222 -1286
rect 414986 -1842 415222 -1606
rect 418586 -3402 418822 -3166
rect 418586 -3722 418822 -3486
rect 422186 -5282 422422 -5046
rect 422186 -5602 422422 -5366
rect 407786 -6222 408022 -5986
rect 407786 -6542 408022 -6306
rect 432986 2208 433222 2406
rect 432986 2170 432992 2208
rect 432992 2170 433056 2208
rect 433056 2170 433072 2208
rect 433072 2170 433136 2208
rect 433136 2170 433152 2208
rect 433152 2170 433216 2208
rect 433216 2170 433222 2208
rect 432986 1850 433222 2086
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436586 -2462 436822 -2226
rect 436586 -2782 436822 -2546
rect 440186 -4342 440422 -4106
rect 440186 -4662 440422 -4426
rect 425786 -7162 426022 -6926
rect 425786 -7482 426022 -7246
rect 450986 -1522 451222 -1286
rect 450986 -1842 451222 -1606
rect 454586 -3402 454822 -3166
rect 454586 -3722 454822 -3486
rect 458186 -5282 458422 -5046
rect 458186 -5602 458422 -5366
rect 443786 -6222 444022 -5986
rect 443786 -6542 444022 -6306
rect 468986 2208 469222 2406
rect 468986 2170 468992 2208
rect 468992 2170 469056 2208
rect 469056 2170 469072 2208
rect 469072 2170 469136 2208
rect 469136 2170 469152 2208
rect 469152 2170 469216 2208
rect 469216 2170 469222 2208
rect 468986 1850 469222 2086
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472586 -2462 472822 -2226
rect 472586 -2782 472822 -2546
rect 476186 -4342 476422 -4106
rect 476186 -4662 476422 -4426
rect 461786 -7162 462022 -6926
rect 461786 -7482 462022 -7246
rect 486986 -1522 487222 -1286
rect 486986 -1842 487222 -1606
rect 490586 -3402 490822 -3166
rect 490586 -3722 490822 -3486
rect 494186 -5282 494422 -5046
rect 494186 -5602 494422 -5366
rect 479786 -6222 480022 -5986
rect 479786 -6542 480022 -6306
rect 504986 2208 505222 2406
rect 504986 2170 504992 2208
rect 504992 2170 505056 2208
rect 505056 2170 505072 2208
rect 505072 2170 505136 2208
rect 505136 2170 505152 2208
rect 505152 2170 505216 2208
rect 505216 2170 505222 2208
rect 504986 1850 505222 2086
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508586 -2462 508822 -2226
rect 508586 -2782 508822 -2546
rect 512186 -4342 512422 -4106
rect 512186 -4662 512422 -4426
rect 497786 -7162 498022 -6926
rect 497786 -7482 498022 -7246
rect 522986 -1522 523222 -1286
rect 522986 -1842 523222 -1606
rect 526586 -3402 526822 -3166
rect 526586 -3722 526822 -3486
rect 530186 -5282 530422 -5046
rect 530186 -5602 530422 -5366
rect 515786 -6222 516022 -5986
rect 515786 -6542 516022 -6306
rect 540986 2208 541222 2406
rect 540986 2170 540992 2208
rect 540992 2170 541056 2208
rect 541056 2170 541072 2208
rect 541072 2170 541136 2208
rect 541136 2170 541152 2208
rect 541152 2170 541216 2208
rect 541216 2170 541222 2208
rect 540986 1850 541222 2086
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544586 -2462 544822 -2226
rect 544586 -2782 544822 -2546
rect 548186 -4342 548422 -4106
rect 548186 -4662 548422 -4426
rect 533786 -7162 534022 -6926
rect 533786 -7482 534022 -7246
rect 558986 -1522 559222 -1286
rect 558986 -1842 559222 -1606
rect 562586 -3402 562822 -3166
rect 562586 -3722 562822 -3486
rect 566186 -5282 566422 -5046
rect 566186 -5602 566422 -5366
rect 551786 -6222 552022 -5986
rect 551786 -6542 552022 -6306
rect 576986 2208 577222 2406
rect 576986 2170 576992 2208
rect 576992 2170 577056 2208
rect 577056 2170 577072 2208
rect 577072 2170 577136 2208
rect 577136 2170 577152 2208
rect 577152 2170 577216 2208
rect 577216 2170 577222 2208
rect 576986 1850 577222 2086
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 580586 5818 580822 6054
rect 580586 5498 580822 5734
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686170 585738 686406
rect 585502 685850 585738 686086
rect 585502 650170 585738 650406
rect 585502 649850 585738 650086
rect 585502 614170 585738 614406
rect 585502 613850 585738 614086
rect 585502 578170 585738 578406
rect 585502 577850 585738 578086
rect 585502 542170 585738 542406
rect 585502 541850 585738 542086
rect 585502 506170 585738 506406
rect 585502 505850 585738 506086
rect 585502 470170 585738 470406
rect 585502 469850 585738 470086
rect 585502 434170 585738 434406
rect 585502 433850 585738 434086
rect 585502 398170 585738 398406
rect 585502 397850 585738 398086
rect 585502 362170 585738 362406
rect 585502 361850 585738 362086
rect 585502 326170 585738 326406
rect 585502 325850 585738 326086
rect 585502 290170 585738 290406
rect 585502 289850 585738 290086
rect 585502 254170 585738 254406
rect 585502 253850 585738 254086
rect 585502 218170 585738 218406
rect 585502 217850 585738 218086
rect 585502 182170 585738 182406
rect 585502 181850 585738 182086
rect 585502 146170 585738 146406
rect 585502 145850 585738 146086
rect 585502 110170 585738 110406
rect 585502 109850 585738 110086
rect 585502 74170 585738 74406
rect 585502 73850 585738 74086
rect 585502 38170 585738 38406
rect 585502 37850 585738 38086
rect 585502 2170 585738 2406
rect 585502 1850 585738 2086
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586442 668170 586678 668406
rect 586442 667850 586678 668086
rect 586442 632170 586678 632406
rect 586442 631850 586678 632086
rect 586442 596170 586678 596406
rect 586442 595850 586678 596086
rect 586442 560170 586678 560406
rect 586442 559850 586678 560086
rect 586442 524170 586678 524406
rect 586442 523850 586678 524086
rect 586442 488170 586678 488406
rect 586442 487850 586678 488086
rect 586442 452170 586678 452406
rect 586442 451850 586678 452086
rect 586442 416170 586678 416406
rect 586442 415850 586678 416086
rect 586442 380170 586678 380406
rect 586442 379850 586678 380086
rect 586442 344170 586678 344406
rect 586442 343850 586678 344086
rect 586442 308170 586678 308406
rect 586442 307850 586678 308086
rect 586442 272170 586678 272406
rect 586442 271850 586678 272086
rect 586442 236170 586678 236406
rect 586442 235850 586678 236086
rect 586442 200170 586678 200406
rect 586442 199850 586678 200086
rect 586442 164170 586678 164406
rect 586442 163850 586678 164086
rect 586442 128170 586678 128406
rect 586442 127850 586678 128086
rect 586442 92170 586678 92406
rect 586442 91850 586678 92086
rect 586442 56170 586678 56406
rect 586442 55850 586678 56086
rect 586442 20170 586678 20406
rect 586442 19850 586678 20086
rect 586442 -1522 586678 -1286
rect 586442 -1842 586678 -1606
rect 587382 689818 587618 690054
rect 587382 689498 587618 689734
rect 587382 653818 587618 654054
rect 587382 653498 587618 653734
rect 587382 617818 587618 618054
rect 587382 617498 587618 617734
rect 587382 581818 587618 582054
rect 587382 581498 587618 581734
rect 587382 545818 587618 546054
rect 587382 545498 587618 545734
rect 587382 509818 587618 510054
rect 587382 509498 587618 509734
rect 587382 473818 587618 474054
rect 587382 473498 587618 473734
rect 587382 437818 587618 438054
rect 587382 437498 587618 437734
rect 587382 401818 587618 402054
rect 587382 401498 587618 401734
rect 587382 365818 587618 366054
rect 587382 365498 587618 365734
rect 587382 329818 587618 330054
rect 587382 329498 587618 329734
rect 587382 293818 587618 294054
rect 587382 293498 587618 293734
rect 587382 257818 587618 258054
rect 587382 257498 587618 257734
rect 587382 221818 587618 222054
rect 587382 221498 587618 221734
rect 587382 185818 587618 186054
rect 587382 185498 587618 185734
rect 587382 149818 587618 150054
rect 587382 149498 587618 149734
rect 587382 113818 587618 114054
rect 587382 113498 587618 113734
rect 587382 77818 587618 78054
rect 587382 77498 587618 77734
rect 587382 41818 587618 42054
rect 587382 41498 587618 41734
rect 587382 5818 587618 6054
rect 587382 5498 587618 5734
rect 580586 -2462 580822 -2226
rect 580586 -2782 580822 -2546
rect 587382 -2462 587618 -2226
rect 587382 -2782 587618 -2546
rect 588322 671818 588558 672054
rect 588322 671498 588558 671734
rect 588322 635818 588558 636054
rect 588322 635498 588558 635734
rect 588322 599818 588558 600054
rect 588322 599498 588558 599734
rect 588322 563818 588558 564054
rect 588322 563498 588558 563734
rect 588322 527818 588558 528054
rect 588322 527498 588558 527734
rect 588322 491818 588558 492054
rect 588322 491498 588558 491734
rect 588322 455818 588558 456054
rect 588322 455498 588558 455734
rect 588322 419818 588558 420054
rect 588322 419498 588558 419734
rect 588322 383818 588558 384054
rect 588322 383498 588558 383734
rect 588322 347818 588558 348054
rect 588322 347498 588558 347734
rect 588322 311818 588558 312054
rect 588322 311498 588558 311734
rect 588322 275818 588558 276054
rect 588322 275498 588558 275734
rect 588322 239818 588558 240054
rect 588322 239498 588558 239734
rect 588322 203818 588558 204054
rect 588322 203498 588558 203734
rect 588322 167818 588558 168054
rect 588322 167498 588558 167734
rect 588322 131818 588558 132054
rect 588322 131498 588558 131734
rect 588322 95818 588558 96054
rect 588322 95498 588558 95734
rect 588322 59818 588558 60054
rect 588322 59498 588558 59734
rect 588322 23818 588558 24054
rect 588322 23498 588558 23734
rect 588322 -3402 588558 -3166
rect 588322 -3722 588558 -3486
rect 589262 693418 589498 693654
rect 589262 693098 589498 693334
rect 589262 657418 589498 657654
rect 589262 657098 589498 657334
rect 589262 621418 589498 621654
rect 589262 621098 589498 621334
rect 589262 585418 589498 585654
rect 589262 585098 589498 585334
rect 589262 549418 589498 549654
rect 589262 549098 589498 549334
rect 589262 513418 589498 513654
rect 589262 513098 589498 513334
rect 589262 477418 589498 477654
rect 589262 477098 589498 477334
rect 589262 441418 589498 441654
rect 589262 441098 589498 441334
rect 589262 405418 589498 405654
rect 589262 405098 589498 405334
rect 589262 369418 589498 369654
rect 589262 369098 589498 369334
rect 589262 333418 589498 333654
rect 589262 333098 589498 333334
rect 589262 297418 589498 297654
rect 589262 297098 589498 297334
rect 589262 261418 589498 261654
rect 589262 261098 589498 261334
rect 589262 225418 589498 225654
rect 589262 225098 589498 225334
rect 589262 189418 589498 189654
rect 589262 189098 589498 189334
rect 589262 153418 589498 153654
rect 589262 153098 589498 153334
rect 589262 117418 589498 117654
rect 589262 117098 589498 117334
rect 589262 81418 589498 81654
rect 589262 81098 589498 81334
rect 589262 45418 589498 45654
rect 589262 45098 589498 45334
rect 589262 9418 589498 9654
rect 589262 9098 589498 9334
rect 589262 -4342 589498 -4106
rect 589262 -4662 589498 -4426
rect 590202 675418 590438 675654
rect 590202 675098 590438 675334
rect 590202 639418 590438 639654
rect 590202 639098 590438 639334
rect 590202 603418 590438 603654
rect 590202 603098 590438 603334
rect 590202 567418 590438 567654
rect 590202 567098 590438 567334
rect 590202 531418 590438 531654
rect 590202 531098 590438 531334
rect 590202 495418 590438 495654
rect 590202 495098 590438 495334
rect 590202 459418 590438 459654
rect 590202 459098 590438 459334
rect 590202 423418 590438 423654
rect 590202 423098 590438 423334
rect 590202 387418 590438 387654
rect 590202 387098 590438 387334
rect 590202 351418 590438 351654
rect 590202 351098 590438 351334
rect 590202 315418 590438 315654
rect 590202 315098 590438 315334
rect 590202 279418 590438 279654
rect 590202 279098 590438 279334
rect 590202 243418 590438 243654
rect 590202 243098 590438 243334
rect 590202 207418 590438 207654
rect 590202 207098 590438 207334
rect 590202 171418 590438 171654
rect 590202 171098 590438 171334
rect 590202 135418 590438 135654
rect 590202 135098 590438 135334
rect 590202 99418 590438 99654
rect 590202 99098 590438 99334
rect 590202 63418 590438 63654
rect 590202 63098 590438 63334
rect 590202 27418 590438 27654
rect 590202 27098 590438 27334
rect 590202 -5282 590438 -5046
rect 590202 -5602 590438 -5366
rect 591142 697018 591378 697254
rect 591142 696698 591378 696934
rect 591142 661018 591378 661254
rect 591142 660698 591378 660934
rect 591142 625018 591378 625254
rect 591142 624698 591378 624934
rect 591142 589018 591378 589254
rect 591142 588698 591378 588934
rect 591142 553018 591378 553254
rect 591142 552698 591378 552934
rect 591142 517018 591378 517254
rect 591142 516698 591378 516934
rect 591142 481018 591378 481254
rect 591142 480698 591378 480934
rect 591142 445018 591378 445254
rect 591142 444698 591378 444934
rect 591142 409018 591378 409254
rect 591142 408698 591378 408934
rect 591142 373018 591378 373254
rect 591142 372698 591378 372934
rect 591142 337018 591378 337254
rect 591142 336698 591378 336934
rect 591142 301018 591378 301254
rect 591142 300698 591378 300934
rect 591142 265018 591378 265254
rect 591142 264698 591378 264934
rect 591142 229018 591378 229254
rect 591142 228698 591378 228934
rect 591142 193018 591378 193254
rect 591142 192698 591378 192934
rect 591142 157018 591378 157254
rect 591142 156698 591378 156934
rect 591142 121018 591378 121254
rect 591142 120698 591378 120934
rect 591142 85018 591378 85254
rect 591142 84698 591378 84934
rect 591142 49018 591378 49254
rect 591142 48698 591378 48934
rect 591142 13018 591378 13254
rect 591142 12698 591378 12934
rect 591142 -6222 591378 -5986
rect 591142 -6542 591378 -6306
rect 592082 679018 592318 679254
rect 592082 678698 592318 678934
rect 592082 643018 592318 643254
rect 592082 642698 592318 642934
rect 592082 607018 592318 607254
rect 592082 606698 592318 606934
rect 592082 571018 592318 571254
rect 592082 570698 592318 570934
rect 592082 535018 592318 535254
rect 592082 534698 592318 534934
rect 592082 499018 592318 499254
rect 592082 498698 592318 498934
rect 592082 463018 592318 463254
rect 592082 462698 592318 462934
rect 592082 427018 592318 427254
rect 592082 426698 592318 426934
rect 592082 391018 592318 391254
rect 592082 390698 592318 390934
rect 592082 355018 592318 355254
rect 592082 354698 592318 354934
rect 592082 319018 592318 319254
rect 592082 318698 592318 318934
rect 592082 283018 592318 283254
rect 592082 282698 592318 282934
rect 592082 247018 592318 247254
rect 592082 246698 592318 246934
rect 592082 211018 592318 211254
rect 592082 210698 592318 210934
rect 592082 175018 592318 175254
rect 592082 174698 592318 174934
rect 592082 139018 592318 139254
rect 592082 138698 592318 138934
rect 592082 103018 592318 103254
rect 592082 102698 592318 102934
rect 592082 67018 592318 67254
rect 592082 66698 592318 66934
rect 592082 31018 592318 31254
rect 592082 30698 592318 30934
rect 569786 -7162 570022 -6926
rect 569786 -7482 570022 -7246
rect 592082 -7162 592318 -6926
rect 592082 -7482 592318 -7246
<< metal5 >>
rect -8576 711440 -7976 711442
rect 29604 711440 30204 711442
rect 65604 711440 66204 711442
rect 101604 711440 102204 711442
rect 137604 711440 138204 711442
rect 173604 711440 174204 711442
rect 209604 711440 210204 711442
rect 245604 711440 246204 711442
rect 281604 711440 282204 711442
rect 317604 711440 318204 711442
rect 353604 711440 354204 711442
rect 389604 711440 390204 711442
rect 425604 711440 426204 711442
rect 461604 711440 462204 711442
rect 497604 711440 498204 711442
rect 533604 711440 534204 711442
rect 569604 711440 570204 711442
rect 591900 711440 592500 711442
rect -8576 711418 592500 711440
rect -8576 711182 -8394 711418
rect -8158 711182 29786 711418
rect 30022 711182 65786 711418
rect 66022 711182 101786 711418
rect 102022 711182 137786 711418
rect 138022 711182 173786 711418
rect 174022 711182 209786 711418
rect 210022 711182 245786 711418
rect 246022 711182 281786 711418
rect 282022 711182 317786 711418
rect 318022 711182 353786 711418
rect 354022 711182 389786 711418
rect 390022 711182 425786 711418
rect 426022 711182 461786 711418
rect 462022 711182 497786 711418
rect 498022 711182 533786 711418
rect 534022 711182 569786 711418
rect 570022 711182 592082 711418
rect 592318 711182 592500 711418
rect -8576 711098 592500 711182
rect -8576 710862 -8394 711098
rect -8158 710862 29786 711098
rect 30022 710862 65786 711098
rect 66022 710862 101786 711098
rect 102022 710862 137786 711098
rect 138022 710862 173786 711098
rect 174022 710862 209786 711098
rect 210022 710862 245786 711098
rect 246022 710862 281786 711098
rect 282022 710862 317786 711098
rect 318022 710862 353786 711098
rect 354022 710862 389786 711098
rect 390022 710862 425786 711098
rect 426022 710862 461786 711098
rect 462022 710862 497786 711098
rect 498022 710862 533786 711098
rect 534022 710862 569786 711098
rect 570022 710862 592082 711098
rect 592318 710862 592500 711098
rect -8576 710840 592500 710862
rect -8576 710838 -7976 710840
rect 29604 710838 30204 710840
rect 65604 710838 66204 710840
rect 101604 710838 102204 710840
rect 137604 710838 138204 710840
rect 173604 710838 174204 710840
rect 209604 710838 210204 710840
rect 245604 710838 246204 710840
rect 281604 710838 282204 710840
rect 317604 710838 318204 710840
rect 353604 710838 354204 710840
rect 389604 710838 390204 710840
rect 425604 710838 426204 710840
rect 461604 710838 462204 710840
rect 497604 710838 498204 710840
rect 533604 710838 534204 710840
rect 569604 710838 570204 710840
rect 591900 710838 592500 710840
rect -7636 710500 -7036 710502
rect 11604 710500 12204 710502
rect 47604 710500 48204 710502
rect 83604 710500 84204 710502
rect 119604 710500 120204 710502
rect 155604 710500 156204 710502
rect 191604 710500 192204 710502
rect 227604 710500 228204 710502
rect 263604 710500 264204 710502
rect 299604 710500 300204 710502
rect 335604 710500 336204 710502
rect 371604 710500 372204 710502
rect 407604 710500 408204 710502
rect 443604 710500 444204 710502
rect 479604 710500 480204 710502
rect 515604 710500 516204 710502
rect 551604 710500 552204 710502
rect 590960 710500 591560 710502
rect -7636 710478 591560 710500
rect -7636 710242 -7454 710478
rect -7218 710242 11786 710478
rect 12022 710242 47786 710478
rect 48022 710242 83786 710478
rect 84022 710242 119786 710478
rect 120022 710242 155786 710478
rect 156022 710242 191786 710478
rect 192022 710242 227786 710478
rect 228022 710242 263786 710478
rect 264022 710242 299786 710478
rect 300022 710242 335786 710478
rect 336022 710242 371786 710478
rect 372022 710242 407786 710478
rect 408022 710242 443786 710478
rect 444022 710242 479786 710478
rect 480022 710242 515786 710478
rect 516022 710242 551786 710478
rect 552022 710242 591142 710478
rect 591378 710242 591560 710478
rect -7636 710158 591560 710242
rect -7636 709922 -7454 710158
rect -7218 709922 11786 710158
rect 12022 709922 47786 710158
rect 48022 709922 83786 710158
rect 84022 709922 119786 710158
rect 120022 709922 155786 710158
rect 156022 709922 191786 710158
rect 192022 709922 227786 710158
rect 228022 709922 263786 710158
rect 264022 709922 299786 710158
rect 300022 709922 335786 710158
rect 336022 709922 371786 710158
rect 372022 709922 407786 710158
rect 408022 709922 443786 710158
rect 444022 709922 479786 710158
rect 480022 709922 515786 710158
rect 516022 709922 551786 710158
rect 552022 709922 591142 710158
rect 591378 709922 591560 710158
rect -7636 709900 591560 709922
rect -7636 709898 -7036 709900
rect 11604 709898 12204 709900
rect 47604 709898 48204 709900
rect 83604 709898 84204 709900
rect 119604 709898 120204 709900
rect 155604 709898 156204 709900
rect 191604 709898 192204 709900
rect 227604 709898 228204 709900
rect 263604 709898 264204 709900
rect 299604 709898 300204 709900
rect 335604 709898 336204 709900
rect 371604 709898 372204 709900
rect 407604 709898 408204 709900
rect 443604 709898 444204 709900
rect 479604 709898 480204 709900
rect 515604 709898 516204 709900
rect 551604 709898 552204 709900
rect 590960 709898 591560 709900
rect -6696 709560 -6096 709562
rect 26004 709560 26604 709562
rect 62004 709560 62604 709562
rect 98004 709560 98604 709562
rect 134004 709560 134604 709562
rect 170004 709560 170604 709562
rect 206004 709560 206604 709562
rect 242004 709560 242604 709562
rect 278004 709560 278604 709562
rect 314004 709560 314604 709562
rect 350004 709560 350604 709562
rect 386004 709560 386604 709562
rect 422004 709560 422604 709562
rect 458004 709560 458604 709562
rect 494004 709560 494604 709562
rect 530004 709560 530604 709562
rect 566004 709560 566604 709562
rect 590020 709560 590620 709562
rect -6696 709538 590620 709560
rect -6696 709302 -6514 709538
rect -6278 709302 26186 709538
rect 26422 709302 62186 709538
rect 62422 709302 98186 709538
rect 98422 709302 134186 709538
rect 134422 709302 170186 709538
rect 170422 709302 206186 709538
rect 206422 709302 242186 709538
rect 242422 709302 278186 709538
rect 278422 709302 314186 709538
rect 314422 709302 350186 709538
rect 350422 709302 386186 709538
rect 386422 709302 422186 709538
rect 422422 709302 458186 709538
rect 458422 709302 494186 709538
rect 494422 709302 530186 709538
rect 530422 709302 566186 709538
rect 566422 709302 590202 709538
rect 590438 709302 590620 709538
rect -6696 709218 590620 709302
rect -6696 708982 -6514 709218
rect -6278 708982 26186 709218
rect 26422 708982 62186 709218
rect 62422 708982 98186 709218
rect 98422 708982 134186 709218
rect 134422 708982 170186 709218
rect 170422 708982 206186 709218
rect 206422 708982 242186 709218
rect 242422 708982 278186 709218
rect 278422 708982 314186 709218
rect 314422 708982 350186 709218
rect 350422 708982 386186 709218
rect 386422 708982 422186 709218
rect 422422 708982 458186 709218
rect 458422 708982 494186 709218
rect 494422 708982 530186 709218
rect 530422 708982 566186 709218
rect 566422 708982 590202 709218
rect 590438 708982 590620 709218
rect -6696 708960 590620 708982
rect -6696 708958 -6096 708960
rect 26004 708958 26604 708960
rect 62004 708958 62604 708960
rect 98004 708958 98604 708960
rect 134004 708958 134604 708960
rect 170004 708958 170604 708960
rect 206004 708958 206604 708960
rect 242004 708958 242604 708960
rect 278004 708958 278604 708960
rect 314004 708958 314604 708960
rect 350004 708958 350604 708960
rect 386004 708958 386604 708960
rect 422004 708958 422604 708960
rect 458004 708958 458604 708960
rect 494004 708958 494604 708960
rect 530004 708958 530604 708960
rect 566004 708958 566604 708960
rect 590020 708958 590620 708960
rect -5756 708620 -5156 708622
rect 8004 708620 8604 708622
rect 44004 708620 44604 708622
rect 80004 708620 80604 708622
rect 116004 708620 116604 708622
rect 152004 708620 152604 708622
rect 188004 708620 188604 708622
rect 224004 708620 224604 708622
rect 260004 708620 260604 708622
rect 296004 708620 296604 708622
rect 332004 708620 332604 708622
rect 368004 708620 368604 708622
rect 404004 708620 404604 708622
rect 440004 708620 440604 708622
rect 476004 708620 476604 708622
rect 512004 708620 512604 708622
rect 548004 708620 548604 708622
rect 589080 708620 589680 708622
rect -5756 708598 589680 708620
rect -5756 708362 -5574 708598
rect -5338 708362 8186 708598
rect 8422 708362 44186 708598
rect 44422 708362 80186 708598
rect 80422 708362 116186 708598
rect 116422 708362 152186 708598
rect 152422 708362 188186 708598
rect 188422 708362 224186 708598
rect 224422 708362 260186 708598
rect 260422 708362 296186 708598
rect 296422 708362 332186 708598
rect 332422 708362 368186 708598
rect 368422 708362 404186 708598
rect 404422 708362 440186 708598
rect 440422 708362 476186 708598
rect 476422 708362 512186 708598
rect 512422 708362 548186 708598
rect 548422 708362 589262 708598
rect 589498 708362 589680 708598
rect -5756 708278 589680 708362
rect -5756 708042 -5574 708278
rect -5338 708042 8186 708278
rect 8422 708042 44186 708278
rect 44422 708042 80186 708278
rect 80422 708042 116186 708278
rect 116422 708042 152186 708278
rect 152422 708042 188186 708278
rect 188422 708042 224186 708278
rect 224422 708042 260186 708278
rect 260422 708042 296186 708278
rect 296422 708042 332186 708278
rect 332422 708042 368186 708278
rect 368422 708042 404186 708278
rect 404422 708042 440186 708278
rect 440422 708042 476186 708278
rect 476422 708042 512186 708278
rect 512422 708042 548186 708278
rect 548422 708042 589262 708278
rect 589498 708042 589680 708278
rect -5756 708020 589680 708042
rect -5756 708018 -5156 708020
rect 8004 708018 8604 708020
rect 44004 708018 44604 708020
rect 80004 708018 80604 708020
rect 116004 708018 116604 708020
rect 152004 708018 152604 708020
rect 188004 708018 188604 708020
rect 224004 708018 224604 708020
rect 260004 708018 260604 708020
rect 296004 708018 296604 708020
rect 332004 708018 332604 708020
rect 368004 708018 368604 708020
rect 404004 708018 404604 708020
rect 440004 708018 440604 708020
rect 476004 708018 476604 708020
rect 512004 708018 512604 708020
rect 548004 708018 548604 708020
rect 589080 708018 589680 708020
rect -4816 707680 -4216 707682
rect 22404 707680 23004 707682
rect 58404 707680 59004 707682
rect 94404 707680 95004 707682
rect 130404 707680 131004 707682
rect 166404 707680 167004 707682
rect 202404 707680 203004 707682
rect 238404 707680 239004 707682
rect 274404 707680 275004 707682
rect 310404 707680 311004 707682
rect 346404 707680 347004 707682
rect 382404 707680 383004 707682
rect 418404 707680 419004 707682
rect 454404 707680 455004 707682
rect 490404 707680 491004 707682
rect 526404 707680 527004 707682
rect 562404 707680 563004 707682
rect 588140 707680 588740 707682
rect -4816 707658 588740 707680
rect -4816 707422 -4634 707658
rect -4398 707422 22586 707658
rect 22822 707422 58586 707658
rect 58822 707422 94586 707658
rect 94822 707422 130586 707658
rect 130822 707422 166586 707658
rect 166822 707422 202586 707658
rect 202822 707422 238586 707658
rect 238822 707422 274586 707658
rect 274822 707422 310586 707658
rect 310822 707422 346586 707658
rect 346822 707422 382586 707658
rect 382822 707422 418586 707658
rect 418822 707422 454586 707658
rect 454822 707422 490586 707658
rect 490822 707422 526586 707658
rect 526822 707422 562586 707658
rect 562822 707422 588322 707658
rect 588558 707422 588740 707658
rect -4816 707338 588740 707422
rect -4816 707102 -4634 707338
rect -4398 707102 22586 707338
rect 22822 707102 58586 707338
rect 58822 707102 94586 707338
rect 94822 707102 130586 707338
rect 130822 707102 166586 707338
rect 166822 707102 202586 707338
rect 202822 707102 238586 707338
rect 238822 707102 274586 707338
rect 274822 707102 310586 707338
rect 310822 707102 346586 707338
rect 346822 707102 382586 707338
rect 382822 707102 418586 707338
rect 418822 707102 454586 707338
rect 454822 707102 490586 707338
rect 490822 707102 526586 707338
rect 526822 707102 562586 707338
rect 562822 707102 588322 707338
rect 588558 707102 588740 707338
rect -4816 707080 588740 707102
rect -4816 707078 -4216 707080
rect 22404 707078 23004 707080
rect 58404 707078 59004 707080
rect 94404 707078 95004 707080
rect 130404 707078 131004 707080
rect 166404 707078 167004 707080
rect 202404 707078 203004 707080
rect 238404 707078 239004 707080
rect 274404 707078 275004 707080
rect 310404 707078 311004 707080
rect 346404 707078 347004 707080
rect 382404 707078 383004 707080
rect 418404 707078 419004 707080
rect 454404 707078 455004 707080
rect 490404 707078 491004 707080
rect 526404 707078 527004 707080
rect 562404 707078 563004 707080
rect 588140 707078 588740 707080
rect -3876 706740 -3276 706742
rect 4404 706740 5004 706742
rect 40404 706740 41004 706742
rect 76404 706740 77004 706742
rect 112404 706740 113004 706742
rect 148404 706740 149004 706742
rect 184404 706740 185004 706742
rect 220404 706740 221004 706742
rect 256404 706740 257004 706742
rect 292404 706740 293004 706742
rect 328404 706740 329004 706742
rect 364404 706740 365004 706742
rect 400404 706740 401004 706742
rect 436404 706740 437004 706742
rect 472404 706740 473004 706742
rect 508404 706740 509004 706742
rect 544404 706740 545004 706742
rect 580404 706740 581004 706742
rect 587200 706740 587800 706742
rect -3876 706718 587800 706740
rect -3876 706482 -3694 706718
rect -3458 706482 4586 706718
rect 4822 706482 40586 706718
rect 40822 706482 76586 706718
rect 76822 706482 112586 706718
rect 112822 706482 148586 706718
rect 148822 706482 184586 706718
rect 184822 706482 220586 706718
rect 220822 706482 256586 706718
rect 256822 706482 292586 706718
rect 292822 706482 328586 706718
rect 328822 706482 364586 706718
rect 364822 706482 400586 706718
rect 400822 706482 436586 706718
rect 436822 706482 472586 706718
rect 472822 706482 508586 706718
rect 508822 706482 544586 706718
rect 544822 706482 580586 706718
rect 580822 706482 587382 706718
rect 587618 706482 587800 706718
rect -3876 706398 587800 706482
rect -3876 706162 -3694 706398
rect -3458 706162 4586 706398
rect 4822 706162 40586 706398
rect 40822 706162 76586 706398
rect 76822 706162 112586 706398
rect 112822 706162 148586 706398
rect 148822 706162 184586 706398
rect 184822 706162 220586 706398
rect 220822 706162 256586 706398
rect 256822 706162 292586 706398
rect 292822 706162 328586 706398
rect 328822 706162 364586 706398
rect 364822 706162 400586 706398
rect 400822 706162 436586 706398
rect 436822 706162 472586 706398
rect 472822 706162 508586 706398
rect 508822 706162 544586 706398
rect 544822 706162 580586 706398
rect 580822 706162 587382 706398
rect 587618 706162 587800 706398
rect -3876 706140 587800 706162
rect -3876 706138 -3276 706140
rect 4404 706138 5004 706140
rect 40404 706138 41004 706140
rect 76404 706138 77004 706140
rect 112404 706138 113004 706140
rect 148404 706138 149004 706140
rect 184404 706138 185004 706140
rect 220404 706138 221004 706140
rect 256404 706138 257004 706140
rect 292404 706138 293004 706140
rect 328404 706138 329004 706140
rect 364404 706138 365004 706140
rect 400404 706138 401004 706140
rect 436404 706138 437004 706140
rect 472404 706138 473004 706140
rect 508404 706138 509004 706140
rect 544404 706138 545004 706140
rect 580404 706138 581004 706140
rect 587200 706138 587800 706140
rect -2936 705800 -2336 705802
rect 18804 705800 19404 705802
rect 54804 705800 55404 705802
rect 90804 705800 91404 705802
rect 126804 705800 127404 705802
rect 162804 705800 163404 705802
rect 198804 705800 199404 705802
rect 234804 705800 235404 705802
rect 270804 705800 271404 705802
rect 306804 705800 307404 705802
rect 342804 705800 343404 705802
rect 378804 705800 379404 705802
rect 414804 705800 415404 705802
rect 450804 705800 451404 705802
rect 486804 705800 487404 705802
rect 522804 705800 523404 705802
rect 558804 705800 559404 705802
rect 586260 705800 586860 705802
rect -2936 705778 586860 705800
rect -2936 705542 -2754 705778
rect -2518 705542 18986 705778
rect 19222 705542 54986 705778
rect 55222 705542 90986 705778
rect 91222 705542 126986 705778
rect 127222 705542 162986 705778
rect 163222 705542 198986 705778
rect 199222 705542 234986 705778
rect 235222 705542 270986 705778
rect 271222 705542 306986 705778
rect 307222 705542 342986 705778
rect 343222 705542 378986 705778
rect 379222 705542 414986 705778
rect 415222 705542 450986 705778
rect 451222 705542 486986 705778
rect 487222 705542 522986 705778
rect 523222 705542 558986 705778
rect 559222 705542 586442 705778
rect 586678 705542 586860 705778
rect -2936 705458 586860 705542
rect -2936 705222 -2754 705458
rect -2518 705222 18986 705458
rect 19222 705222 54986 705458
rect 55222 705222 90986 705458
rect 91222 705222 126986 705458
rect 127222 705222 162986 705458
rect 163222 705222 198986 705458
rect 199222 705222 234986 705458
rect 235222 705222 270986 705458
rect 271222 705222 306986 705458
rect 307222 705222 342986 705458
rect 343222 705222 378986 705458
rect 379222 705222 414986 705458
rect 415222 705222 450986 705458
rect 451222 705222 486986 705458
rect 487222 705222 522986 705458
rect 523222 705222 558986 705458
rect 559222 705222 586442 705458
rect 586678 705222 586860 705458
rect -2936 705200 586860 705222
rect -2936 705198 -2336 705200
rect 18804 705198 19404 705200
rect 54804 705198 55404 705200
rect 90804 705198 91404 705200
rect 126804 705198 127404 705200
rect 162804 705198 163404 705200
rect 198804 705198 199404 705200
rect 234804 705198 235404 705200
rect 270804 705198 271404 705200
rect 306804 705198 307404 705200
rect 342804 705198 343404 705200
rect 378804 705198 379404 705200
rect 414804 705198 415404 705200
rect 450804 705198 451404 705200
rect 486804 705198 487404 705200
rect 522804 705198 523404 705200
rect 558804 705198 559404 705200
rect 586260 705198 586860 705200
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -7636 697276 -7036 697278
rect 590960 697276 591560 697278
rect -8576 697254 592500 697276
rect -8576 697018 -7454 697254
rect -7218 697018 591142 697254
rect 591378 697018 592500 697254
rect -8576 696934 592500 697018
rect -8576 696698 -7454 696934
rect -7218 696698 591142 696934
rect 591378 696698 592500 696934
rect -8576 696676 592500 696698
rect -7636 696674 -7036 696676
rect 590960 696674 591560 696676
rect -5756 693676 -5156 693678
rect 589080 693676 589680 693678
rect -6696 693654 590620 693676
rect -6696 693418 -5574 693654
rect -5338 693418 589262 693654
rect 589498 693418 590620 693654
rect -6696 693334 590620 693418
rect -6696 693098 -5574 693334
rect -5338 693098 589262 693334
rect 589498 693098 590620 693334
rect -6696 693076 590620 693098
rect -5756 693074 -5156 693076
rect 589080 693074 589680 693076
rect 18884 692698 27300 692740
rect 18884 692462 18926 692698
rect 19162 692462 27022 692698
rect 27258 692462 27300 692698
rect 18884 692420 27300 692462
rect 76844 692698 85444 692740
rect 76844 692462 76886 692698
rect 77122 692462 85166 692698
rect 85402 692462 85444 692698
rect 76844 692420 85444 692462
rect -3876 690076 -3276 690078
rect 4404 690076 5004 690078
rect 580404 690076 581004 690078
rect 587200 690076 587800 690078
rect -4816 690054 588740 690076
rect -4816 689818 -3694 690054
rect -3458 689818 4586 690054
rect 4822 689818 580586 690054
rect 580822 689818 587382 690054
rect 587618 689818 588740 690054
rect -4816 689734 588740 689818
rect -4816 689498 -3694 689734
rect -3458 689498 4586 689734
rect 4822 689498 580586 689734
rect 580822 689498 587382 689734
rect 587618 689498 588740 689734
rect -4816 689476 588740 689498
rect -3876 689474 -3276 689476
rect 4404 689474 5004 689476
rect 580404 689474 581004 689476
rect 587200 689474 587800 689476
rect -1996 686428 -1396 686430
rect 804 686428 1404 686430
rect 585320 686428 585920 686430
rect -2936 686406 586860 686428
rect -2936 686170 -1814 686406
rect -1578 686170 986 686406
rect 1222 686170 585502 686406
rect 585738 686170 586860 686406
rect -2936 686086 586860 686170
rect -2936 685850 -1814 686086
rect -1578 685850 986 686086
rect 1222 685850 585502 686086
rect 585738 685850 586860 686086
rect -2936 685828 586860 685850
rect -1996 685826 -1396 685828
rect 804 685826 1404 685828
rect 585320 685826 585920 685828
rect -8576 679276 -7976 679278
rect 591900 679276 592500 679278
rect -8576 679254 592500 679276
rect -8576 679018 -8394 679254
rect -8158 679018 592082 679254
rect 592318 679018 592500 679254
rect -8576 678934 592500 679018
rect -8576 678698 -8394 678934
rect -8158 678698 592082 678934
rect 592318 678698 592500 678934
rect -8576 678676 592500 678698
rect -8576 678674 -7976 678676
rect 591900 678674 592500 678676
rect -6696 675676 -6096 675678
rect 590020 675676 590620 675678
rect -6696 675654 590620 675676
rect -6696 675418 -6514 675654
rect -6278 675418 590202 675654
rect 590438 675418 590620 675654
rect -6696 675334 590620 675418
rect -6696 675098 -6514 675334
rect -6278 675098 590202 675334
rect 590438 675098 590620 675334
rect -6696 675076 590620 675098
rect -6696 675074 -6096 675076
rect 590020 675074 590620 675076
rect -4816 672076 -4216 672078
rect 588140 672076 588740 672078
rect -4816 672054 588740 672076
rect -4816 671818 -4634 672054
rect -4398 671818 588322 672054
rect 588558 671818 588740 672054
rect -4816 671734 588740 671818
rect -4816 671498 -4634 671734
rect -4398 671498 588322 671734
rect 588558 671498 588740 671734
rect -4816 671476 588740 671498
rect -4816 671474 -4216 671476
rect 588140 671474 588740 671476
rect -2936 668428 -2336 668430
rect 586260 668428 586860 668430
rect -2936 668406 586860 668428
rect -2936 668170 -2754 668406
rect -2518 668170 586442 668406
rect 586678 668170 586860 668406
rect -2936 668086 586860 668170
rect -2936 667850 -2754 668086
rect -2518 667850 586442 668086
rect 586678 667850 586860 668086
rect -2936 667828 586860 667850
rect -2936 667826 -2336 667828
rect 586260 667826 586860 667828
rect -7636 661276 -7036 661278
rect 590960 661276 591560 661278
rect -8576 661254 592500 661276
rect -8576 661018 -7454 661254
rect -7218 661018 591142 661254
rect 591378 661018 592500 661254
rect -8576 660934 592500 661018
rect -8576 660698 -7454 660934
rect -7218 660698 591142 660934
rect 591378 660698 592500 660934
rect -8576 660676 592500 660698
rect -7636 660674 -7036 660676
rect 590960 660674 591560 660676
rect -5756 657676 -5156 657678
rect 589080 657676 589680 657678
rect -6696 657654 590620 657676
rect -6696 657418 -5574 657654
rect -5338 657418 589262 657654
rect 589498 657418 590620 657654
rect -6696 657334 590620 657418
rect -6696 657098 -5574 657334
rect -5338 657098 589262 657334
rect 589498 657098 590620 657334
rect -6696 657076 590620 657098
rect -5756 657074 -5156 657076
rect 589080 657074 589680 657076
rect -3876 654076 -3276 654078
rect 4404 654076 5004 654078
rect 580404 654076 581004 654078
rect 587200 654076 587800 654078
rect -4816 654054 588740 654076
rect -4816 653818 -3694 654054
rect -3458 653818 4586 654054
rect 4822 653818 580586 654054
rect 580822 653818 587382 654054
rect 587618 653818 588740 654054
rect -4816 653734 588740 653818
rect -4816 653498 -3694 653734
rect -3458 653498 4586 653734
rect 4822 653498 580586 653734
rect 580822 653498 587382 653734
rect 587618 653498 588740 653734
rect -4816 653476 588740 653498
rect -3876 653474 -3276 653476
rect 4404 653474 5004 653476
rect 580404 653474 581004 653476
rect 587200 653474 587800 653476
rect -1996 650428 -1396 650430
rect 804 650428 1404 650430
rect 585320 650428 585920 650430
rect -2936 650406 586860 650428
rect -2936 650170 -1814 650406
rect -1578 650170 986 650406
rect 1222 650170 585502 650406
rect 585738 650170 586860 650406
rect -2936 650086 586860 650170
rect -2936 649850 -1814 650086
rect -1578 649850 986 650086
rect 1222 649850 585502 650086
rect 585738 649850 586860 650086
rect -2936 649828 586860 649850
rect -1996 649826 -1396 649828
rect 804 649826 1404 649828
rect 585320 649826 585920 649828
rect -8576 643276 -7976 643278
rect 591900 643276 592500 643278
rect -8576 643254 592500 643276
rect -8576 643018 -8394 643254
rect -8158 643018 592082 643254
rect 592318 643018 592500 643254
rect -8576 642934 592500 643018
rect -8576 642698 -8394 642934
rect -8158 642698 592082 642934
rect 592318 642698 592500 642934
rect -8576 642676 592500 642698
rect -8576 642674 -7976 642676
rect 591900 642674 592500 642676
rect -6696 639676 -6096 639678
rect 590020 639676 590620 639678
rect -6696 639654 590620 639676
rect -6696 639418 -6514 639654
rect -6278 639418 590202 639654
rect 590438 639418 590620 639654
rect -6696 639334 590620 639418
rect -6696 639098 -6514 639334
rect -6278 639098 590202 639334
rect 590438 639098 590620 639334
rect -6696 639076 590620 639098
rect -6696 639074 -6096 639076
rect 590020 639074 590620 639076
rect -4816 636076 -4216 636078
rect 588140 636076 588740 636078
rect -4816 636054 588740 636076
rect -4816 635818 -4634 636054
rect -4398 635818 588322 636054
rect 588558 635818 588740 636054
rect -4816 635734 588740 635818
rect -4816 635498 -4634 635734
rect -4398 635498 588322 635734
rect 588558 635498 588740 635734
rect -4816 635476 588740 635498
rect -4816 635474 -4216 635476
rect 588140 635474 588740 635476
rect -2936 632428 -2336 632430
rect 586260 632428 586860 632430
rect -2936 632406 586860 632428
rect -2936 632170 -2754 632406
rect -2518 632170 586442 632406
rect 586678 632170 586860 632406
rect -2936 632086 586860 632170
rect -2936 631850 -2754 632086
rect -2518 631850 586442 632086
rect 586678 631850 586860 632086
rect -2936 631828 586860 631850
rect -2936 631826 -2336 631828
rect 586260 631826 586860 631828
rect -7636 625276 -7036 625278
rect 590960 625276 591560 625278
rect -8576 625254 592500 625276
rect -8576 625018 -7454 625254
rect -7218 625018 591142 625254
rect 591378 625018 592500 625254
rect -8576 624934 592500 625018
rect -8576 624698 -7454 624934
rect -7218 624698 591142 624934
rect 591378 624698 592500 624934
rect -8576 624676 592500 624698
rect -7636 624674 -7036 624676
rect 590960 624674 591560 624676
rect -5756 621676 -5156 621678
rect 589080 621676 589680 621678
rect -6696 621654 590620 621676
rect -6696 621418 -5574 621654
rect -5338 621418 589262 621654
rect 589498 621418 590620 621654
rect -6696 621334 590620 621418
rect -6696 621098 -5574 621334
rect -5338 621098 589262 621334
rect 589498 621098 590620 621334
rect -6696 621076 590620 621098
rect -5756 621074 -5156 621076
rect 589080 621074 589680 621076
rect -3876 618076 -3276 618078
rect 4404 618076 5004 618078
rect 580404 618076 581004 618078
rect 587200 618076 587800 618078
rect -4816 618054 588740 618076
rect -4816 617818 -3694 618054
rect -3458 617818 4586 618054
rect 4822 617818 580586 618054
rect 580822 617818 587382 618054
rect 587618 617818 588740 618054
rect -4816 617734 588740 617818
rect -4816 617498 -3694 617734
rect -3458 617498 4586 617734
rect 4822 617498 580586 617734
rect 580822 617498 587382 617734
rect 587618 617498 588740 617734
rect -4816 617476 588740 617498
rect -3876 617474 -3276 617476
rect 4404 617474 5004 617476
rect 580404 617474 581004 617476
rect 587200 617474 587800 617476
rect -1996 614428 -1396 614430
rect 804 614428 1404 614430
rect 585320 614428 585920 614430
rect -2936 614406 586860 614428
rect -2936 614170 -1814 614406
rect -1578 614170 986 614406
rect 1222 614170 585502 614406
rect 585738 614170 586860 614406
rect -2936 614086 586860 614170
rect -2936 613850 -1814 614086
rect -1578 613850 986 614086
rect 1222 613850 585502 614086
rect 585738 613850 586860 614086
rect -2936 613828 586860 613850
rect -1996 613826 -1396 613828
rect 804 613826 1404 613828
rect 585320 613826 585920 613828
rect -8576 607276 -7976 607278
rect 591900 607276 592500 607278
rect -8576 607254 592500 607276
rect -8576 607018 -8394 607254
rect -8158 607018 592082 607254
rect 592318 607018 592500 607254
rect -8576 606934 592500 607018
rect -8576 606698 -8394 606934
rect -8158 606698 592082 606934
rect 592318 606698 592500 606934
rect -8576 606676 592500 606698
rect -8576 606674 -7976 606676
rect 591900 606674 592500 606676
rect -6696 603676 -6096 603678
rect 590020 603676 590620 603678
rect -6696 603654 590620 603676
rect -6696 603418 -6514 603654
rect -6278 603418 590202 603654
rect 590438 603418 590620 603654
rect -6696 603334 590620 603418
rect -6696 603098 -6514 603334
rect -6278 603098 590202 603334
rect 590438 603098 590620 603334
rect -6696 603076 590620 603098
rect -6696 603074 -6096 603076
rect 590020 603074 590620 603076
rect -4816 600076 -4216 600078
rect 588140 600076 588740 600078
rect -4816 600054 588740 600076
rect -4816 599818 -4634 600054
rect -4398 599818 588322 600054
rect 588558 599818 588740 600054
rect -4816 599734 588740 599818
rect -4816 599498 -4634 599734
rect -4398 599498 588322 599734
rect 588558 599498 588740 599734
rect -4816 599476 588740 599498
rect -4816 599474 -4216 599476
rect 588140 599474 588740 599476
rect -2936 596428 -2336 596430
rect 586260 596428 586860 596430
rect -2936 596406 586860 596428
rect -2936 596170 -2754 596406
rect -2518 596170 586442 596406
rect 586678 596170 586860 596406
rect -2936 596086 586860 596170
rect -2936 595850 -2754 596086
rect -2518 595850 586442 596086
rect 586678 595850 586860 596086
rect -2936 595828 586860 595850
rect -2936 595826 -2336 595828
rect 586260 595826 586860 595828
rect -7636 589276 -7036 589278
rect 590960 589276 591560 589278
rect -8576 589254 592500 589276
rect -8576 589018 -7454 589254
rect -7218 589018 591142 589254
rect 591378 589018 592500 589254
rect -8576 588934 592500 589018
rect -8576 588698 -7454 588934
rect -7218 588698 591142 588934
rect 591378 588698 592500 588934
rect -8576 588676 592500 588698
rect -7636 588674 -7036 588676
rect 590960 588674 591560 588676
rect -5756 585676 -5156 585678
rect 589080 585676 589680 585678
rect -6696 585654 590620 585676
rect -6696 585418 -5574 585654
rect -5338 585418 589262 585654
rect 589498 585418 590620 585654
rect -6696 585334 590620 585418
rect -6696 585098 -5574 585334
rect -5338 585098 589262 585334
rect 589498 585098 590620 585334
rect -6696 585076 590620 585098
rect -5756 585074 -5156 585076
rect 589080 585074 589680 585076
rect -3876 582076 -3276 582078
rect 4404 582076 5004 582078
rect 580404 582076 581004 582078
rect 587200 582076 587800 582078
rect -4816 582054 588740 582076
rect -4816 581818 -3694 582054
rect -3458 581818 4586 582054
rect 4822 581818 580586 582054
rect 580822 581818 587382 582054
rect 587618 581818 588740 582054
rect -4816 581734 588740 581818
rect -4816 581498 -3694 581734
rect -3458 581498 4586 581734
rect 4822 581498 580586 581734
rect 580822 581498 587382 581734
rect 587618 581498 588740 581734
rect -4816 581476 588740 581498
rect -3876 581474 -3276 581476
rect 4404 581474 5004 581476
rect 580404 581474 581004 581476
rect 587200 581474 587800 581476
rect -1996 578428 -1396 578430
rect 804 578428 1404 578430
rect 585320 578428 585920 578430
rect -2936 578406 586860 578428
rect -2936 578170 -1814 578406
rect -1578 578170 986 578406
rect 1222 578170 585502 578406
rect 585738 578170 586860 578406
rect -2936 578086 586860 578170
rect -2936 577850 -1814 578086
rect -1578 577850 986 578086
rect 1222 577850 585502 578086
rect 585738 577850 586860 578086
rect -2936 577828 586860 577850
rect -1996 577826 -1396 577828
rect 804 577826 1404 577828
rect 585320 577826 585920 577828
rect -8576 571276 -7976 571278
rect 591900 571276 592500 571278
rect -8576 571254 592500 571276
rect -8576 571018 -8394 571254
rect -8158 571018 592082 571254
rect 592318 571018 592500 571254
rect -8576 570934 592500 571018
rect -8576 570698 -8394 570934
rect -8158 570698 592082 570934
rect 592318 570698 592500 570934
rect -8576 570676 592500 570698
rect -8576 570674 -7976 570676
rect 591900 570674 592500 570676
rect -6696 567676 -6096 567678
rect 590020 567676 590620 567678
rect -6696 567654 590620 567676
rect -6696 567418 -6514 567654
rect -6278 567418 590202 567654
rect 590438 567418 590620 567654
rect -6696 567334 590620 567418
rect -6696 567098 -6514 567334
rect -6278 567098 590202 567334
rect 590438 567098 590620 567334
rect -6696 567076 590620 567098
rect -6696 567074 -6096 567076
rect 590020 567074 590620 567076
rect -4816 564076 -4216 564078
rect 588140 564076 588740 564078
rect -4816 564054 588740 564076
rect -4816 563818 -4634 564054
rect -4398 563818 588322 564054
rect 588558 563818 588740 564054
rect -4816 563734 588740 563818
rect -4816 563498 -4634 563734
rect -4398 563498 588322 563734
rect 588558 563498 588740 563734
rect -4816 563476 588740 563498
rect -4816 563474 -4216 563476
rect 588140 563474 588740 563476
rect -2936 560428 -2336 560430
rect 586260 560428 586860 560430
rect -2936 560406 586860 560428
rect -2936 560170 -2754 560406
rect -2518 560170 586442 560406
rect 586678 560170 586860 560406
rect -2936 560086 586860 560170
rect -2936 559850 -2754 560086
rect -2518 559850 586442 560086
rect 586678 559850 586860 560086
rect -2936 559828 586860 559850
rect -2936 559826 -2336 559828
rect 586260 559826 586860 559828
rect -7636 553276 -7036 553278
rect 590960 553276 591560 553278
rect -8576 553254 592500 553276
rect -8576 553018 -7454 553254
rect -7218 553018 591142 553254
rect 591378 553018 592500 553254
rect -8576 552934 592500 553018
rect -8576 552698 -7454 552934
rect -7218 552698 591142 552934
rect 591378 552698 592500 552934
rect -8576 552676 592500 552698
rect -7636 552674 -7036 552676
rect 590960 552674 591560 552676
rect -5756 549676 -5156 549678
rect 589080 549676 589680 549678
rect -6696 549654 590620 549676
rect -6696 549418 -5574 549654
rect -5338 549418 589262 549654
rect 589498 549418 590620 549654
rect -6696 549334 590620 549418
rect -6696 549098 -5574 549334
rect -5338 549098 589262 549334
rect 589498 549098 590620 549334
rect -6696 549076 590620 549098
rect -5756 549074 -5156 549076
rect 589080 549074 589680 549076
rect -3876 546076 -3276 546078
rect 4404 546076 5004 546078
rect 580404 546076 581004 546078
rect 587200 546076 587800 546078
rect -4816 546054 588740 546076
rect -4816 545818 -3694 546054
rect -3458 545818 4586 546054
rect 4822 545818 580586 546054
rect 580822 545818 587382 546054
rect 587618 545818 588740 546054
rect -4816 545734 588740 545818
rect -4816 545498 -3694 545734
rect -3458 545498 4586 545734
rect 4822 545498 580586 545734
rect 580822 545498 587382 545734
rect 587618 545498 588740 545734
rect -4816 545476 588740 545498
rect -3876 545474 -3276 545476
rect 4404 545474 5004 545476
rect 580404 545474 581004 545476
rect 587200 545474 587800 545476
rect -1996 542428 -1396 542430
rect 804 542428 1404 542430
rect 585320 542428 585920 542430
rect -2936 542406 586860 542428
rect -2936 542170 -1814 542406
rect -1578 542170 986 542406
rect 1222 542170 585502 542406
rect 585738 542170 586860 542406
rect -2936 542086 586860 542170
rect -2936 541850 -1814 542086
rect -1578 541850 986 542086
rect 1222 541850 585502 542086
rect 585738 541850 586860 542086
rect -2936 541828 586860 541850
rect -1996 541826 -1396 541828
rect 804 541826 1404 541828
rect 585320 541826 585920 541828
rect -8576 535276 -7976 535278
rect 591900 535276 592500 535278
rect -8576 535254 592500 535276
rect -8576 535018 -8394 535254
rect -8158 535018 592082 535254
rect 592318 535018 592500 535254
rect -8576 534934 592500 535018
rect -8576 534698 -8394 534934
rect -8158 534698 592082 534934
rect 592318 534698 592500 534934
rect -8576 534676 592500 534698
rect -8576 534674 -7976 534676
rect 591900 534674 592500 534676
rect -6696 531676 -6096 531678
rect 590020 531676 590620 531678
rect -6696 531654 590620 531676
rect -6696 531418 -6514 531654
rect -6278 531418 590202 531654
rect 590438 531418 590620 531654
rect -6696 531334 590620 531418
rect -6696 531098 -6514 531334
rect -6278 531098 590202 531334
rect 590438 531098 590620 531334
rect -6696 531076 590620 531098
rect -6696 531074 -6096 531076
rect 590020 531074 590620 531076
rect -4816 528076 -4216 528078
rect 588140 528076 588740 528078
rect -4816 528054 588740 528076
rect -4816 527818 -4634 528054
rect -4398 527818 588322 528054
rect 588558 527818 588740 528054
rect -4816 527734 588740 527818
rect -4816 527498 -4634 527734
rect -4398 527498 588322 527734
rect 588558 527498 588740 527734
rect -4816 527476 588740 527498
rect -4816 527474 -4216 527476
rect 588140 527474 588740 527476
rect -2936 524428 -2336 524430
rect 586260 524428 586860 524430
rect -2936 524406 586860 524428
rect -2936 524170 -2754 524406
rect -2518 524170 586442 524406
rect 586678 524170 586860 524406
rect -2936 524086 586860 524170
rect -2936 523850 -2754 524086
rect -2518 523850 586442 524086
rect 586678 523850 586860 524086
rect -2936 523828 586860 523850
rect -2936 523826 -2336 523828
rect 586260 523826 586860 523828
rect -7636 517276 -7036 517278
rect 590960 517276 591560 517278
rect -8576 517254 592500 517276
rect -8576 517018 -7454 517254
rect -7218 517018 591142 517254
rect 591378 517018 592500 517254
rect -8576 516934 592500 517018
rect -8576 516698 -7454 516934
rect -7218 516698 591142 516934
rect 591378 516698 592500 516934
rect -8576 516676 592500 516698
rect -7636 516674 -7036 516676
rect 590960 516674 591560 516676
rect -5756 513676 -5156 513678
rect 589080 513676 589680 513678
rect -6696 513654 590620 513676
rect -6696 513418 -5574 513654
rect -5338 513418 589262 513654
rect 589498 513418 590620 513654
rect -6696 513334 590620 513418
rect -6696 513098 -5574 513334
rect -5338 513098 589262 513334
rect 589498 513098 590620 513334
rect -6696 513076 590620 513098
rect -5756 513074 -5156 513076
rect 589080 513074 589680 513076
rect -3876 510076 -3276 510078
rect 4404 510076 5004 510078
rect 580404 510076 581004 510078
rect 587200 510076 587800 510078
rect -4816 510054 588740 510076
rect -4816 509818 -3694 510054
rect -3458 509818 4586 510054
rect 4822 509818 580586 510054
rect 580822 509818 587382 510054
rect 587618 509818 588740 510054
rect -4816 509734 588740 509818
rect -4816 509498 -3694 509734
rect -3458 509498 4586 509734
rect 4822 509498 580586 509734
rect 580822 509498 587382 509734
rect 587618 509498 588740 509734
rect -4816 509476 588740 509498
rect -3876 509474 -3276 509476
rect 4404 509474 5004 509476
rect 580404 509474 581004 509476
rect 587200 509474 587800 509476
rect -1996 506428 -1396 506430
rect 804 506428 1404 506430
rect 585320 506428 585920 506430
rect -2936 506406 586860 506428
rect -2936 506170 -1814 506406
rect -1578 506170 986 506406
rect 1222 506170 585502 506406
rect 585738 506170 586860 506406
rect -2936 506086 586860 506170
rect -2936 505850 -1814 506086
rect -1578 505850 986 506086
rect 1222 505850 585502 506086
rect 585738 505850 586860 506086
rect -2936 505828 586860 505850
rect -1996 505826 -1396 505828
rect 804 505826 1404 505828
rect 585320 505826 585920 505828
rect -8576 499276 -7976 499278
rect 591900 499276 592500 499278
rect -8576 499254 592500 499276
rect -8576 499018 -8394 499254
rect -8158 499018 592082 499254
rect 592318 499018 592500 499254
rect -8576 498934 592500 499018
rect -8576 498698 -8394 498934
rect -8158 498698 592082 498934
rect 592318 498698 592500 498934
rect -8576 498676 592500 498698
rect -8576 498674 -7976 498676
rect 591900 498674 592500 498676
rect -6696 495676 -6096 495678
rect 590020 495676 590620 495678
rect -6696 495654 590620 495676
rect -6696 495418 -6514 495654
rect -6278 495418 590202 495654
rect 590438 495418 590620 495654
rect -6696 495334 590620 495418
rect -6696 495098 -6514 495334
rect -6278 495098 590202 495334
rect 590438 495098 590620 495334
rect -6696 495076 590620 495098
rect -6696 495074 -6096 495076
rect 590020 495074 590620 495076
rect -4816 492076 -4216 492078
rect 588140 492076 588740 492078
rect -4816 492054 588740 492076
rect -4816 491818 -4634 492054
rect -4398 491818 588322 492054
rect 588558 491818 588740 492054
rect -4816 491734 588740 491818
rect -4816 491498 -4634 491734
rect -4398 491498 588322 491734
rect 588558 491498 588740 491734
rect -4816 491476 588740 491498
rect -4816 491474 -4216 491476
rect 588140 491474 588740 491476
rect -2936 488428 -2336 488430
rect 586260 488428 586860 488430
rect -2936 488406 586860 488428
rect -2936 488170 -2754 488406
rect -2518 488170 586442 488406
rect 586678 488170 586860 488406
rect -2936 488086 586860 488170
rect -2936 487850 -2754 488086
rect -2518 487850 586442 488086
rect 586678 487850 586860 488086
rect -2936 487828 586860 487850
rect -2936 487826 -2336 487828
rect 586260 487826 586860 487828
rect -7636 481276 -7036 481278
rect 590960 481276 591560 481278
rect -8576 481254 592500 481276
rect -8576 481018 -7454 481254
rect -7218 481018 591142 481254
rect 591378 481018 592500 481254
rect -8576 480934 592500 481018
rect -8576 480698 -7454 480934
rect -7218 480698 591142 480934
rect 591378 480698 592500 480934
rect -8576 480676 592500 480698
rect -7636 480674 -7036 480676
rect 590960 480674 591560 480676
rect -5756 477676 -5156 477678
rect 589080 477676 589680 477678
rect -6696 477654 590620 477676
rect -6696 477418 -5574 477654
rect -5338 477418 589262 477654
rect 589498 477418 590620 477654
rect -6696 477334 590620 477418
rect -6696 477098 -5574 477334
rect -5338 477098 589262 477334
rect 589498 477098 590620 477334
rect -6696 477076 590620 477098
rect -5756 477074 -5156 477076
rect 589080 477074 589680 477076
rect -3876 474076 -3276 474078
rect 4404 474076 5004 474078
rect 580404 474076 581004 474078
rect 587200 474076 587800 474078
rect -4816 474054 588740 474076
rect -4816 473818 -3694 474054
rect -3458 473818 4586 474054
rect 4822 473818 580586 474054
rect 580822 473818 587382 474054
rect 587618 473818 588740 474054
rect -4816 473734 588740 473818
rect -4816 473498 -3694 473734
rect -3458 473498 4586 473734
rect 4822 473498 580586 473734
rect 580822 473498 587382 473734
rect 587618 473498 588740 473734
rect -4816 473476 588740 473498
rect -3876 473474 -3276 473476
rect 4404 473474 5004 473476
rect 580404 473474 581004 473476
rect 587200 473474 587800 473476
rect -1996 470428 -1396 470430
rect 804 470428 1404 470430
rect 585320 470428 585920 470430
rect -2936 470406 586860 470428
rect -2936 470170 -1814 470406
rect -1578 470170 986 470406
rect 1222 470170 585502 470406
rect 585738 470170 586860 470406
rect -2936 470086 586860 470170
rect -2936 469850 -1814 470086
rect -1578 469850 986 470086
rect 1222 469850 585502 470086
rect 585738 469850 586860 470086
rect -2936 469828 586860 469850
rect -1996 469826 -1396 469828
rect 804 469826 1404 469828
rect 585320 469826 585920 469828
rect -8576 463276 -7976 463278
rect 591900 463276 592500 463278
rect -8576 463254 592500 463276
rect -8576 463018 -8394 463254
rect -8158 463018 592082 463254
rect 592318 463018 592500 463254
rect -8576 462934 592500 463018
rect -8576 462698 -8394 462934
rect -8158 462698 592082 462934
rect 592318 462698 592500 462934
rect -8576 462676 592500 462698
rect -8576 462674 -7976 462676
rect 591900 462674 592500 462676
rect -6696 459676 -6096 459678
rect 590020 459676 590620 459678
rect -6696 459654 590620 459676
rect -6696 459418 -6514 459654
rect -6278 459418 590202 459654
rect 590438 459418 590620 459654
rect -6696 459334 590620 459418
rect -6696 459098 -6514 459334
rect -6278 459098 590202 459334
rect 590438 459098 590620 459334
rect -6696 459076 590620 459098
rect -6696 459074 -6096 459076
rect 590020 459074 590620 459076
rect -4816 456076 -4216 456078
rect 588140 456076 588740 456078
rect -4816 456054 588740 456076
rect -4816 455818 -4634 456054
rect -4398 455818 588322 456054
rect 588558 455818 588740 456054
rect -4816 455734 588740 455818
rect -4816 455498 -4634 455734
rect -4398 455498 588322 455734
rect 588558 455498 588740 455734
rect -4816 455476 588740 455498
rect -4816 455474 -4216 455476
rect 588140 455474 588740 455476
rect -2936 452428 -2336 452430
rect 586260 452428 586860 452430
rect -2936 452406 586860 452428
rect -2936 452170 -2754 452406
rect -2518 452170 586442 452406
rect 586678 452170 586860 452406
rect -2936 452086 586860 452170
rect -2936 451850 -2754 452086
rect -2518 451850 586442 452086
rect 586678 451850 586860 452086
rect -2936 451828 586860 451850
rect -2936 451826 -2336 451828
rect 586260 451826 586860 451828
rect -7636 445276 -7036 445278
rect 590960 445276 591560 445278
rect -8576 445254 592500 445276
rect -8576 445018 -7454 445254
rect -7218 445018 591142 445254
rect 591378 445018 592500 445254
rect -8576 444934 592500 445018
rect -8576 444698 -7454 444934
rect -7218 444698 591142 444934
rect 591378 444698 592500 444934
rect -8576 444676 592500 444698
rect -7636 444674 -7036 444676
rect 590960 444674 591560 444676
rect -5756 441676 -5156 441678
rect 589080 441676 589680 441678
rect -6696 441654 590620 441676
rect -6696 441418 -5574 441654
rect -5338 441418 589262 441654
rect 589498 441418 590620 441654
rect -6696 441334 590620 441418
rect -6696 441098 -5574 441334
rect -5338 441098 589262 441334
rect 589498 441098 590620 441334
rect -6696 441076 590620 441098
rect -5756 441074 -5156 441076
rect 589080 441074 589680 441076
rect -3876 438076 -3276 438078
rect 4404 438076 5004 438078
rect 580404 438076 581004 438078
rect 587200 438076 587800 438078
rect -4816 438054 588740 438076
rect -4816 437818 -3694 438054
rect -3458 437818 4586 438054
rect 4822 437818 580586 438054
rect 580822 437818 587382 438054
rect 587618 437818 588740 438054
rect -4816 437734 588740 437818
rect -4816 437498 -3694 437734
rect -3458 437498 4586 437734
rect 4822 437498 580586 437734
rect 580822 437498 587382 437734
rect 587618 437498 588740 437734
rect -4816 437476 588740 437498
rect -3876 437474 -3276 437476
rect 4404 437474 5004 437476
rect 580404 437474 581004 437476
rect 587200 437474 587800 437476
rect -1996 434428 -1396 434430
rect 804 434428 1404 434430
rect 585320 434428 585920 434430
rect -2936 434406 586860 434428
rect -2936 434170 -1814 434406
rect -1578 434170 986 434406
rect 1222 434170 585502 434406
rect 585738 434170 586860 434406
rect -2936 434086 586860 434170
rect -2936 433850 -1814 434086
rect -1578 433850 986 434086
rect 1222 433850 585502 434086
rect 585738 433850 586860 434086
rect -2936 433828 586860 433850
rect -1996 433826 -1396 433828
rect 804 433826 1404 433828
rect 585320 433826 585920 433828
rect -8576 427276 -7976 427278
rect 591900 427276 592500 427278
rect -8576 427254 592500 427276
rect -8576 427018 -8394 427254
rect -8158 427018 592082 427254
rect 592318 427018 592500 427254
rect -8576 426934 592500 427018
rect -8576 426698 -8394 426934
rect -8158 426698 592082 426934
rect 592318 426698 592500 426934
rect -8576 426676 592500 426698
rect -8576 426674 -7976 426676
rect 591900 426674 592500 426676
rect -6696 423676 -6096 423678
rect 590020 423676 590620 423678
rect -6696 423654 590620 423676
rect -6696 423418 -6514 423654
rect -6278 423418 590202 423654
rect 590438 423418 590620 423654
rect -6696 423334 590620 423418
rect -6696 423098 -6514 423334
rect -6278 423098 590202 423334
rect 590438 423098 590620 423334
rect -6696 423076 590620 423098
rect -6696 423074 -6096 423076
rect 590020 423074 590620 423076
rect -4816 420076 -4216 420078
rect 588140 420076 588740 420078
rect -4816 420054 588740 420076
rect -4816 419818 -4634 420054
rect -4398 419818 588322 420054
rect 588558 419818 588740 420054
rect -4816 419734 588740 419818
rect -4816 419498 -4634 419734
rect -4398 419498 588322 419734
rect 588558 419498 588740 419734
rect -4816 419476 588740 419498
rect -4816 419474 -4216 419476
rect 588140 419474 588740 419476
rect -2936 416428 -2336 416430
rect 586260 416428 586860 416430
rect -2936 416406 586860 416428
rect -2936 416170 -2754 416406
rect -2518 416170 586442 416406
rect 586678 416170 586860 416406
rect -2936 416086 586860 416170
rect -2936 415850 -2754 416086
rect -2518 415850 586442 416086
rect 586678 415850 586860 416086
rect -2936 415828 586860 415850
rect -2936 415826 -2336 415828
rect 586260 415826 586860 415828
rect -7636 409276 -7036 409278
rect 590960 409276 591560 409278
rect -8576 409254 592500 409276
rect -8576 409018 -7454 409254
rect -7218 409018 591142 409254
rect 591378 409018 592500 409254
rect -8576 408934 592500 409018
rect -8576 408698 -7454 408934
rect -7218 408698 591142 408934
rect 591378 408698 592500 408934
rect -8576 408676 592500 408698
rect -7636 408674 -7036 408676
rect 590960 408674 591560 408676
rect -5756 405676 -5156 405678
rect 589080 405676 589680 405678
rect -6696 405654 590620 405676
rect -6696 405418 -5574 405654
rect -5338 405418 589262 405654
rect 589498 405418 590620 405654
rect -6696 405334 590620 405418
rect -6696 405098 -5574 405334
rect -5338 405098 589262 405334
rect 589498 405098 590620 405334
rect -6696 405076 590620 405098
rect -5756 405074 -5156 405076
rect 589080 405074 589680 405076
rect -3876 402076 -3276 402078
rect 4404 402076 5004 402078
rect 580404 402076 581004 402078
rect 587200 402076 587800 402078
rect -4816 402054 588740 402076
rect -4816 401818 -3694 402054
rect -3458 401818 4586 402054
rect 4822 401818 580586 402054
rect 580822 401818 587382 402054
rect 587618 401818 588740 402054
rect -4816 401734 588740 401818
rect -4816 401498 -3694 401734
rect -3458 401498 4586 401734
rect 4822 401498 580586 401734
rect 580822 401498 587382 401734
rect 587618 401498 588740 401734
rect -4816 401476 588740 401498
rect -3876 401474 -3276 401476
rect 4404 401474 5004 401476
rect 580404 401474 581004 401476
rect 587200 401474 587800 401476
rect -1996 398428 -1396 398430
rect 804 398428 1404 398430
rect 585320 398428 585920 398430
rect -2936 398406 586860 398428
rect -2936 398170 -1814 398406
rect -1578 398170 986 398406
rect 1222 398170 585502 398406
rect 585738 398170 586860 398406
rect -2936 398086 586860 398170
rect -2936 397850 -1814 398086
rect -1578 397850 986 398086
rect 1222 397850 585502 398086
rect 585738 397850 586860 398086
rect -2936 397828 586860 397850
rect -1996 397826 -1396 397828
rect 804 397826 1404 397828
rect 585320 397826 585920 397828
rect -8576 391276 -7976 391278
rect 591900 391276 592500 391278
rect -8576 391254 592500 391276
rect -8576 391018 -8394 391254
rect -8158 391018 592082 391254
rect 592318 391018 592500 391254
rect -8576 390934 592500 391018
rect -8576 390698 -8394 390934
rect -8158 390698 592082 390934
rect 592318 390698 592500 390934
rect -8576 390676 592500 390698
rect -8576 390674 -7976 390676
rect 591900 390674 592500 390676
rect -6696 387676 -6096 387678
rect 590020 387676 590620 387678
rect -6696 387654 590620 387676
rect -6696 387418 -6514 387654
rect -6278 387418 590202 387654
rect 590438 387418 590620 387654
rect -6696 387334 590620 387418
rect -6696 387098 -6514 387334
rect -6278 387098 590202 387334
rect 590438 387098 590620 387334
rect -6696 387076 590620 387098
rect -6696 387074 -6096 387076
rect 590020 387074 590620 387076
rect -4816 384076 -4216 384078
rect 588140 384076 588740 384078
rect -4816 384054 588740 384076
rect -4816 383818 -4634 384054
rect -4398 383818 588322 384054
rect 588558 383818 588740 384054
rect -4816 383734 588740 383818
rect -4816 383498 -4634 383734
rect -4398 383498 588322 383734
rect 588558 383498 588740 383734
rect -4816 383476 588740 383498
rect -4816 383474 -4216 383476
rect 588140 383474 588740 383476
rect -2936 380428 -2336 380430
rect 586260 380428 586860 380430
rect -2936 380406 586860 380428
rect -2936 380170 -2754 380406
rect -2518 380170 586442 380406
rect 586678 380170 586860 380406
rect -2936 380086 586860 380170
rect -2936 379850 -2754 380086
rect -2518 379850 586442 380086
rect 586678 379850 586860 380086
rect -2936 379828 586860 379850
rect -2936 379826 -2336 379828
rect 586260 379826 586860 379828
rect -7636 373276 -7036 373278
rect 590960 373276 591560 373278
rect -8576 373254 592500 373276
rect -8576 373018 -7454 373254
rect -7218 373018 591142 373254
rect 591378 373018 592500 373254
rect -8576 372934 592500 373018
rect -8576 372698 -7454 372934
rect -7218 372698 591142 372934
rect 591378 372698 592500 372934
rect -8576 372676 592500 372698
rect -7636 372674 -7036 372676
rect 590960 372674 591560 372676
rect -5756 369676 -5156 369678
rect 589080 369676 589680 369678
rect -6696 369654 590620 369676
rect -6696 369418 -5574 369654
rect -5338 369418 589262 369654
rect 589498 369418 590620 369654
rect -6696 369334 590620 369418
rect -6696 369098 -5574 369334
rect -5338 369098 589262 369334
rect 589498 369098 590620 369334
rect -6696 369076 590620 369098
rect -5756 369074 -5156 369076
rect 589080 369074 589680 369076
rect -3876 366076 -3276 366078
rect 4404 366076 5004 366078
rect 580404 366076 581004 366078
rect 587200 366076 587800 366078
rect -4816 366054 588740 366076
rect -4816 365818 -3694 366054
rect -3458 365818 4586 366054
rect 4822 365818 580586 366054
rect 580822 365818 587382 366054
rect 587618 365818 588740 366054
rect -4816 365734 588740 365818
rect -4816 365498 -3694 365734
rect -3458 365498 4586 365734
rect 4822 365498 580586 365734
rect 580822 365498 587382 365734
rect 587618 365498 588740 365734
rect -4816 365476 588740 365498
rect -3876 365474 -3276 365476
rect 4404 365474 5004 365476
rect 580404 365474 581004 365476
rect 587200 365474 587800 365476
rect -1996 362428 -1396 362430
rect 804 362428 1404 362430
rect 585320 362428 585920 362430
rect -2936 362406 586860 362428
rect -2936 362170 -1814 362406
rect -1578 362170 986 362406
rect 1222 362170 585502 362406
rect 585738 362170 586860 362406
rect -2936 362086 586860 362170
rect -2936 361850 -1814 362086
rect -1578 361850 986 362086
rect 1222 361850 585502 362086
rect 585738 361850 586860 362086
rect -2936 361828 586860 361850
rect -1996 361826 -1396 361828
rect 804 361826 1404 361828
rect 585320 361826 585920 361828
rect -8576 355276 -7976 355278
rect 591900 355276 592500 355278
rect -8576 355254 592500 355276
rect -8576 355018 -8394 355254
rect -8158 355018 592082 355254
rect 592318 355018 592500 355254
rect -8576 354934 592500 355018
rect -8576 354698 -8394 354934
rect -8158 354698 592082 354934
rect 592318 354698 592500 354934
rect -8576 354676 592500 354698
rect -8576 354674 -7976 354676
rect 591900 354674 592500 354676
rect -6696 351676 -6096 351678
rect 590020 351676 590620 351678
rect -6696 351654 590620 351676
rect -6696 351418 -6514 351654
rect -6278 351418 590202 351654
rect 590438 351418 590620 351654
rect -6696 351334 590620 351418
rect -6696 351098 -6514 351334
rect -6278 351098 590202 351334
rect 590438 351098 590620 351334
rect -6696 351076 590620 351098
rect -6696 351074 -6096 351076
rect 590020 351074 590620 351076
rect -4816 348076 -4216 348078
rect 588140 348076 588740 348078
rect -4816 348054 588740 348076
rect -4816 347818 -4634 348054
rect -4398 347818 588322 348054
rect 588558 347818 588740 348054
rect -4816 347734 588740 347818
rect -4816 347498 -4634 347734
rect -4398 347498 588322 347734
rect 588558 347498 588740 347734
rect -4816 347476 588740 347498
rect -4816 347474 -4216 347476
rect 588140 347474 588740 347476
rect -2936 344428 -2336 344430
rect 586260 344428 586860 344430
rect -2936 344406 586860 344428
rect -2936 344170 -2754 344406
rect -2518 344170 586442 344406
rect 586678 344170 586860 344406
rect -2936 344086 586860 344170
rect -2936 343850 -2754 344086
rect -2518 343850 586442 344086
rect 586678 343850 586860 344086
rect -2936 343828 586860 343850
rect -2936 343826 -2336 343828
rect 586260 343826 586860 343828
rect -7636 337276 -7036 337278
rect 590960 337276 591560 337278
rect -8576 337254 592500 337276
rect -8576 337018 -7454 337254
rect -7218 337018 591142 337254
rect 591378 337018 592500 337254
rect -8576 336934 592500 337018
rect -8576 336698 -7454 336934
rect -7218 336698 591142 336934
rect 591378 336698 592500 336934
rect -8576 336676 592500 336698
rect -7636 336674 -7036 336676
rect 590960 336674 591560 336676
rect -5756 333676 -5156 333678
rect 589080 333676 589680 333678
rect -6696 333654 590620 333676
rect -6696 333418 -5574 333654
rect -5338 333418 589262 333654
rect 589498 333418 590620 333654
rect -6696 333334 590620 333418
rect -6696 333098 -5574 333334
rect -5338 333098 589262 333334
rect 589498 333098 590620 333334
rect -6696 333076 590620 333098
rect -5756 333074 -5156 333076
rect 589080 333074 589680 333076
rect -3876 330076 -3276 330078
rect 4404 330076 5004 330078
rect 580404 330076 581004 330078
rect 587200 330076 587800 330078
rect -4816 330054 588740 330076
rect -4816 329818 -3694 330054
rect -3458 329818 4586 330054
rect 4822 329818 580586 330054
rect 580822 329818 587382 330054
rect 587618 329818 588740 330054
rect -4816 329734 588740 329818
rect -4816 329498 -3694 329734
rect -3458 329498 4586 329734
rect 4822 329498 580586 329734
rect 580822 329498 587382 329734
rect 587618 329498 588740 329734
rect -4816 329476 588740 329498
rect -3876 329474 -3276 329476
rect 4404 329474 5004 329476
rect 580404 329474 581004 329476
rect 587200 329474 587800 329476
rect -1996 326428 -1396 326430
rect 804 326428 1404 326430
rect 585320 326428 585920 326430
rect -2936 326406 586860 326428
rect -2936 326170 -1814 326406
rect -1578 326170 986 326406
rect 1222 326170 585502 326406
rect 585738 326170 586860 326406
rect -2936 326086 586860 326170
rect -2936 325850 -1814 326086
rect -1578 325850 986 326086
rect 1222 325850 585502 326086
rect 585738 325850 586860 326086
rect -2936 325828 586860 325850
rect -1996 325826 -1396 325828
rect 804 325826 1404 325828
rect 585320 325826 585920 325828
rect -8576 319276 -7976 319278
rect 591900 319276 592500 319278
rect -8576 319254 592500 319276
rect -8576 319018 -8394 319254
rect -8158 319018 592082 319254
rect 592318 319018 592500 319254
rect -8576 318934 592500 319018
rect -8576 318698 -8394 318934
rect -8158 318698 592082 318934
rect 592318 318698 592500 318934
rect -8576 318676 592500 318698
rect -8576 318674 -7976 318676
rect 591900 318674 592500 318676
rect -6696 315676 -6096 315678
rect 590020 315676 590620 315678
rect -6696 315654 590620 315676
rect -6696 315418 -6514 315654
rect -6278 315418 590202 315654
rect 590438 315418 590620 315654
rect -6696 315334 590620 315418
rect -6696 315098 -6514 315334
rect -6278 315098 590202 315334
rect 590438 315098 590620 315334
rect -6696 315076 590620 315098
rect -6696 315074 -6096 315076
rect 590020 315074 590620 315076
rect -4816 312076 -4216 312078
rect 588140 312076 588740 312078
rect -4816 312054 588740 312076
rect -4816 311818 -4634 312054
rect -4398 311818 588322 312054
rect 588558 311818 588740 312054
rect -4816 311734 588740 311818
rect -4816 311498 -4634 311734
rect -4398 311498 588322 311734
rect 588558 311498 588740 311734
rect -4816 311476 588740 311498
rect -4816 311474 -4216 311476
rect 588140 311474 588740 311476
rect -2936 308428 -2336 308430
rect 586260 308428 586860 308430
rect -2936 308406 586860 308428
rect -2936 308170 -2754 308406
rect -2518 308170 586442 308406
rect 586678 308170 586860 308406
rect -2936 308086 586860 308170
rect -2936 307850 -2754 308086
rect -2518 307850 586442 308086
rect 586678 307850 586860 308086
rect -2936 307828 586860 307850
rect -2936 307826 -2336 307828
rect 586260 307826 586860 307828
rect -7636 301276 -7036 301278
rect 590960 301276 591560 301278
rect -8576 301254 592500 301276
rect -8576 301018 -7454 301254
rect -7218 301018 591142 301254
rect 591378 301018 592500 301254
rect -8576 300934 592500 301018
rect -8576 300698 -7454 300934
rect -7218 300698 591142 300934
rect 591378 300698 592500 300934
rect -8576 300676 592500 300698
rect -7636 300674 -7036 300676
rect 590960 300674 591560 300676
rect -5756 297676 -5156 297678
rect 589080 297676 589680 297678
rect -6696 297654 590620 297676
rect -6696 297418 -5574 297654
rect -5338 297418 589262 297654
rect 589498 297418 590620 297654
rect -6696 297334 590620 297418
rect -6696 297098 -5574 297334
rect -5338 297098 589262 297334
rect 589498 297098 590620 297334
rect -6696 297076 590620 297098
rect -5756 297074 -5156 297076
rect 589080 297074 589680 297076
rect -3876 294076 -3276 294078
rect 4404 294076 5004 294078
rect 580404 294076 581004 294078
rect 587200 294076 587800 294078
rect -4816 294054 588740 294076
rect -4816 293818 -3694 294054
rect -3458 293818 4586 294054
rect 4822 293818 580586 294054
rect 580822 293818 587382 294054
rect 587618 293818 588740 294054
rect -4816 293734 588740 293818
rect -4816 293498 -3694 293734
rect -3458 293498 4586 293734
rect 4822 293498 580586 293734
rect 580822 293498 587382 293734
rect 587618 293498 588740 293734
rect -4816 293476 588740 293498
rect -3876 293474 -3276 293476
rect 4404 293474 5004 293476
rect 580404 293474 581004 293476
rect 587200 293474 587800 293476
rect -1996 290428 -1396 290430
rect 804 290428 1404 290430
rect 585320 290428 585920 290430
rect -2936 290406 586860 290428
rect -2936 290170 -1814 290406
rect -1578 290170 986 290406
rect 1222 290170 585502 290406
rect 585738 290170 586860 290406
rect -2936 290086 586860 290170
rect -2936 289850 -1814 290086
rect -1578 289850 986 290086
rect 1222 289850 585502 290086
rect 585738 289850 586860 290086
rect -2936 289828 586860 289850
rect -1996 289826 -1396 289828
rect 804 289826 1404 289828
rect 585320 289826 585920 289828
rect -8576 283276 -7976 283278
rect 591900 283276 592500 283278
rect -8576 283254 592500 283276
rect -8576 283018 -8394 283254
rect -8158 283018 592082 283254
rect 592318 283018 592500 283254
rect -8576 282934 592500 283018
rect -8576 282698 -8394 282934
rect -8158 282698 592082 282934
rect 592318 282698 592500 282934
rect -8576 282676 592500 282698
rect -8576 282674 -7976 282676
rect 591900 282674 592500 282676
rect -6696 279676 -6096 279678
rect 590020 279676 590620 279678
rect -6696 279654 590620 279676
rect -6696 279418 -6514 279654
rect -6278 279418 590202 279654
rect 590438 279418 590620 279654
rect -6696 279334 590620 279418
rect -6696 279098 -6514 279334
rect -6278 279098 590202 279334
rect 590438 279098 590620 279334
rect -6696 279076 590620 279098
rect -6696 279074 -6096 279076
rect 590020 279074 590620 279076
rect -4816 276076 -4216 276078
rect 588140 276076 588740 276078
rect -4816 276054 588740 276076
rect -4816 275818 -4634 276054
rect -4398 275818 588322 276054
rect 588558 275818 588740 276054
rect -4816 275734 588740 275818
rect -4816 275498 -4634 275734
rect -4398 275498 588322 275734
rect 588558 275498 588740 275734
rect -4816 275476 588740 275498
rect -4816 275474 -4216 275476
rect 588140 275474 588740 275476
rect -2936 272428 -2336 272430
rect 586260 272428 586860 272430
rect -2936 272406 586860 272428
rect -2936 272170 -2754 272406
rect -2518 272170 586442 272406
rect 586678 272170 586860 272406
rect -2936 272086 586860 272170
rect -2936 271850 -2754 272086
rect -2518 271850 586442 272086
rect 586678 271850 586860 272086
rect -2936 271828 586860 271850
rect -2936 271826 -2336 271828
rect 586260 271826 586860 271828
rect -7636 265276 -7036 265278
rect 590960 265276 591560 265278
rect -8576 265254 592500 265276
rect -8576 265018 -7454 265254
rect -7218 265018 591142 265254
rect 591378 265018 592500 265254
rect -8576 264934 592500 265018
rect -8576 264698 -7454 264934
rect -7218 264698 591142 264934
rect 591378 264698 592500 264934
rect -8576 264676 592500 264698
rect -7636 264674 -7036 264676
rect 590960 264674 591560 264676
rect -5756 261676 -5156 261678
rect 589080 261676 589680 261678
rect -6696 261654 590620 261676
rect -6696 261418 -5574 261654
rect -5338 261418 589262 261654
rect 589498 261418 590620 261654
rect -6696 261334 590620 261418
rect -6696 261098 -5574 261334
rect -5338 261098 589262 261334
rect 589498 261098 590620 261334
rect -6696 261076 590620 261098
rect -5756 261074 -5156 261076
rect 589080 261074 589680 261076
rect -3876 258076 -3276 258078
rect 4404 258076 5004 258078
rect 580404 258076 581004 258078
rect 587200 258076 587800 258078
rect -4816 258054 588740 258076
rect -4816 257818 -3694 258054
rect -3458 257818 4586 258054
rect 4822 257818 580586 258054
rect 580822 257818 587382 258054
rect 587618 257818 588740 258054
rect -4816 257734 588740 257818
rect -4816 257498 -3694 257734
rect -3458 257498 4586 257734
rect 4822 257498 580586 257734
rect 580822 257498 587382 257734
rect 587618 257498 588740 257734
rect -4816 257476 588740 257498
rect -3876 257474 -3276 257476
rect 4404 257474 5004 257476
rect 580404 257474 581004 257476
rect 587200 257474 587800 257476
rect -1996 254428 -1396 254430
rect 804 254428 1404 254430
rect 585320 254428 585920 254430
rect -2936 254406 586860 254428
rect -2936 254170 -1814 254406
rect -1578 254170 986 254406
rect 1222 254170 585502 254406
rect 585738 254170 586860 254406
rect -2936 254086 586860 254170
rect -2936 253850 -1814 254086
rect -1578 253850 986 254086
rect 1222 253850 585502 254086
rect 585738 253850 586860 254086
rect -2936 253828 586860 253850
rect -1996 253826 -1396 253828
rect 804 253826 1404 253828
rect 585320 253826 585920 253828
rect -8576 247276 -7976 247278
rect 591900 247276 592500 247278
rect -8576 247254 592500 247276
rect -8576 247018 -8394 247254
rect -8158 247018 592082 247254
rect 592318 247018 592500 247254
rect -8576 246934 592500 247018
rect -8576 246698 -8394 246934
rect -8158 246698 592082 246934
rect 592318 246698 592500 246934
rect -8576 246676 592500 246698
rect -8576 246674 -7976 246676
rect 591900 246674 592500 246676
rect -6696 243676 -6096 243678
rect 590020 243676 590620 243678
rect -6696 243654 590620 243676
rect -6696 243418 -6514 243654
rect -6278 243418 590202 243654
rect 590438 243418 590620 243654
rect -6696 243334 590620 243418
rect -6696 243098 -6514 243334
rect -6278 243098 590202 243334
rect 590438 243098 590620 243334
rect -6696 243076 590620 243098
rect -6696 243074 -6096 243076
rect 590020 243074 590620 243076
rect -4816 240076 -4216 240078
rect 588140 240076 588740 240078
rect -4816 240054 588740 240076
rect -4816 239818 -4634 240054
rect -4398 239818 588322 240054
rect 588558 239818 588740 240054
rect -4816 239734 588740 239818
rect -4816 239498 -4634 239734
rect -4398 239498 588322 239734
rect 588558 239498 588740 239734
rect -4816 239476 588740 239498
rect -4816 239474 -4216 239476
rect 588140 239474 588740 239476
rect -2936 236428 -2336 236430
rect 586260 236428 586860 236430
rect -2936 236406 586860 236428
rect -2936 236170 -2754 236406
rect -2518 236170 586442 236406
rect 586678 236170 586860 236406
rect -2936 236086 586860 236170
rect -2936 235850 -2754 236086
rect -2518 235850 586442 236086
rect 586678 235850 586860 236086
rect -2936 235828 586860 235850
rect -2936 235826 -2336 235828
rect 586260 235826 586860 235828
rect -7636 229276 -7036 229278
rect 590960 229276 591560 229278
rect -8576 229254 592500 229276
rect -8576 229018 -7454 229254
rect -7218 229018 591142 229254
rect 591378 229018 592500 229254
rect -8576 228934 592500 229018
rect -8576 228698 -7454 228934
rect -7218 228698 591142 228934
rect 591378 228698 592500 228934
rect -8576 228676 592500 228698
rect -7636 228674 -7036 228676
rect 590960 228674 591560 228676
rect -5756 225676 -5156 225678
rect 589080 225676 589680 225678
rect -6696 225654 590620 225676
rect -6696 225418 -5574 225654
rect -5338 225418 589262 225654
rect 589498 225418 590620 225654
rect -6696 225334 590620 225418
rect -6696 225098 -5574 225334
rect -5338 225098 589262 225334
rect 589498 225098 590620 225334
rect -6696 225076 590620 225098
rect -5756 225074 -5156 225076
rect 589080 225074 589680 225076
rect -3876 222076 -3276 222078
rect 4404 222076 5004 222078
rect 580404 222076 581004 222078
rect 587200 222076 587800 222078
rect -4816 222054 588740 222076
rect -4816 221818 -3694 222054
rect -3458 221818 4586 222054
rect 4822 221818 580586 222054
rect 580822 221818 587382 222054
rect 587618 221818 588740 222054
rect -4816 221734 588740 221818
rect -4816 221498 -3694 221734
rect -3458 221498 4586 221734
rect 4822 221498 580586 221734
rect 580822 221498 587382 221734
rect 587618 221498 588740 221734
rect -4816 221476 588740 221498
rect -3876 221474 -3276 221476
rect 4404 221474 5004 221476
rect 580404 221474 581004 221476
rect 587200 221474 587800 221476
rect -1996 218428 -1396 218430
rect 804 218428 1404 218430
rect 585320 218428 585920 218430
rect -2936 218406 586860 218428
rect -2936 218170 -1814 218406
rect -1578 218170 986 218406
rect 1222 218170 585502 218406
rect 585738 218170 586860 218406
rect -2936 218086 586860 218170
rect -2936 217850 -1814 218086
rect -1578 217850 986 218086
rect 1222 217850 585502 218086
rect 585738 217850 586860 218086
rect -2936 217828 586860 217850
rect -1996 217826 -1396 217828
rect 804 217826 1404 217828
rect 585320 217826 585920 217828
rect -8576 211276 -7976 211278
rect 591900 211276 592500 211278
rect -8576 211254 592500 211276
rect -8576 211018 -8394 211254
rect -8158 211018 592082 211254
rect 592318 211018 592500 211254
rect -8576 210934 592500 211018
rect -8576 210698 -8394 210934
rect -8158 210698 592082 210934
rect 592318 210698 592500 210934
rect -8576 210676 592500 210698
rect -8576 210674 -7976 210676
rect 591900 210674 592500 210676
rect -6696 207676 -6096 207678
rect 590020 207676 590620 207678
rect -6696 207654 590620 207676
rect -6696 207418 -6514 207654
rect -6278 207418 590202 207654
rect 590438 207418 590620 207654
rect -6696 207334 590620 207418
rect -6696 207098 -6514 207334
rect -6278 207098 590202 207334
rect 590438 207098 590620 207334
rect -6696 207076 590620 207098
rect -6696 207074 -6096 207076
rect 590020 207074 590620 207076
rect -4816 204076 -4216 204078
rect 588140 204076 588740 204078
rect -4816 204054 588740 204076
rect -4816 203818 -4634 204054
rect -4398 203818 588322 204054
rect 588558 203818 588740 204054
rect -4816 203734 588740 203818
rect -4816 203498 -4634 203734
rect -4398 203498 588322 203734
rect 588558 203498 588740 203734
rect -4816 203476 588740 203498
rect -4816 203474 -4216 203476
rect 588140 203474 588740 203476
rect -2936 200428 -2336 200430
rect 586260 200428 586860 200430
rect -2936 200406 586860 200428
rect -2936 200170 -2754 200406
rect -2518 200170 586442 200406
rect 586678 200170 586860 200406
rect -2936 200086 586860 200170
rect -2936 199850 -2754 200086
rect -2518 199850 586442 200086
rect 586678 199850 586860 200086
rect -2936 199828 586860 199850
rect -2936 199826 -2336 199828
rect 586260 199826 586860 199828
rect -7636 193276 -7036 193278
rect 590960 193276 591560 193278
rect -8576 193254 592500 193276
rect -8576 193018 -7454 193254
rect -7218 193018 591142 193254
rect 591378 193018 592500 193254
rect -8576 192934 592500 193018
rect -8576 192698 -7454 192934
rect -7218 192698 591142 192934
rect 591378 192698 592500 192934
rect -8576 192676 592500 192698
rect -7636 192674 -7036 192676
rect 590960 192674 591560 192676
rect -5756 189676 -5156 189678
rect 589080 189676 589680 189678
rect -6696 189654 590620 189676
rect -6696 189418 -5574 189654
rect -5338 189418 589262 189654
rect 589498 189418 590620 189654
rect -6696 189334 590620 189418
rect -6696 189098 -5574 189334
rect -5338 189098 589262 189334
rect 589498 189098 590620 189334
rect -6696 189076 590620 189098
rect -5756 189074 -5156 189076
rect 589080 189074 589680 189076
rect -3876 186076 -3276 186078
rect 4404 186076 5004 186078
rect 580404 186076 581004 186078
rect 587200 186076 587800 186078
rect -4816 186054 588740 186076
rect -4816 185818 -3694 186054
rect -3458 185818 4586 186054
rect 4822 185818 580586 186054
rect 580822 185818 587382 186054
rect 587618 185818 588740 186054
rect -4816 185734 588740 185818
rect -4816 185498 -3694 185734
rect -3458 185498 4586 185734
rect 4822 185498 580586 185734
rect 580822 185498 587382 185734
rect 587618 185498 588740 185734
rect -4816 185476 588740 185498
rect -3876 185474 -3276 185476
rect 4404 185474 5004 185476
rect 580404 185474 581004 185476
rect 587200 185474 587800 185476
rect -1996 182428 -1396 182430
rect 804 182428 1404 182430
rect 585320 182428 585920 182430
rect -2936 182406 586860 182428
rect -2936 182170 -1814 182406
rect -1578 182170 986 182406
rect 1222 182170 585502 182406
rect 585738 182170 586860 182406
rect -2936 182086 586860 182170
rect -2936 181850 -1814 182086
rect -1578 181850 986 182086
rect 1222 181850 585502 182086
rect 585738 181850 586860 182086
rect -2936 181828 586860 181850
rect -1996 181826 -1396 181828
rect 804 181826 1404 181828
rect 585320 181826 585920 181828
rect -8576 175276 -7976 175278
rect 591900 175276 592500 175278
rect -8576 175254 592500 175276
rect -8576 175018 -8394 175254
rect -8158 175018 592082 175254
rect 592318 175018 592500 175254
rect -8576 174934 592500 175018
rect -8576 174698 -8394 174934
rect -8158 174698 592082 174934
rect 592318 174698 592500 174934
rect -8576 174676 592500 174698
rect -8576 174674 -7976 174676
rect 591900 174674 592500 174676
rect -6696 171676 -6096 171678
rect 590020 171676 590620 171678
rect -6696 171654 590620 171676
rect -6696 171418 -6514 171654
rect -6278 171418 590202 171654
rect 590438 171418 590620 171654
rect -6696 171334 590620 171418
rect -6696 171098 -6514 171334
rect -6278 171098 590202 171334
rect 590438 171098 590620 171334
rect -6696 171076 590620 171098
rect -6696 171074 -6096 171076
rect 590020 171074 590620 171076
rect -4816 168076 -4216 168078
rect 588140 168076 588740 168078
rect -4816 168054 588740 168076
rect -4816 167818 -4634 168054
rect -4398 167818 588322 168054
rect 588558 167818 588740 168054
rect -4816 167734 588740 167818
rect -4816 167498 -4634 167734
rect -4398 167498 588322 167734
rect 588558 167498 588740 167734
rect -4816 167476 588740 167498
rect -4816 167474 -4216 167476
rect 588140 167474 588740 167476
rect -2936 164428 -2336 164430
rect 586260 164428 586860 164430
rect -2936 164406 586860 164428
rect -2936 164170 -2754 164406
rect -2518 164170 586442 164406
rect 586678 164170 586860 164406
rect -2936 164086 586860 164170
rect -2936 163850 -2754 164086
rect -2518 163850 586442 164086
rect 586678 163850 586860 164086
rect -2936 163828 586860 163850
rect -2936 163826 -2336 163828
rect 586260 163826 586860 163828
rect -7636 157276 -7036 157278
rect 590960 157276 591560 157278
rect -8576 157254 592500 157276
rect -8576 157018 -7454 157254
rect -7218 157018 591142 157254
rect 591378 157018 592500 157254
rect -8576 156934 592500 157018
rect -8576 156698 -7454 156934
rect -7218 156698 591142 156934
rect 591378 156698 592500 156934
rect -8576 156676 592500 156698
rect -7636 156674 -7036 156676
rect 590960 156674 591560 156676
rect -5756 153676 -5156 153678
rect 589080 153676 589680 153678
rect -6696 153654 590620 153676
rect -6696 153418 -5574 153654
rect -5338 153418 589262 153654
rect 589498 153418 590620 153654
rect -6696 153334 590620 153418
rect -6696 153098 -5574 153334
rect -5338 153098 589262 153334
rect 589498 153098 590620 153334
rect -6696 153076 590620 153098
rect -5756 153074 -5156 153076
rect 589080 153074 589680 153076
rect -3876 150076 -3276 150078
rect 4404 150076 5004 150078
rect 580404 150076 581004 150078
rect 587200 150076 587800 150078
rect -4816 150054 588740 150076
rect -4816 149818 -3694 150054
rect -3458 149818 4586 150054
rect 4822 149818 580586 150054
rect 580822 149818 587382 150054
rect 587618 149818 588740 150054
rect -4816 149734 588740 149818
rect -4816 149498 -3694 149734
rect -3458 149498 4586 149734
rect 4822 149498 580586 149734
rect 580822 149498 587382 149734
rect 587618 149498 588740 149734
rect -4816 149476 588740 149498
rect -3876 149474 -3276 149476
rect 4404 149474 5004 149476
rect 580404 149474 581004 149476
rect 587200 149474 587800 149476
rect -1996 146428 -1396 146430
rect 804 146428 1404 146430
rect 585320 146428 585920 146430
rect -2936 146406 586860 146428
rect -2936 146170 -1814 146406
rect -1578 146170 986 146406
rect 1222 146170 585502 146406
rect 585738 146170 586860 146406
rect -2936 146086 586860 146170
rect -2936 145850 -1814 146086
rect -1578 145850 986 146086
rect 1222 145850 585502 146086
rect 585738 145850 586860 146086
rect -2936 145828 586860 145850
rect -1996 145826 -1396 145828
rect 804 145826 1404 145828
rect 585320 145826 585920 145828
rect -8576 139276 -7976 139278
rect 591900 139276 592500 139278
rect -8576 139254 592500 139276
rect -8576 139018 -8394 139254
rect -8158 139018 592082 139254
rect 592318 139018 592500 139254
rect -8576 138934 592500 139018
rect -8576 138698 -8394 138934
rect -8158 138698 592082 138934
rect 592318 138698 592500 138934
rect -8576 138676 592500 138698
rect -8576 138674 -7976 138676
rect 591900 138674 592500 138676
rect -6696 135676 -6096 135678
rect 590020 135676 590620 135678
rect -6696 135654 590620 135676
rect -6696 135418 -6514 135654
rect -6278 135418 590202 135654
rect 590438 135418 590620 135654
rect -6696 135334 590620 135418
rect -6696 135098 -6514 135334
rect -6278 135098 590202 135334
rect 590438 135098 590620 135334
rect -6696 135076 590620 135098
rect -6696 135074 -6096 135076
rect 590020 135074 590620 135076
rect -4816 132076 -4216 132078
rect 588140 132076 588740 132078
rect -4816 132054 588740 132076
rect -4816 131818 -4634 132054
rect -4398 131818 588322 132054
rect 588558 131818 588740 132054
rect -4816 131734 588740 131818
rect -4816 131498 -4634 131734
rect -4398 131498 588322 131734
rect 588558 131498 588740 131734
rect -4816 131476 588740 131498
rect -4816 131474 -4216 131476
rect 588140 131474 588740 131476
rect -2936 128428 -2336 128430
rect 586260 128428 586860 128430
rect -2936 128406 586860 128428
rect -2936 128170 -2754 128406
rect -2518 128170 586442 128406
rect 586678 128170 586860 128406
rect -2936 128086 586860 128170
rect -2936 127850 -2754 128086
rect -2518 127850 586442 128086
rect 586678 127850 586860 128086
rect -2936 127828 586860 127850
rect -2936 127826 -2336 127828
rect 586260 127826 586860 127828
rect -7636 121276 -7036 121278
rect 590960 121276 591560 121278
rect -8576 121254 592500 121276
rect -8576 121018 -7454 121254
rect -7218 121018 591142 121254
rect 591378 121018 592500 121254
rect -8576 120934 592500 121018
rect -8576 120698 -7454 120934
rect -7218 120698 591142 120934
rect 591378 120698 592500 120934
rect -8576 120676 592500 120698
rect -7636 120674 -7036 120676
rect 590960 120674 591560 120676
rect -5756 117676 -5156 117678
rect 589080 117676 589680 117678
rect -6696 117654 590620 117676
rect -6696 117418 -5574 117654
rect -5338 117418 589262 117654
rect 589498 117418 590620 117654
rect -6696 117334 590620 117418
rect -6696 117098 -5574 117334
rect -5338 117098 589262 117334
rect 589498 117098 590620 117334
rect -6696 117076 590620 117098
rect -5756 117074 -5156 117076
rect 589080 117074 589680 117076
rect -3876 114076 -3276 114078
rect 4404 114076 5004 114078
rect 580404 114076 581004 114078
rect 587200 114076 587800 114078
rect -4816 114054 588740 114076
rect -4816 113818 -3694 114054
rect -3458 113818 4586 114054
rect 4822 113818 580586 114054
rect 580822 113818 587382 114054
rect 587618 113818 588740 114054
rect -4816 113734 588740 113818
rect -4816 113498 -3694 113734
rect -3458 113498 4586 113734
rect 4822 113498 580586 113734
rect 580822 113498 587382 113734
rect 587618 113498 588740 113734
rect -4816 113476 588740 113498
rect -3876 113474 -3276 113476
rect 4404 113474 5004 113476
rect 580404 113474 581004 113476
rect 587200 113474 587800 113476
rect -1996 110428 -1396 110430
rect 804 110428 1404 110430
rect 585320 110428 585920 110430
rect -2936 110406 586860 110428
rect -2936 110170 -1814 110406
rect -1578 110170 986 110406
rect 1222 110170 585502 110406
rect 585738 110170 586860 110406
rect -2936 110086 586860 110170
rect -2936 109850 -1814 110086
rect -1578 109850 986 110086
rect 1222 109850 585502 110086
rect 585738 109850 586860 110086
rect -2936 109828 586860 109850
rect -1996 109826 -1396 109828
rect 804 109826 1404 109828
rect 585320 109826 585920 109828
rect -8576 103276 -7976 103278
rect 591900 103276 592500 103278
rect -8576 103254 592500 103276
rect -8576 103018 -8394 103254
rect -8158 103018 592082 103254
rect 592318 103018 592500 103254
rect -8576 102934 592500 103018
rect -8576 102698 -8394 102934
rect -8158 102698 592082 102934
rect 592318 102698 592500 102934
rect -8576 102676 592500 102698
rect -8576 102674 -7976 102676
rect 591900 102674 592500 102676
rect -6696 99676 -6096 99678
rect 590020 99676 590620 99678
rect -6696 99654 590620 99676
rect -6696 99418 -6514 99654
rect -6278 99418 590202 99654
rect 590438 99418 590620 99654
rect -6696 99334 590620 99418
rect -6696 99098 -6514 99334
rect -6278 99098 590202 99334
rect 590438 99098 590620 99334
rect -6696 99076 590620 99098
rect -6696 99074 -6096 99076
rect 590020 99074 590620 99076
rect -4816 96076 -4216 96078
rect 588140 96076 588740 96078
rect -4816 96054 588740 96076
rect -4816 95818 -4634 96054
rect -4398 95818 588322 96054
rect 588558 95818 588740 96054
rect -4816 95734 588740 95818
rect -4816 95498 -4634 95734
rect -4398 95498 588322 95734
rect 588558 95498 588740 95734
rect -4816 95476 588740 95498
rect -4816 95474 -4216 95476
rect 588140 95474 588740 95476
rect -2936 92428 -2336 92430
rect 586260 92428 586860 92430
rect -2936 92406 586860 92428
rect -2936 92170 -2754 92406
rect -2518 92170 586442 92406
rect 586678 92170 586860 92406
rect -2936 92086 586860 92170
rect -2936 91850 -2754 92086
rect -2518 91850 586442 92086
rect 586678 91850 586860 92086
rect -2936 91828 586860 91850
rect -2936 91826 -2336 91828
rect 586260 91826 586860 91828
rect -7636 85276 -7036 85278
rect 590960 85276 591560 85278
rect -8576 85254 592500 85276
rect -8576 85018 -7454 85254
rect -7218 85018 591142 85254
rect 591378 85018 592500 85254
rect -8576 84934 592500 85018
rect -8576 84698 -7454 84934
rect -7218 84698 591142 84934
rect 591378 84698 592500 84934
rect -8576 84676 592500 84698
rect -7636 84674 -7036 84676
rect 590960 84674 591560 84676
rect -5756 81676 -5156 81678
rect 589080 81676 589680 81678
rect -6696 81654 590620 81676
rect -6696 81418 -5574 81654
rect -5338 81418 589262 81654
rect 589498 81418 590620 81654
rect -6696 81334 590620 81418
rect -6696 81098 -5574 81334
rect -5338 81098 589262 81334
rect 589498 81098 590620 81334
rect -6696 81076 590620 81098
rect -5756 81074 -5156 81076
rect 589080 81074 589680 81076
rect -3876 78076 -3276 78078
rect 4404 78076 5004 78078
rect 580404 78076 581004 78078
rect 587200 78076 587800 78078
rect -4816 78054 588740 78076
rect -4816 77818 -3694 78054
rect -3458 77818 4586 78054
rect 4822 77818 580586 78054
rect 580822 77818 587382 78054
rect 587618 77818 588740 78054
rect -4816 77734 588740 77818
rect -4816 77498 -3694 77734
rect -3458 77498 4586 77734
rect 4822 77498 580586 77734
rect 580822 77498 587382 77734
rect 587618 77498 588740 77734
rect -4816 77476 588740 77498
rect -3876 77474 -3276 77476
rect 4404 77474 5004 77476
rect 580404 77474 581004 77476
rect 587200 77474 587800 77476
rect -1996 74428 -1396 74430
rect 804 74428 1404 74430
rect 585320 74428 585920 74430
rect -2936 74406 586860 74428
rect -2936 74170 -1814 74406
rect -1578 74170 986 74406
rect 1222 74170 585502 74406
rect 585738 74170 586860 74406
rect -2936 74086 586860 74170
rect -2936 73850 -1814 74086
rect -1578 73850 986 74086
rect 1222 73850 585502 74086
rect 585738 73850 586860 74086
rect -2936 73828 586860 73850
rect -1996 73826 -1396 73828
rect 804 73826 1404 73828
rect 585320 73826 585920 73828
rect -8576 67276 -7976 67278
rect 591900 67276 592500 67278
rect -8576 67254 592500 67276
rect -8576 67018 -8394 67254
rect -8158 67018 592082 67254
rect 592318 67018 592500 67254
rect -8576 66934 592500 67018
rect -8576 66698 -8394 66934
rect -8158 66698 592082 66934
rect 592318 66698 592500 66934
rect -8576 66676 592500 66698
rect -8576 66674 -7976 66676
rect 591900 66674 592500 66676
rect -6696 63676 -6096 63678
rect 590020 63676 590620 63678
rect -6696 63654 590620 63676
rect -6696 63418 -6514 63654
rect -6278 63418 590202 63654
rect 590438 63418 590620 63654
rect -6696 63334 590620 63418
rect -6696 63098 -6514 63334
rect -6278 63098 590202 63334
rect 590438 63098 590620 63334
rect -6696 63076 590620 63098
rect -6696 63074 -6096 63076
rect 590020 63074 590620 63076
rect -4816 60076 -4216 60078
rect 588140 60076 588740 60078
rect -4816 60054 588740 60076
rect -4816 59818 -4634 60054
rect -4398 59818 588322 60054
rect 588558 59818 588740 60054
rect -4816 59734 588740 59818
rect -4816 59498 -4634 59734
rect -4398 59498 588322 59734
rect 588558 59498 588740 59734
rect -4816 59476 588740 59498
rect -4816 59474 -4216 59476
rect 588140 59474 588740 59476
rect -2936 56428 -2336 56430
rect 586260 56428 586860 56430
rect -2936 56406 586860 56428
rect -2936 56170 -2754 56406
rect -2518 56170 586442 56406
rect 586678 56170 586860 56406
rect -2936 56086 586860 56170
rect -2936 55850 -2754 56086
rect -2518 55850 586442 56086
rect 586678 55850 586860 56086
rect -2936 55828 586860 55850
rect -2936 55826 -2336 55828
rect 586260 55826 586860 55828
rect -7636 49276 -7036 49278
rect 590960 49276 591560 49278
rect -8576 49254 592500 49276
rect -8576 49018 -7454 49254
rect -7218 49018 591142 49254
rect 591378 49018 592500 49254
rect -8576 48934 592500 49018
rect -8576 48698 -7454 48934
rect -7218 48698 591142 48934
rect 591378 48698 592500 48934
rect -8576 48676 592500 48698
rect -7636 48674 -7036 48676
rect 590960 48674 591560 48676
rect -5756 45676 -5156 45678
rect 589080 45676 589680 45678
rect -6696 45654 590620 45676
rect -6696 45418 -5574 45654
rect -5338 45418 589262 45654
rect 589498 45418 590620 45654
rect -6696 45334 590620 45418
rect -6696 45098 -5574 45334
rect -5338 45098 589262 45334
rect 589498 45098 590620 45334
rect -6696 45076 590620 45098
rect -5756 45074 -5156 45076
rect 589080 45074 589680 45076
rect -3876 42076 -3276 42078
rect 4404 42076 5004 42078
rect 580404 42076 581004 42078
rect 587200 42076 587800 42078
rect -4816 42054 588740 42076
rect -4816 41818 -3694 42054
rect -3458 41818 4586 42054
rect 4822 41818 580586 42054
rect 580822 41818 587382 42054
rect 587618 41818 588740 42054
rect -4816 41734 588740 41818
rect -4816 41498 -3694 41734
rect -3458 41498 4586 41734
rect 4822 41498 580586 41734
rect 580822 41498 587382 41734
rect 587618 41498 588740 41734
rect -4816 41476 588740 41498
rect -3876 41474 -3276 41476
rect 4404 41474 5004 41476
rect 580404 41474 581004 41476
rect 587200 41474 587800 41476
rect -1996 38428 -1396 38430
rect 804 38428 1404 38430
rect 585320 38428 585920 38430
rect -2936 38406 586860 38428
rect -2936 38170 -1814 38406
rect -1578 38170 986 38406
rect 1222 38170 585502 38406
rect 585738 38170 586860 38406
rect -2936 38086 586860 38170
rect -2936 37850 -1814 38086
rect -1578 37850 986 38086
rect 1222 37850 585502 38086
rect 585738 37850 586860 38086
rect -2936 37828 586860 37850
rect -1996 37826 -1396 37828
rect 804 37826 1404 37828
rect 585320 37826 585920 37828
rect -8576 31276 -7976 31278
rect 591900 31276 592500 31278
rect -8576 31254 592500 31276
rect -8576 31018 -8394 31254
rect -8158 31018 592082 31254
rect 592318 31018 592500 31254
rect -8576 30934 592500 31018
rect -8576 30698 -8394 30934
rect -8158 30698 592082 30934
rect 592318 30698 592500 30934
rect -8576 30676 592500 30698
rect -8576 30674 -7976 30676
rect 591900 30674 592500 30676
rect -6696 27676 -6096 27678
rect 590020 27676 590620 27678
rect -6696 27654 590620 27676
rect -6696 27418 -6514 27654
rect -6278 27418 590202 27654
rect 590438 27418 590620 27654
rect -6696 27334 590620 27418
rect -6696 27098 -6514 27334
rect -6278 27098 590202 27334
rect 590438 27098 590620 27334
rect -6696 27076 590620 27098
rect -6696 27074 -6096 27076
rect 590020 27074 590620 27076
rect -4816 24076 -4216 24078
rect 588140 24076 588740 24078
rect -4816 24054 588740 24076
rect -4816 23818 -4634 24054
rect -4398 23818 588322 24054
rect 588558 23818 588740 24054
rect -4816 23734 588740 23818
rect -4816 23498 -4634 23734
rect -4398 23498 588322 23734
rect 588558 23498 588740 23734
rect -4816 23476 588740 23498
rect -4816 23474 -4216 23476
rect 588140 23474 588740 23476
rect -2936 20428 -2336 20430
rect 586260 20428 586860 20430
rect -2936 20406 586860 20428
rect -2936 20170 -2754 20406
rect -2518 20170 586442 20406
rect 586678 20170 586860 20406
rect -2936 20086 586860 20170
rect -2936 19850 -2754 20086
rect -2518 19850 586442 20086
rect 586678 19850 586860 20086
rect -2936 19828 586860 19850
rect -2936 19826 -2336 19828
rect 586260 19826 586860 19828
rect -7636 13276 -7036 13278
rect 590960 13276 591560 13278
rect -8576 13254 592500 13276
rect -8576 13018 -7454 13254
rect -7218 13018 591142 13254
rect 591378 13018 592500 13254
rect -8576 12934 592500 13018
rect -8576 12698 -7454 12934
rect -7218 12698 591142 12934
rect 591378 12698 592500 12934
rect -8576 12676 592500 12698
rect -7636 12674 -7036 12676
rect 590960 12674 591560 12676
rect -5756 9676 -5156 9678
rect 589080 9676 589680 9678
rect -6696 9654 590620 9676
rect -6696 9418 -5574 9654
rect -5338 9418 589262 9654
rect 589498 9418 590620 9654
rect -6696 9334 590620 9418
rect -6696 9098 -5574 9334
rect -5338 9098 589262 9334
rect 589498 9098 590620 9334
rect -6696 9076 590620 9098
rect -5756 9074 -5156 9076
rect 589080 9074 589680 9076
rect -3876 6076 -3276 6078
rect 4404 6076 5004 6078
rect 580404 6076 581004 6078
rect 587200 6076 587800 6078
rect -4816 6054 588740 6076
rect -4816 5818 -3694 6054
rect -3458 5818 4586 6054
rect 4822 5818 580586 6054
rect 580822 5818 587382 6054
rect 587618 5818 588740 6054
rect -4816 5734 588740 5818
rect -4816 5498 -3694 5734
rect -3458 5498 4586 5734
rect 4822 5498 580586 5734
rect 580822 5498 587382 5734
rect 587618 5498 588740 5734
rect -4816 5476 588740 5498
rect -3876 5474 -3276 5476
rect 4404 5474 5004 5476
rect 580404 5474 581004 5476
rect 587200 5474 587800 5476
rect -1996 2428 -1396 2430
rect 804 2428 1404 2430
rect 36804 2428 37404 2430
rect 72804 2428 73404 2430
rect 108804 2428 109404 2430
rect 144804 2428 145404 2430
rect 180804 2428 181404 2430
rect 216804 2428 217404 2430
rect 252804 2428 253404 2430
rect 288804 2428 289404 2430
rect 324804 2428 325404 2430
rect 360804 2428 361404 2430
rect 396804 2428 397404 2430
rect 432804 2428 433404 2430
rect 468804 2428 469404 2430
rect 504804 2428 505404 2430
rect 540804 2428 541404 2430
rect 576804 2428 577404 2430
rect 585320 2428 585920 2430
rect -2936 2406 586860 2428
rect -2936 2170 -1814 2406
rect -1578 2170 986 2406
rect 1222 2170 36986 2406
rect 37222 2170 72986 2406
rect 73222 2170 108986 2406
rect 109222 2170 144986 2406
rect 145222 2170 180986 2406
rect 181222 2170 216986 2406
rect 217222 2170 252986 2406
rect 253222 2170 288986 2406
rect 289222 2170 324986 2406
rect 325222 2170 360986 2406
rect 361222 2170 396986 2406
rect 397222 2170 432986 2406
rect 433222 2170 468986 2406
rect 469222 2170 504986 2406
rect 505222 2170 540986 2406
rect 541222 2170 576986 2406
rect 577222 2170 585502 2406
rect 585738 2170 586860 2406
rect -2936 2086 586860 2170
rect -2936 1850 -1814 2086
rect -1578 1850 986 2086
rect 1222 1850 36986 2086
rect 37222 1850 72986 2086
rect 73222 1850 108986 2086
rect 109222 1850 144986 2086
rect 145222 1850 180986 2086
rect 181222 1850 216986 2086
rect 217222 1850 252986 2086
rect 253222 1850 288986 2086
rect 289222 1850 324986 2086
rect 325222 1850 360986 2086
rect 361222 1850 396986 2086
rect 397222 1850 432986 2086
rect 433222 1850 468986 2086
rect 469222 1850 504986 2086
rect 505222 1850 540986 2086
rect 541222 1850 576986 2086
rect 577222 1850 585502 2086
rect 585738 1850 586860 2086
rect -2936 1828 586860 1850
rect -1996 1826 -1396 1828
rect 804 1826 1404 1828
rect 36804 1826 37404 1828
rect 72804 1826 73404 1828
rect 108804 1826 109404 1828
rect 144804 1826 145404 1828
rect 180804 1826 181404 1828
rect 216804 1826 217404 1828
rect 252804 1826 253404 1828
rect 288804 1826 289404 1828
rect 324804 1826 325404 1828
rect 360804 1826 361404 1828
rect 396804 1826 397404 1828
rect 432804 1826 433404 1828
rect 468804 1826 469404 1828
rect 504804 1826 505404 1828
rect 540804 1826 541404 1828
rect 576804 1826 577404 1828
rect 585320 1826 585920 1828
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2936 -1264 -2336 -1262
rect 18804 -1264 19404 -1262
rect 54804 -1264 55404 -1262
rect 90804 -1264 91404 -1262
rect 126804 -1264 127404 -1262
rect 162804 -1264 163404 -1262
rect 198804 -1264 199404 -1262
rect 234804 -1264 235404 -1262
rect 270804 -1264 271404 -1262
rect 306804 -1264 307404 -1262
rect 342804 -1264 343404 -1262
rect 378804 -1264 379404 -1262
rect 414804 -1264 415404 -1262
rect 450804 -1264 451404 -1262
rect 486804 -1264 487404 -1262
rect 522804 -1264 523404 -1262
rect 558804 -1264 559404 -1262
rect 586260 -1264 586860 -1262
rect -2936 -1286 586860 -1264
rect -2936 -1522 -2754 -1286
rect -2518 -1522 18986 -1286
rect 19222 -1522 54986 -1286
rect 55222 -1522 90986 -1286
rect 91222 -1522 126986 -1286
rect 127222 -1522 162986 -1286
rect 163222 -1522 198986 -1286
rect 199222 -1522 234986 -1286
rect 235222 -1522 270986 -1286
rect 271222 -1522 306986 -1286
rect 307222 -1522 342986 -1286
rect 343222 -1522 378986 -1286
rect 379222 -1522 414986 -1286
rect 415222 -1522 450986 -1286
rect 451222 -1522 486986 -1286
rect 487222 -1522 522986 -1286
rect 523222 -1522 558986 -1286
rect 559222 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect -2936 -1606 586860 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 18986 -1606
rect 19222 -1842 54986 -1606
rect 55222 -1842 90986 -1606
rect 91222 -1842 126986 -1606
rect 127222 -1842 162986 -1606
rect 163222 -1842 198986 -1606
rect 199222 -1842 234986 -1606
rect 235222 -1842 270986 -1606
rect 271222 -1842 306986 -1606
rect 307222 -1842 342986 -1606
rect 343222 -1842 378986 -1606
rect 379222 -1842 414986 -1606
rect 415222 -1842 450986 -1606
rect 451222 -1842 486986 -1606
rect 487222 -1842 522986 -1606
rect 523222 -1842 558986 -1606
rect 559222 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect -2936 -1864 586860 -1842
rect -2936 -1866 -2336 -1864
rect 18804 -1866 19404 -1864
rect 54804 -1866 55404 -1864
rect 90804 -1866 91404 -1864
rect 126804 -1866 127404 -1864
rect 162804 -1866 163404 -1864
rect 198804 -1866 199404 -1864
rect 234804 -1866 235404 -1864
rect 270804 -1866 271404 -1864
rect 306804 -1866 307404 -1864
rect 342804 -1866 343404 -1864
rect 378804 -1866 379404 -1864
rect 414804 -1866 415404 -1864
rect 450804 -1866 451404 -1864
rect 486804 -1866 487404 -1864
rect 522804 -1866 523404 -1864
rect 558804 -1866 559404 -1864
rect 586260 -1866 586860 -1864
rect -3876 -2204 -3276 -2202
rect 4404 -2204 5004 -2202
rect 40404 -2204 41004 -2202
rect 76404 -2204 77004 -2202
rect 112404 -2204 113004 -2202
rect 148404 -2204 149004 -2202
rect 184404 -2204 185004 -2202
rect 220404 -2204 221004 -2202
rect 256404 -2204 257004 -2202
rect 292404 -2204 293004 -2202
rect 328404 -2204 329004 -2202
rect 364404 -2204 365004 -2202
rect 400404 -2204 401004 -2202
rect 436404 -2204 437004 -2202
rect 472404 -2204 473004 -2202
rect 508404 -2204 509004 -2202
rect 544404 -2204 545004 -2202
rect 580404 -2204 581004 -2202
rect 587200 -2204 587800 -2202
rect -3876 -2226 587800 -2204
rect -3876 -2462 -3694 -2226
rect -3458 -2462 4586 -2226
rect 4822 -2462 40586 -2226
rect 40822 -2462 76586 -2226
rect 76822 -2462 112586 -2226
rect 112822 -2462 148586 -2226
rect 148822 -2462 184586 -2226
rect 184822 -2462 220586 -2226
rect 220822 -2462 256586 -2226
rect 256822 -2462 292586 -2226
rect 292822 -2462 328586 -2226
rect 328822 -2462 364586 -2226
rect 364822 -2462 400586 -2226
rect 400822 -2462 436586 -2226
rect 436822 -2462 472586 -2226
rect 472822 -2462 508586 -2226
rect 508822 -2462 544586 -2226
rect 544822 -2462 580586 -2226
rect 580822 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect -3876 -2546 587800 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 4586 -2546
rect 4822 -2782 40586 -2546
rect 40822 -2782 76586 -2546
rect 76822 -2782 112586 -2546
rect 112822 -2782 148586 -2546
rect 148822 -2782 184586 -2546
rect 184822 -2782 220586 -2546
rect 220822 -2782 256586 -2546
rect 256822 -2782 292586 -2546
rect 292822 -2782 328586 -2546
rect 328822 -2782 364586 -2546
rect 364822 -2782 400586 -2546
rect 400822 -2782 436586 -2546
rect 436822 -2782 472586 -2546
rect 472822 -2782 508586 -2546
rect 508822 -2782 544586 -2546
rect 544822 -2782 580586 -2546
rect 580822 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect -3876 -2804 587800 -2782
rect -3876 -2806 -3276 -2804
rect 4404 -2806 5004 -2804
rect 40404 -2806 41004 -2804
rect 76404 -2806 77004 -2804
rect 112404 -2806 113004 -2804
rect 148404 -2806 149004 -2804
rect 184404 -2806 185004 -2804
rect 220404 -2806 221004 -2804
rect 256404 -2806 257004 -2804
rect 292404 -2806 293004 -2804
rect 328404 -2806 329004 -2804
rect 364404 -2806 365004 -2804
rect 400404 -2806 401004 -2804
rect 436404 -2806 437004 -2804
rect 472404 -2806 473004 -2804
rect 508404 -2806 509004 -2804
rect 544404 -2806 545004 -2804
rect 580404 -2806 581004 -2804
rect 587200 -2806 587800 -2804
rect -4816 -3144 -4216 -3142
rect 22404 -3144 23004 -3142
rect 58404 -3144 59004 -3142
rect 94404 -3144 95004 -3142
rect 130404 -3144 131004 -3142
rect 166404 -3144 167004 -3142
rect 202404 -3144 203004 -3142
rect 238404 -3144 239004 -3142
rect 274404 -3144 275004 -3142
rect 310404 -3144 311004 -3142
rect 346404 -3144 347004 -3142
rect 382404 -3144 383004 -3142
rect 418404 -3144 419004 -3142
rect 454404 -3144 455004 -3142
rect 490404 -3144 491004 -3142
rect 526404 -3144 527004 -3142
rect 562404 -3144 563004 -3142
rect 588140 -3144 588740 -3142
rect -4816 -3166 588740 -3144
rect -4816 -3402 -4634 -3166
rect -4398 -3402 22586 -3166
rect 22822 -3402 58586 -3166
rect 58822 -3402 94586 -3166
rect 94822 -3402 130586 -3166
rect 130822 -3402 166586 -3166
rect 166822 -3402 202586 -3166
rect 202822 -3402 238586 -3166
rect 238822 -3402 274586 -3166
rect 274822 -3402 310586 -3166
rect 310822 -3402 346586 -3166
rect 346822 -3402 382586 -3166
rect 382822 -3402 418586 -3166
rect 418822 -3402 454586 -3166
rect 454822 -3402 490586 -3166
rect 490822 -3402 526586 -3166
rect 526822 -3402 562586 -3166
rect 562822 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect -4816 -3486 588740 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 22586 -3486
rect 22822 -3722 58586 -3486
rect 58822 -3722 94586 -3486
rect 94822 -3722 130586 -3486
rect 130822 -3722 166586 -3486
rect 166822 -3722 202586 -3486
rect 202822 -3722 238586 -3486
rect 238822 -3722 274586 -3486
rect 274822 -3722 310586 -3486
rect 310822 -3722 346586 -3486
rect 346822 -3722 382586 -3486
rect 382822 -3722 418586 -3486
rect 418822 -3722 454586 -3486
rect 454822 -3722 490586 -3486
rect 490822 -3722 526586 -3486
rect 526822 -3722 562586 -3486
rect 562822 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect -4816 -3744 588740 -3722
rect -4816 -3746 -4216 -3744
rect 22404 -3746 23004 -3744
rect 58404 -3746 59004 -3744
rect 94404 -3746 95004 -3744
rect 130404 -3746 131004 -3744
rect 166404 -3746 167004 -3744
rect 202404 -3746 203004 -3744
rect 238404 -3746 239004 -3744
rect 274404 -3746 275004 -3744
rect 310404 -3746 311004 -3744
rect 346404 -3746 347004 -3744
rect 382404 -3746 383004 -3744
rect 418404 -3746 419004 -3744
rect 454404 -3746 455004 -3744
rect 490404 -3746 491004 -3744
rect 526404 -3746 527004 -3744
rect 562404 -3746 563004 -3744
rect 588140 -3746 588740 -3744
rect -5756 -4084 -5156 -4082
rect 8004 -4084 8604 -4082
rect 44004 -4084 44604 -4082
rect 80004 -4084 80604 -4082
rect 116004 -4084 116604 -4082
rect 152004 -4084 152604 -4082
rect 188004 -4084 188604 -4082
rect 224004 -4084 224604 -4082
rect 260004 -4084 260604 -4082
rect 296004 -4084 296604 -4082
rect 332004 -4084 332604 -4082
rect 368004 -4084 368604 -4082
rect 404004 -4084 404604 -4082
rect 440004 -4084 440604 -4082
rect 476004 -4084 476604 -4082
rect 512004 -4084 512604 -4082
rect 548004 -4084 548604 -4082
rect 589080 -4084 589680 -4082
rect -5756 -4106 589680 -4084
rect -5756 -4342 -5574 -4106
rect -5338 -4342 8186 -4106
rect 8422 -4342 44186 -4106
rect 44422 -4342 80186 -4106
rect 80422 -4342 116186 -4106
rect 116422 -4342 152186 -4106
rect 152422 -4342 188186 -4106
rect 188422 -4342 224186 -4106
rect 224422 -4342 260186 -4106
rect 260422 -4342 296186 -4106
rect 296422 -4342 332186 -4106
rect 332422 -4342 368186 -4106
rect 368422 -4342 404186 -4106
rect 404422 -4342 440186 -4106
rect 440422 -4342 476186 -4106
rect 476422 -4342 512186 -4106
rect 512422 -4342 548186 -4106
rect 548422 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect -5756 -4426 589680 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 8186 -4426
rect 8422 -4662 44186 -4426
rect 44422 -4662 80186 -4426
rect 80422 -4662 116186 -4426
rect 116422 -4662 152186 -4426
rect 152422 -4662 188186 -4426
rect 188422 -4662 224186 -4426
rect 224422 -4662 260186 -4426
rect 260422 -4662 296186 -4426
rect 296422 -4662 332186 -4426
rect 332422 -4662 368186 -4426
rect 368422 -4662 404186 -4426
rect 404422 -4662 440186 -4426
rect 440422 -4662 476186 -4426
rect 476422 -4662 512186 -4426
rect 512422 -4662 548186 -4426
rect 548422 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect -5756 -4684 589680 -4662
rect -5756 -4686 -5156 -4684
rect 8004 -4686 8604 -4684
rect 44004 -4686 44604 -4684
rect 80004 -4686 80604 -4684
rect 116004 -4686 116604 -4684
rect 152004 -4686 152604 -4684
rect 188004 -4686 188604 -4684
rect 224004 -4686 224604 -4684
rect 260004 -4686 260604 -4684
rect 296004 -4686 296604 -4684
rect 332004 -4686 332604 -4684
rect 368004 -4686 368604 -4684
rect 404004 -4686 404604 -4684
rect 440004 -4686 440604 -4684
rect 476004 -4686 476604 -4684
rect 512004 -4686 512604 -4684
rect 548004 -4686 548604 -4684
rect 589080 -4686 589680 -4684
rect -6696 -5024 -6096 -5022
rect 26004 -5024 26604 -5022
rect 62004 -5024 62604 -5022
rect 98004 -5024 98604 -5022
rect 134004 -5024 134604 -5022
rect 170004 -5024 170604 -5022
rect 206004 -5024 206604 -5022
rect 242004 -5024 242604 -5022
rect 278004 -5024 278604 -5022
rect 314004 -5024 314604 -5022
rect 350004 -5024 350604 -5022
rect 386004 -5024 386604 -5022
rect 422004 -5024 422604 -5022
rect 458004 -5024 458604 -5022
rect 494004 -5024 494604 -5022
rect 530004 -5024 530604 -5022
rect 566004 -5024 566604 -5022
rect 590020 -5024 590620 -5022
rect -6696 -5046 590620 -5024
rect -6696 -5282 -6514 -5046
rect -6278 -5282 26186 -5046
rect 26422 -5282 62186 -5046
rect 62422 -5282 98186 -5046
rect 98422 -5282 134186 -5046
rect 134422 -5282 170186 -5046
rect 170422 -5282 206186 -5046
rect 206422 -5282 242186 -5046
rect 242422 -5282 278186 -5046
rect 278422 -5282 314186 -5046
rect 314422 -5282 350186 -5046
rect 350422 -5282 386186 -5046
rect 386422 -5282 422186 -5046
rect 422422 -5282 458186 -5046
rect 458422 -5282 494186 -5046
rect 494422 -5282 530186 -5046
rect 530422 -5282 566186 -5046
rect 566422 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect -6696 -5366 590620 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 26186 -5366
rect 26422 -5602 62186 -5366
rect 62422 -5602 98186 -5366
rect 98422 -5602 134186 -5366
rect 134422 -5602 170186 -5366
rect 170422 -5602 206186 -5366
rect 206422 -5602 242186 -5366
rect 242422 -5602 278186 -5366
rect 278422 -5602 314186 -5366
rect 314422 -5602 350186 -5366
rect 350422 -5602 386186 -5366
rect 386422 -5602 422186 -5366
rect 422422 -5602 458186 -5366
rect 458422 -5602 494186 -5366
rect 494422 -5602 530186 -5366
rect 530422 -5602 566186 -5366
rect 566422 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect -6696 -5624 590620 -5602
rect -6696 -5626 -6096 -5624
rect 26004 -5626 26604 -5624
rect 62004 -5626 62604 -5624
rect 98004 -5626 98604 -5624
rect 134004 -5626 134604 -5624
rect 170004 -5626 170604 -5624
rect 206004 -5626 206604 -5624
rect 242004 -5626 242604 -5624
rect 278004 -5626 278604 -5624
rect 314004 -5626 314604 -5624
rect 350004 -5626 350604 -5624
rect 386004 -5626 386604 -5624
rect 422004 -5626 422604 -5624
rect 458004 -5626 458604 -5624
rect 494004 -5626 494604 -5624
rect 530004 -5626 530604 -5624
rect 566004 -5626 566604 -5624
rect 590020 -5626 590620 -5624
rect -7636 -5964 -7036 -5962
rect 11604 -5964 12204 -5962
rect 47604 -5964 48204 -5962
rect 83604 -5964 84204 -5962
rect 119604 -5964 120204 -5962
rect 155604 -5964 156204 -5962
rect 191604 -5964 192204 -5962
rect 227604 -5964 228204 -5962
rect 263604 -5964 264204 -5962
rect 299604 -5964 300204 -5962
rect 335604 -5964 336204 -5962
rect 371604 -5964 372204 -5962
rect 407604 -5964 408204 -5962
rect 443604 -5964 444204 -5962
rect 479604 -5964 480204 -5962
rect 515604 -5964 516204 -5962
rect 551604 -5964 552204 -5962
rect 590960 -5964 591560 -5962
rect -7636 -5986 591560 -5964
rect -7636 -6222 -7454 -5986
rect -7218 -6222 11786 -5986
rect 12022 -6222 47786 -5986
rect 48022 -6222 83786 -5986
rect 84022 -6222 119786 -5986
rect 120022 -6222 155786 -5986
rect 156022 -6222 191786 -5986
rect 192022 -6222 227786 -5986
rect 228022 -6222 263786 -5986
rect 264022 -6222 299786 -5986
rect 300022 -6222 335786 -5986
rect 336022 -6222 371786 -5986
rect 372022 -6222 407786 -5986
rect 408022 -6222 443786 -5986
rect 444022 -6222 479786 -5986
rect 480022 -6222 515786 -5986
rect 516022 -6222 551786 -5986
rect 552022 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect -7636 -6306 591560 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 11786 -6306
rect 12022 -6542 47786 -6306
rect 48022 -6542 83786 -6306
rect 84022 -6542 119786 -6306
rect 120022 -6542 155786 -6306
rect 156022 -6542 191786 -6306
rect 192022 -6542 227786 -6306
rect 228022 -6542 263786 -6306
rect 264022 -6542 299786 -6306
rect 300022 -6542 335786 -6306
rect 336022 -6542 371786 -6306
rect 372022 -6542 407786 -6306
rect 408022 -6542 443786 -6306
rect 444022 -6542 479786 -6306
rect 480022 -6542 515786 -6306
rect 516022 -6542 551786 -6306
rect 552022 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect -7636 -6564 591560 -6542
rect -7636 -6566 -7036 -6564
rect 11604 -6566 12204 -6564
rect 47604 -6566 48204 -6564
rect 83604 -6566 84204 -6564
rect 119604 -6566 120204 -6564
rect 155604 -6566 156204 -6564
rect 191604 -6566 192204 -6564
rect 227604 -6566 228204 -6564
rect 263604 -6566 264204 -6564
rect 299604 -6566 300204 -6564
rect 335604 -6566 336204 -6564
rect 371604 -6566 372204 -6564
rect 407604 -6566 408204 -6564
rect 443604 -6566 444204 -6564
rect 479604 -6566 480204 -6564
rect 515604 -6566 516204 -6564
rect 551604 -6566 552204 -6564
rect 590960 -6566 591560 -6564
rect -8576 -6904 -7976 -6902
rect 29604 -6904 30204 -6902
rect 65604 -6904 66204 -6902
rect 101604 -6904 102204 -6902
rect 137604 -6904 138204 -6902
rect 173604 -6904 174204 -6902
rect 209604 -6904 210204 -6902
rect 245604 -6904 246204 -6902
rect 281604 -6904 282204 -6902
rect 317604 -6904 318204 -6902
rect 353604 -6904 354204 -6902
rect 389604 -6904 390204 -6902
rect 425604 -6904 426204 -6902
rect 461604 -6904 462204 -6902
rect 497604 -6904 498204 -6902
rect 533604 -6904 534204 -6902
rect 569604 -6904 570204 -6902
rect 591900 -6904 592500 -6902
rect -8576 -6926 592500 -6904
rect -8576 -7162 -8394 -6926
rect -8158 -7162 29786 -6926
rect 30022 -7162 65786 -6926
rect 66022 -7162 101786 -6926
rect 102022 -7162 137786 -6926
rect 138022 -7162 173786 -6926
rect 174022 -7162 209786 -6926
rect 210022 -7162 245786 -6926
rect 246022 -7162 281786 -6926
rect 282022 -7162 317786 -6926
rect 318022 -7162 353786 -6926
rect 354022 -7162 389786 -6926
rect 390022 -7162 425786 -6926
rect 426022 -7162 461786 -6926
rect 462022 -7162 497786 -6926
rect 498022 -7162 533786 -6926
rect 534022 -7162 569786 -6926
rect 570022 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect -8576 -7246 592500 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 29786 -7246
rect 30022 -7482 65786 -7246
rect 66022 -7482 101786 -7246
rect 102022 -7482 137786 -7246
rect 138022 -7482 173786 -7246
rect 174022 -7482 209786 -7246
rect 210022 -7482 245786 -7246
rect 246022 -7482 281786 -7246
rect 282022 -7482 317786 -7246
rect 318022 -7482 353786 -7246
rect 354022 -7482 389786 -7246
rect 390022 -7482 425786 -7246
rect 426022 -7482 461786 -7246
rect 462022 -7482 497786 -7246
rect 498022 -7482 533786 -7246
rect 534022 -7482 569786 -7246
rect 570022 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect -8576 -7504 592500 -7482
rect -8576 -7506 -7976 -7504
rect 29604 -7506 30204 -7504
rect 65604 -7506 66204 -7504
rect 101604 -7506 102204 -7504
rect 137604 -7506 138204 -7504
rect 173604 -7506 174204 -7504
rect 209604 -7506 210204 -7504
rect 245604 -7506 246204 -7504
rect 281604 -7506 282204 -7504
rect 317604 -7506 318204 -7504
rect 353604 -7506 354204 -7504
rect 389604 -7506 390204 -7504
rect 425604 -7506 426204 -7504
rect 461604 -7506 462204 -7504
rect 497604 -7506 498204 -7504
rect 533604 -7506 534204 -7504
rect 569604 -7506 570204 -7504
rect 591900 -7506 592500 -7504
use user_proj_example  mprj
timestamp 1608616637
transform 1 0 8000 0 1 8000
box 0 0 568000 688000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew signal bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew signal bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew signal bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew signal bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew signal input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew signal input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew signal input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew signal input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew signal input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew signal input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew signal input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew signal input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew signal input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew signal input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew signal input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew signal input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew signal input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew signal input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew signal input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew signal input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew signal input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew signal input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew signal input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew signal input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew signal input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew signal input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew signal input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew signal input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew signal input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew signal input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew signal input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew signal input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew signal input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew signal tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew signal tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew signal tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew signal tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew signal tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew signal tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew signal tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew signal tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew signal tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew signal tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew signal tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew signal tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew signal tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew signal tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew signal tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew signal tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew signal tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew signal tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew signal tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew signal tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew signal tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew signal tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew signal tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew signal tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew signal tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew signal tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew signal tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew signal tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew signal tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew signal tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew signal tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew signal tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew signal tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew signal tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew signal tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew signal tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew signal tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew signal tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew signal tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew signal tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew signal tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew signal tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew signal tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew signal tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew signal tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew signal tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew signal tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew signal tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew signal tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew signal tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew signal tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew signal tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew signal tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew signal tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew signal tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew signal tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew signal tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew signal tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew signal input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew signal input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew signal input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew signal input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew signal input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew signal input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew signal input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew signal input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew signal input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew signal input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew signal input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew signal input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew signal input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew signal input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew signal input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew signal input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew signal input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew signal input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew signal input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew signal input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew signal input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew signal input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew signal input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew signal input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew signal input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew signal input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew signal input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew signal input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew signal input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew signal input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew signal input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew signal input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew signal input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew signal input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew signal input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew signal input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew signal input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew signal input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew signal input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew signal input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew signal input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew signal input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew signal input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew signal input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew signal input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew signal input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew signal input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew signal input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew signal input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew signal input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew signal input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew signal input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew signal input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew signal input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew signal input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew signal input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew signal input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew signal input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew signal input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew signal input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew signal input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew signal input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew signal input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew signal input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew signal input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew signal input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew signal input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew signal input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew signal input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew signal input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew signal input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew signal input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew signal input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew signal input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew signal input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew signal input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew signal input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew signal input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew signal input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew signal input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew signal input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew signal input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew signal input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew signal input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew signal input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew signal input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew signal input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew signal input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew signal input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew signal input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew signal input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew signal input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew signal input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew signal input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew signal input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew signal input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew signal input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew signal input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew signal input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew signal input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew signal input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew signal input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew signal input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew signal input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew signal input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew signal input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew signal input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew signal input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew signal input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew signal input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew signal input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew signal input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew signal input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew signal input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew signal input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew signal input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew signal input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew signal input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew signal input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew signal input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew signal input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew signal input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew signal tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew signal tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew signal tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew signal tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew signal tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew signal tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew signal tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew signal tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew signal tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew signal tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew signal tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew signal tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew signal tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew signal tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew signal tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew signal tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew signal tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew signal tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew signal tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew signal tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew signal tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew signal tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew signal tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew signal tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew signal tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew signal tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew signal tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew signal tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew signal tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew signal tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew signal tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew signal tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew signal tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew signal tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew signal tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew signal tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew signal tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew signal tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew signal tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew signal tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew signal tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew signal tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew signal tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew signal tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew signal tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew signal tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew signal tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew signal tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew signal tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew signal tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew signal tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew signal tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew signal tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew signal tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew signal tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew signal tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew signal tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew signal tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew signal tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew signal tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew signal tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew signal tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew signal tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew signal tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew signal tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew signal tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew signal tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew signal tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew signal tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew signal tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew signal tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew signal tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew signal tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew signal tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew signal tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew signal tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew signal tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew signal tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew signal tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew signal tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew signal tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew signal tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew signal tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew signal tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew signal tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew signal tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew signal tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew signal tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew signal tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew signal tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew signal tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew signal tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew signal tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew signal tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew signal tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew signal tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew signal tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew signal tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew signal tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew signal tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew signal tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew signal tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew signal tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew signal tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew signal tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew signal tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew signal tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew signal tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew signal tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew signal tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew signal tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew signal tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew signal tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew signal tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew signal tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew signal tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew signal tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew signal tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew signal tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew signal tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew signal tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew signal tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew signal tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew signal tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew signal tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew signal tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew signal tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew signal input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew signal input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew signal input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew signal input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew signal input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew signal input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew signal input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew signal input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew signal input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew signal input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew signal input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew signal input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew signal input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew signal input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew signal input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew signal input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew signal input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew signal input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew signal input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew signal input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew signal input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew signal input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew signal input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew signal input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew signal input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew signal input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew signal input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew signal input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew signal input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew signal input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew signal input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew signal input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew signal input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew signal input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew signal input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew signal input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew signal input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew signal input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew signal input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew signal input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew signal input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew signal input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew signal input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew signal input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew signal input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew signal input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew signal input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew signal input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew signal input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew signal input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew signal input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew signal input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew signal input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew signal input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew signal input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew signal input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew signal input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew signal input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew signal input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew signal input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew signal input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew signal input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew signal input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew signal input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew signal input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew signal input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew signal input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew signal input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew signal input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew signal input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew signal input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew signal input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew signal input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew signal input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew signal input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew signal input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew signal input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew signal input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew signal input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew signal input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew signal input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew signal input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew signal input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew signal input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew signal input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew signal input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew signal input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew signal input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew signal input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew signal input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew signal input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew signal input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew signal input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew signal input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew signal input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew signal input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew signal input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew signal input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew signal input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew signal input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew signal input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew signal input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew signal input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew signal input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew signal input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew signal input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew signal input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew signal input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew signal input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew signal input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew signal input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew signal input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew signal input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew signal input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew signal input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew signal input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew signal input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew signal input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew signal input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew signal input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew signal input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew signal input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew signal input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew signal input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew signal input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew signal input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew signal input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew signal input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew signal input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew signal input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew signal input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew signal input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew signal input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew signal input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew signal input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew signal input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew signal input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew signal input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew signal input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew signal input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew signal input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew signal input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew signal input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew signal input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew signal input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew signal input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew signal input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew signal input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew signal input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew signal input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew signal input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew signal input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew signal input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew signal input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew signal input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew signal input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew signal input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew signal input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew signal input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew signal input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew signal input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew signal input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew signal input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew signal input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew signal input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew signal input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew signal input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew signal input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew signal input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew signal input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew signal input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew signal input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew signal input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew signal input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew signal input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew signal input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew signal input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew signal input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew signal input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew signal input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew signal input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew signal input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew signal input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew signal input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew signal input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew signal input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew signal input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew signal input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew signal tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew signal tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew signal tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew signal tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew signal tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew signal tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew signal tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew signal tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew signal tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew signal tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew signal tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew signal tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew signal tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew signal tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew signal tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew signal tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew signal tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew signal tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew signal tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew signal tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew signal tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew signal tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew signal tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew signal tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew signal tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew signal tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew signal tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew signal tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew signal tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew signal tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew signal tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew signal tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew signal input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew signal input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew signal input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew signal input
rlabel metal4 s 576804 697952 577404 705800 6 vccd1
port 636 nsew power bidirectional
rlabel metal4 s 540804 697952 541404 705800 6 vccd1
port 637 nsew power bidirectional
rlabel metal4 s 504804 697952 505404 705800 6 vccd1
port 638 nsew power bidirectional
rlabel metal4 s 468804 697952 469404 705800 6 vccd1
port 639 nsew power bidirectional
rlabel metal4 s 432804 697952 433404 705800 6 vccd1
port 640 nsew power bidirectional
rlabel metal4 s 396804 697952 397404 705800 6 vccd1
port 641 nsew power bidirectional
rlabel metal4 s 360804 697952 361404 705800 6 vccd1
port 642 nsew power bidirectional
rlabel metal4 s 324804 697952 325404 705800 6 vccd1
port 643 nsew power bidirectional
rlabel metal4 s 288804 697952 289404 705800 6 vccd1
port 644 nsew power bidirectional
rlabel metal4 s 252804 697952 253404 705800 6 vccd1
port 645 nsew power bidirectional
rlabel metal4 s 216804 697952 217404 705800 6 vccd1
port 646 nsew power bidirectional
rlabel metal4 s 180804 697952 181404 705800 6 vccd1
port 647 nsew power bidirectional
rlabel metal4 s 144804 697952 145404 705800 6 vccd1
port 648 nsew power bidirectional
rlabel metal4 s 108804 697952 109404 705800 6 vccd1
port 649 nsew power bidirectional
rlabel metal4 s 72804 697952 73404 705800 6 vccd1
port 650 nsew power bidirectional
rlabel metal4 s 36804 697952 37404 705800 6 vccd1
port 651 nsew power bidirectional
rlabel metal4 s 804 -1864 1404 705800 6 vccd1
port 652 nsew power bidirectional
rlabel metal4 s 585320 -924 585920 704860 6 vccd1
port 653 nsew power bidirectional
rlabel metal4 s -1996 -924 -1396 704860 4 vccd1
port 654 nsew power bidirectional
rlabel metal4 s 576804 -1864 577404 6048 6 vccd1
port 655 nsew power bidirectional
rlabel metal4 s 540804 -1864 541404 6048 6 vccd1
port 656 nsew power bidirectional
rlabel metal4 s 504804 -1864 505404 6048 6 vccd1
port 657 nsew power bidirectional
rlabel metal4 s 468804 -1864 469404 6048 6 vccd1
port 658 nsew power bidirectional
rlabel metal4 s 432804 -1864 433404 6048 6 vccd1
port 659 nsew power bidirectional
rlabel metal4 s 396804 -1864 397404 6048 6 vccd1
port 660 nsew power bidirectional
rlabel metal4 s 360804 -1864 361404 6048 6 vccd1
port 661 nsew power bidirectional
rlabel metal4 s 324804 -1864 325404 6048 6 vccd1
port 662 nsew power bidirectional
rlabel metal4 s 288804 -1864 289404 6048 6 vccd1
port 663 nsew power bidirectional
rlabel metal4 s 252804 -1864 253404 6048 6 vccd1
port 664 nsew power bidirectional
rlabel metal4 s 216804 -1864 217404 6048 6 vccd1
port 665 nsew power bidirectional
rlabel metal4 s 180804 -1864 181404 6048 6 vccd1
port 666 nsew power bidirectional
rlabel metal4 s 144804 -1864 145404 6048 6 vccd1
port 667 nsew power bidirectional
rlabel metal4 s 108804 -1864 109404 6048 6 vccd1
port 668 nsew power bidirectional
rlabel metal4 s 72804 -1864 73404 6048 6 vccd1
port 669 nsew power bidirectional
rlabel metal4 s 36804 -1864 37404 6048 6 vccd1
port 670 nsew power bidirectional
rlabel metal5 s -1996 704260 585920 704860 6 vccd1
port 671 nsew power bidirectional
rlabel metal5 s -2936 685828 586860 686428 6 vccd1
port 672 nsew power bidirectional
rlabel metal5 s -2936 649828 586860 650428 6 vccd1
port 673 nsew power bidirectional
rlabel metal5 s -2936 613828 586860 614428 6 vccd1
port 674 nsew power bidirectional
rlabel metal5 s -2936 577828 586860 578428 6 vccd1
port 675 nsew power bidirectional
rlabel metal5 s -2936 541828 586860 542428 6 vccd1
port 676 nsew power bidirectional
rlabel metal5 s -2936 505828 586860 506428 6 vccd1
port 677 nsew power bidirectional
rlabel metal5 s -2936 469828 586860 470428 6 vccd1
port 678 nsew power bidirectional
rlabel metal5 s -2936 433828 586860 434428 6 vccd1
port 679 nsew power bidirectional
rlabel metal5 s -2936 397828 586860 398428 6 vccd1
port 680 nsew power bidirectional
rlabel metal5 s -2936 361828 586860 362428 6 vccd1
port 681 nsew power bidirectional
rlabel metal5 s -2936 325828 586860 326428 6 vccd1
port 682 nsew power bidirectional
rlabel metal5 s -2936 289828 586860 290428 6 vccd1
port 683 nsew power bidirectional
rlabel metal5 s -2936 253828 586860 254428 6 vccd1
port 684 nsew power bidirectional
rlabel metal5 s -2936 217828 586860 218428 6 vccd1
port 685 nsew power bidirectional
rlabel metal5 s -2936 181828 586860 182428 6 vccd1
port 686 nsew power bidirectional
rlabel metal5 s -2936 145828 586860 146428 6 vccd1
port 687 nsew power bidirectional
rlabel metal5 s -2936 109828 586860 110428 6 vccd1
port 688 nsew power bidirectional
rlabel metal5 s -2936 73828 586860 74428 6 vccd1
port 689 nsew power bidirectional
rlabel metal5 s -2936 37828 586860 38428 6 vccd1
port 690 nsew power bidirectional
rlabel metal5 s -2936 1828 586860 2428 6 vccd1
port 691 nsew power bidirectional
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 692 nsew power bidirectional
rlabel metal4 s 586260 -1864 586860 705800 6 vssd1
port 693 nsew ground bidirectional
rlabel metal4 s 558804 697952 559404 705800 6 vssd1
port 694 nsew ground bidirectional
rlabel metal4 s 522804 697952 523404 705800 6 vssd1
port 695 nsew ground bidirectional
rlabel metal4 s 486804 697952 487404 705800 6 vssd1
port 696 nsew ground bidirectional
rlabel metal4 s 450804 697952 451404 705800 6 vssd1
port 697 nsew ground bidirectional
rlabel metal4 s 414804 697952 415404 705800 6 vssd1
port 698 nsew ground bidirectional
rlabel metal4 s 378804 697952 379404 705800 6 vssd1
port 699 nsew ground bidirectional
rlabel metal4 s 342804 697952 343404 705800 6 vssd1
port 700 nsew ground bidirectional
rlabel metal4 s 306804 697952 307404 705800 6 vssd1
port 701 nsew ground bidirectional
rlabel metal4 s 270804 697952 271404 705800 6 vssd1
port 702 nsew ground bidirectional
rlabel metal4 s 234804 697952 235404 705800 6 vssd1
port 703 nsew ground bidirectional
rlabel metal4 s 198804 697952 199404 705800 6 vssd1
port 704 nsew ground bidirectional
rlabel metal4 s 162804 697952 163404 705800 6 vssd1
port 705 nsew ground bidirectional
rlabel metal4 s 126804 697952 127404 705800 6 vssd1
port 706 nsew ground bidirectional
rlabel metal4 s 90804 697952 91404 705800 6 vssd1
port 707 nsew ground bidirectional
rlabel metal4 s 54804 697952 55404 705800 6 vssd1
port 708 nsew ground bidirectional
rlabel metal4 s 18804 697952 19404 705800 6 vssd1
port 709 nsew ground bidirectional
rlabel metal4 s -2936 -1864 -2336 705800 4 vssd1
port 710 nsew ground bidirectional
rlabel metal4 s 558804 -1864 559404 6048 6 vssd1
port 711 nsew ground bidirectional
rlabel metal4 s 522804 -1864 523404 6048 6 vssd1
port 712 nsew ground bidirectional
rlabel metal4 s 486804 -1864 487404 6048 6 vssd1
port 713 nsew ground bidirectional
rlabel metal4 s 450804 -1864 451404 6048 6 vssd1
port 714 nsew ground bidirectional
rlabel metal4 s 414804 -1864 415404 6048 6 vssd1
port 715 nsew ground bidirectional
rlabel metal4 s 378804 -1864 379404 6048 6 vssd1
port 716 nsew ground bidirectional
rlabel metal4 s 342804 -1864 343404 6048 6 vssd1
port 717 nsew ground bidirectional
rlabel metal4 s 306804 -1864 307404 6048 6 vssd1
port 718 nsew ground bidirectional
rlabel metal4 s 270804 -1864 271404 6048 6 vssd1
port 719 nsew ground bidirectional
rlabel metal4 s 234804 -1864 235404 6048 6 vssd1
port 720 nsew ground bidirectional
rlabel metal4 s 198804 -1864 199404 6048 6 vssd1
port 721 nsew ground bidirectional
rlabel metal4 s 162804 -1864 163404 6048 6 vssd1
port 722 nsew ground bidirectional
rlabel metal4 s 126804 -1864 127404 6048 6 vssd1
port 723 nsew ground bidirectional
rlabel metal4 s 90804 -1864 91404 6048 6 vssd1
port 724 nsew ground bidirectional
rlabel metal4 s 54804 -1864 55404 6048 6 vssd1
port 725 nsew ground bidirectional
rlabel metal4 s 18804 -1864 19404 6048 6 vssd1
port 726 nsew ground bidirectional
rlabel metal5 s -2936 705200 586860 705800 6 vssd1
port 727 nsew ground bidirectional
rlabel metal5 s -2936 667828 586860 668428 6 vssd1
port 728 nsew ground bidirectional
rlabel metal5 s -2936 631828 586860 632428 6 vssd1
port 729 nsew ground bidirectional
rlabel metal5 s -2936 595828 586860 596428 6 vssd1
port 730 nsew ground bidirectional
rlabel metal5 s -2936 559828 586860 560428 6 vssd1
port 731 nsew ground bidirectional
rlabel metal5 s -2936 523828 586860 524428 6 vssd1
port 732 nsew ground bidirectional
rlabel metal5 s -2936 487828 586860 488428 6 vssd1
port 733 nsew ground bidirectional
rlabel metal5 s -2936 451828 586860 452428 6 vssd1
port 734 nsew ground bidirectional
rlabel metal5 s -2936 415828 586860 416428 6 vssd1
port 735 nsew ground bidirectional
rlabel metal5 s -2936 379828 586860 380428 6 vssd1
port 736 nsew ground bidirectional
rlabel metal5 s -2936 343828 586860 344428 6 vssd1
port 737 nsew ground bidirectional
rlabel metal5 s -2936 307828 586860 308428 6 vssd1
port 738 nsew ground bidirectional
rlabel metal5 s -2936 271828 586860 272428 6 vssd1
port 739 nsew ground bidirectional
rlabel metal5 s -2936 235828 586860 236428 6 vssd1
port 740 nsew ground bidirectional
rlabel metal5 s -2936 199828 586860 200428 6 vssd1
port 741 nsew ground bidirectional
rlabel metal5 s -2936 163828 586860 164428 6 vssd1
port 742 nsew ground bidirectional
rlabel metal5 s -2936 127828 586860 128428 6 vssd1
port 743 nsew ground bidirectional
rlabel metal5 s -2936 91828 586860 92428 6 vssd1
port 744 nsew ground bidirectional
rlabel metal5 s -2936 55828 586860 56428 6 vssd1
port 745 nsew ground bidirectional
rlabel metal5 s -2936 19828 586860 20428 6 vssd1
port 746 nsew ground bidirectional
rlabel metal5 s -2936 -1864 586860 -1264 8 vssd1
port 747 nsew ground bidirectional
rlabel metal4 s 580404 -3744 581004 707680 6 vccd2
port 748 nsew power bidirectional
rlabel metal4 s 544404 698000 545004 707680 6 vccd2
port 749 nsew power bidirectional
rlabel metal4 s 508404 698000 509004 707680 6 vccd2
port 750 nsew power bidirectional
rlabel metal4 s 472404 698000 473004 707680 6 vccd2
port 751 nsew power bidirectional
rlabel metal4 s 436404 698000 437004 707680 6 vccd2
port 752 nsew power bidirectional
rlabel metal4 s 400404 698000 401004 707680 6 vccd2
port 753 nsew power bidirectional
rlabel metal4 s 364404 698000 365004 707680 6 vccd2
port 754 nsew power bidirectional
rlabel metal4 s 328404 698000 329004 707680 6 vccd2
port 755 nsew power bidirectional
rlabel metal4 s 292404 698000 293004 707680 6 vccd2
port 756 nsew power bidirectional
rlabel metal4 s 256404 698000 257004 707680 6 vccd2
port 757 nsew power bidirectional
rlabel metal4 s 220404 698000 221004 707680 6 vccd2
port 758 nsew power bidirectional
rlabel metal4 s 184404 698000 185004 707680 6 vccd2
port 759 nsew power bidirectional
rlabel metal4 s 148404 698000 149004 707680 6 vccd2
port 760 nsew power bidirectional
rlabel metal4 s 112404 698000 113004 707680 6 vccd2
port 761 nsew power bidirectional
rlabel metal4 s 76404 698000 77004 707680 6 vccd2
port 762 nsew power bidirectional
rlabel metal4 s 40404 698000 41004 707680 6 vccd2
port 763 nsew power bidirectional
rlabel metal4 s 4404 -3744 5004 707680 6 vccd2
port 764 nsew power bidirectional
rlabel metal4 s 587200 -2804 587800 706740 6 vccd2
port 765 nsew power bidirectional
rlabel metal4 s -3876 -2804 -3276 706740 4 vccd2
port 766 nsew power bidirectional
rlabel metal4 s 544404 -3744 545004 6000 6 vccd2
port 767 nsew power bidirectional
rlabel metal4 s 508404 -3744 509004 6000 6 vccd2
port 768 nsew power bidirectional
rlabel metal4 s 472404 -3744 473004 6000 6 vccd2
port 769 nsew power bidirectional
rlabel metal4 s 436404 -3744 437004 6000 6 vccd2
port 770 nsew power bidirectional
rlabel metal4 s 400404 -3744 401004 6000 6 vccd2
port 771 nsew power bidirectional
rlabel metal4 s 364404 -3744 365004 6000 6 vccd2
port 772 nsew power bidirectional
rlabel metal4 s 328404 -3744 329004 6000 6 vccd2
port 773 nsew power bidirectional
rlabel metal4 s 292404 -3744 293004 6000 6 vccd2
port 774 nsew power bidirectional
rlabel metal4 s 256404 -3744 257004 6000 6 vccd2
port 775 nsew power bidirectional
rlabel metal4 s 220404 -3744 221004 6000 6 vccd2
port 776 nsew power bidirectional
rlabel metal4 s 184404 -3744 185004 6000 6 vccd2
port 777 nsew power bidirectional
rlabel metal4 s 148404 -3744 149004 6000 6 vccd2
port 778 nsew power bidirectional
rlabel metal4 s 112404 -3744 113004 6000 6 vccd2
port 779 nsew power bidirectional
rlabel metal4 s 76404 -3744 77004 6000 6 vccd2
port 780 nsew power bidirectional
rlabel metal4 s 40404 -3744 41004 6000 6 vccd2
port 781 nsew power bidirectional
rlabel metal5 s -3876 706140 587800 706740 6 vccd2
port 782 nsew power bidirectional
rlabel metal5 s -4816 689476 588740 690076 6 vccd2
port 783 nsew power bidirectional
rlabel metal5 s -4816 653476 588740 654076 6 vccd2
port 784 nsew power bidirectional
rlabel metal5 s -4816 617476 588740 618076 6 vccd2
port 785 nsew power bidirectional
rlabel metal5 s -4816 581476 588740 582076 6 vccd2
port 786 nsew power bidirectional
rlabel metal5 s -4816 545476 588740 546076 6 vccd2
port 787 nsew power bidirectional
rlabel metal5 s -4816 509476 588740 510076 6 vccd2
port 788 nsew power bidirectional
rlabel metal5 s -4816 473476 588740 474076 6 vccd2
port 789 nsew power bidirectional
rlabel metal5 s -4816 437476 588740 438076 6 vccd2
port 790 nsew power bidirectional
rlabel metal5 s -4816 401476 588740 402076 6 vccd2
port 791 nsew power bidirectional
rlabel metal5 s -4816 365476 588740 366076 6 vccd2
port 792 nsew power bidirectional
rlabel metal5 s -4816 329476 588740 330076 6 vccd2
port 793 nsew power bidirectional
rlabel metal5 s -4816 293476 588740 294076 6 vccd2
port 794 nsew power bidirectional
rlabel metal5 s -4816 257476 588740 258076 6 vccd2
port 795 nsew power bidirectional
rlabel metal5 s -4816 221476 588740 222076 6 vccd2
port 796 nsew power bidirectional
rlabel metal5 s -4816 185476 588740 186076 6 vccd2
port 797 nsew power bidirectional
rlabel metal5 s -4816 149476 588740 150076 6 vccd2
port 798 nsew power bidirectional
rlabel metal5 s -4816 113476 588740 114076 6 vccd2
port 799 nsew power bidirectional
rlabel metal5 s -4816 77476 588740 78076 6 vccd2
port 800 nsew power bidirectional
rlabel metal5 s -4816 41476 588740 42076 6 vccd2
port 801 nsew power bidirectional
rlabel metal5 s -4816 5476 588740 6076 6 vccd2
port 802 nsew power bidirectional
rlabel metal5 s -3876 -2804 587800 -2204 8 vccd2
port 803 nsew power bidirectional
rlabel metal4 s 588140 -3744 588740 707680 6 vssd2
port 804 nsew ground bidirectional
rlabel metal4 s 562404 698000 563004 707680 6 vssd2
port 805 nsew ground bidirectional
rlabel metal4 s 526404 698000 527004 707680 6 vssd2
port 806 nsew ground bidirectional
rlabel metal4 s 490404 698000 491004 707680 6 vssd2
port 807 nsew ground bidirectional
rlabel metal4 s 454404 698000 455004 707680 6 vssd2
port 808 nsew ground bidirectional
rlabel metal4 s 418404 698000 419004 707680 6 vssd2
port 809 nsew ground bidirectional
rlabel metal4 s 382404 698000 383004 707680 6 vssd2
port 810 nsew ground bidirectional
rlabel metal4 s 346404 698000 347004 707680 6 vssd2
port 811 nsew ground bidirectional
rlabel metal4 s 310404 698000 311004 707680 6 vssd2
port 812 nsew ground bidirectional
rlabel metal4 s 274404 698000 275004 707680 6 vssd2
port 813 nsew ground bidirectional
rlabel metal4 s 238404 698000 239004 707680 6 vssd2
port 814 nsew ground bidirectional
rlabel metal4 s 202404 698000 203004 707680 6 vssd2
port 815 nsew ground bidirectional
rlabel metal4 s 166404 698000 167004 707680 6 vssd2
port 816 nsew ground bidirectional
rlabel metal4 s 130404 698000 131004 707680 6 vssd2
port 817 nsew ground bidirectional
rlabel metal4 s 94404 698000 95004 707680 6 vssd2
port 818 nsew ground bidirectional
rlabel metal4 s 58404 698000 59004 707680 6 vssd2
port 819 nsew ground bidirectional
rlabel metal4 s 22404 698000 23004 707680 6 vssd2
port 820 nsew ground bidirectional
rlabel metal4 s -4816 -3744 -4216 707680 4 vssd2
port 821 nsew ground bidirectional
rlabel metal4 s 562404 -3744 563004 6000 6 vssd2
port 822 nsew ground bidirectional
rlabel metal4 s 526404 -3744 527004 6000 6 vssd2
port 823 nsew ground bidirectional
rlabel metal4 s 490404 -3744 491004 6000 6 vssd2
port 824 nsew ground bidirectional
rlabel metal4 s 454404 -3744 455004 6000 6 vssd2
port 825 nsew ground bidirectional
rlabel metal4 s 418404 -3744 419004 6000 6 vssd2
port 826 nsew ground bidirectional
rlabel metal4 s 382404 -3744 383004 6000 6 vssd2
port 827 nsew ground bidirectional
rlabel metal4 s 346404 -3744 347004 6000 6 vssd2
port 828 nsew ground bidirectional
rlabel metal4 s 310404 -3744 311004 6000 6 vssd2
port 829 nsew ground bidirectional
rlabel metal4 s 274404 -3744 275004 6000 6 vssd2
port 830 nsew ground bidirectional
rlabel metal4 s 238404 -3744 239004 6000 6 vssd2
port 831 nsew ground bidirectional
rlabel metal4 s 202404 -3744 203004 6000 6 vssd2
port 832 nsew ground bidirectional
rlabel metal4 s 166404 -3744 167004 6000 6 vssd2
port 833 nsew ground bidirectional
rlabel metal4 s 130404 -3744 131004 6000 6 vssd2
port 834 nsew ground bidirectional
rlabel metal4 s 94404 -3744 95004 6000 6 vssd2
port 835 nsew ground bidirectional
rlabel metal4 s 58404 -3744 59004 6000 6 vssd2
port 836 nsew ground bidirectional
rlabel metal4 s 22404 -3744 23004 6000 6 vssd2
port 837 nsew ground bidirectional
rlabel metal5 s -4816 707080 588740 707680 6 vssd2
port 838 nsew ground bidirectional
rlabel metal5 s -4816 671476 588740 672076 6 vssd2
port 839 nsew ground bidirectional
rlabel metal5 s -4816 635476 588740 636076 6 vssd2
port 840 nsew ground bidirectional
rlabel metal5 s -4816 599476 588740 600076 6 vssd2
port 841 nsew ground bidirectional
rlabel metal5 s -4816 563476 588740 564076 6 vssd2
port 842 nsew ground bidirectional
rlabel metal5 s -4816 527476 588740 528076 6 vssd2
port 843 nsew ground bidirectional
rlabel metal5 s -4816 491476 588740 492076 6 vssd2
port 844 nsew ground bidirectional
rlabel metal5 s -4816 455476 588740 456076 6 vssd2
port 845 nsew ground bidirectional
rlabel metal5 s -4816 419476 588740 420076 6 vssd2
port 846 nsew ground bidirectional
rlabel metal5 s -4816 383476 588740 384076 6 vssd2
port 847 nsew ground bidirectional
rlabel metal5 s -4816 347476 588740 348076 6 vssd2
port 848 nsew ground bidirectional
rlabel metal5 s -4816 311476 588740 312076 6 vssd2
port 849 nsew ground bidirectional
rlabel metal5 s -4816 275476 588740 276076 6 vssd2
port 850 nsew ground bidirectional
rlabel metal5 s -4816 239476 588740 240076 6 vssd2
port 851 nsew ground bidirectional
rlabel metal5 s -4816 203476 588740 204076 6 vssd2
port 852 nsew ground bidirectional
rlabel metal5 s -4816 167476 588740 168076 6 vssd2
port 853 nsew ground bidirectional
rlabel metal5 s -4816 131476 588740 132076 6 vssd2
port 854 nsew ground bidirectional
rlabel metal5 s -4816 95476 588740 96076 6 vssd2
port 855 nsew ground bidirectional
rlabel metal5 s -4816 59476 588740 60076 6 vssd2
port 856 nsew ground bidirectional
rlabel metal5 s -4816 23476 588740 24076 6 vssd2
port 857 nsew ground bidirectional
rlabel metal5 s -4816 -3744 588740 -3144 8 vssd2
port 858 nsew ground bidirectional
rlabel metal4 s 548004 698000 548604 709560 6 vdda1
port 859 nsew power bidirectional
rlabel metal4 s 512004 698000 512604 709560 6 vdda1
port 860 nsew power bidirectional
rlabel metal4 s 476004 698000 476604 709560 6 vdda1
port 861 nsew power bidirectional
rlabel metal4 s 440004 698000 440604 709560 6 vdda1
port 862 nsew power bidirectional
rlabel metal4 s 404004 698000 404604 709560 6 vdda1
port 863 nsew power bidirectional
rlabel metal4 s 368004 698000 368604 709560 6 vdda1
port 864 nsew power bidirectional
rlabel metal4 s 332004 698000 332604 709560 6 vdda1
port 865 nsew power bidirectional
rlabel metal4 s 296004 698000 296604 709560 6 vdda1
port 866 nsew power bidirectional
rlabel metal4 s 260004 698000 260604 709560 6 vdda1
port 867 nsew power bidirectional
rlabel metal4 s 224004 698000 224604 709560 6 vdda1
port 868 nsew power bidirectional
rlabel metal4 s 188004 698000 188604 709560 6 vdda1
port 869 nsew power bidirectional
rlabel metal4 s 152004 698000 152604 709560 6 vdda1
port 870 nsew power bidirectional
rlabel metal4 s 116004 698000 116604 709560 6 vdda1
port 871 nsew power bidirectional
rlabel metal4 s 80004 698000 80604 709560 6 vdda1
port 872 nsew power bidirectional
rlabel metal4 s 44004 698000 44604 709560 6 vdda1
port 873 nsew power bidirectional
rlabel metal4 s 8004 698000 8604 709560 6 vdda1
port 874 nsew power bidirectional
rlabel metal4 s 589080 -4684 589680 708620 6 vdda1
port 875 nsew power bidirectional
rlabel metal4 s -5756 -4684 -5156 708620 4 vdda1
port 876 nsew power bidirectional
rlabel metal4 s 548004 -5624 548604 6000 6 vdda1
port 877 nsew power bidirectional
rlabel metal4 s 512004 -5624 512604 6000 6 vdda1
port 878 nsew power bidirectional
rlabel metal4 s 476004 -5624 476604 6000 6 vdda1
port 879 nsew power bidirectional
rlabel metal4 s 440004 -5624 440604 6000 6 vdda1
port 880 nsew power bidirectional
rlabel metal4 s 404004 -5624 404604 6000 6 vdda1
port 881 nsew power bidirectional
rlabel metal4 s 368004 -5624 368604 6000 6 vdda1
port 882 nsew power bidirectional
rlabel metal4 s 332004 -5624 332604 6000 6 vdda1
port 883 nsew power bidirectional
rlabel metal4 s 296004 -5624 296604 6000 6 vdda1
port 884 nsew power bidirectional
rlabel metal4 s 260004 -5624 260604 6000 6 vdda1
port 885 nsew power bidirectional
rlabel metal4 s 224004 -5624 224604 6000 6 vdda1
port 886 nsew power bidirectional
rlabel metal4 s 188004 -5624 188604 6000 6 vdda1
port 887 nsew power bidirectional
rlabel metal4 s 152004 -5624 152604 6000 6 vdda1
port 888 nsew power bidirectional
rlabel metal4 s 116004 -5624 116604 6000 6 vdda1
port 889 nsew power bidirectional
rlabel metal4 s 80004 -5624 80604 6000 6 vdda1
port 890 nsew power bidirectional
rlabel metal4 s 44004 -5624 44604 6000 6 vdda1
port 891 nsew power bidirectional
rlabel metal4 s 8004 -5624 8604 6000 6 vdda1
port 892 nsew power bidirectional
rlabel metal5 s -5756 708020 589680 708620 6 vdda1
port 893 nsew power bidirectional
rlabel metal5 s -6696 693076 590620 693676 6 vdda1
port 894 nsew power bidirectional
rlabel metal5 s -6696 657076 590620 657676 6 vdda1
port 895 nsew power bidirectional
rlabel metal5 s -6696 621076 590620 621676 6 vdda1
port 896 nsew power bidirectional
rlabel metal5 s -6696 585076 590620 585676 6 vdda1
port 897 nsew power bidirectional
rlabel metal5 s -6696 549076 590620 549676 6 vdda1
port 898 nsew power bidirectional
rlabel metal5 s -6696 513076 590620 513676 6 vdda1
port 899 nsew power bidirectional
rlabel metal5 s -6696 477076 590620 477676 6 vdda1
port 900 nsew power bidirectional
rlabel metal5 s -6696 441076 590620 441676 6 vdda1
port 901 nsew power bidirectional
rlabel metal5 s -6696 405076 590620 405676 6 vdda1
port 902 nsew power bidirectional
rlabel metal5 s -6696 369076 590620 369676 6 vdda1
port 903 nsew power bidirectional
rlabel metal5 s -6696 333076 590620 333676 6 vdda1
port 904 nsew power bidirectional
rlabel metal5 s -6696 297076 590620 297676 6 vdda1
port 905 nsew power bidirectional
rlabel metal5 s -6696 261076 590620 261676 6 vdda1
port 906 nsew power bidirectional
rlabel metal5 s -6696 225076 590620 225676 6 vdda1
port 907 nsew power bidirectional
rlabel metal5 s -6696 189076 590620 189676 6 vdda1
port 908 nsew power bidirectional
rlabel metal5 s -6696 153076 590620 153676 6 vdda1
port 909 nsew power bidirectional
rlabel metal5 s -6696 117076 590620 117676 6 vdda1
port 910 nsew power bidirectional
rlabel metal5 s -6696 81076 590620 81676 6 vdda1
port 911 nsew power bidirectional
rlabel metal5 s -6696 45076 590620 45676 6 vdda1
port 912 nsew power bidirectional
rlabel metal5 s -6696 9076 590620 9676 6 vdda1
port 913 nsew power bidirectional
rlabel metal5 s -5756 -4684 589680 -4084 8 vdda1
port 914 nsew power bidirectional
rlabel metal4 s 590020 -5624 590620 709560 6 vssa1
port 915 nsew ground bidirectional
rlabel metal4 s 566004 698000 566604 709560 6 vssa1
port 916 nsew ground bidirectional
rlabel metal4 s 530004 698000 530604 709560 6 vssa1
port 917 nsew ground bidirectional
rlabel metal4 s 494004 698000 494604 709560 6 vssa1
port 918 nsew ground bidirectional
rlabel metal4 s 458004 698000 458604 709560 6 vssa1
port 919 nsew ground bidirectional
rlabel metal4 s 422004 698000 422604 709560 6 vssa1
port 920 nsew ground bidirectional
rlabel metal4 s 386004 698000 386604 709560 6 vssa1
port 921 nsew ground bidirectional
rlabel metal4 s 350004 698000 350604 709560 6 vssa1
port 922 nsew ground bidirectional
rlabel metal4 s 314004 698000 314604 709560 6 vssa1
port 923 nsew ground bidirectional
rlabel metal4 s 278004 698000 278604 709560 6 vssa1
port 924 nsew ground bidirectional
rlabel metal4 s 242004 698000 242604 709560 6 vssa1
port 925 nsew ground bidirectional
rlabel metal4 s 206004 698000 206604 709560 6 vssa1
port 926 nsew ground bidirectional
rlabel metal4 s 170004 698000 170604 709560 6 vssa1
port 927 nsew ground bidirectional
rlabel metal4 s 134004 698000 134604 709560 6 vssa1
port 928 nsew ground bidirectional
rlabel metal4 s 98004 698000 98604 709560 6 vssa1
port 929 nsew ground bidirectional
rlabel metal4 s 62004 698000 62604 709560 6 vssa1
port 930 nsew ground bidirectional
rlabel metal4 s 26004 698000 26604 709560 6 vssa1
port 931 nsew ground bidirectional
rlabel metal4 s -6696 -5624 -6096 709560 4 vssa1
port 932 nsew ground bidirectional
rlabel metal4 s 566004 -5624 566604 6000 6 vssa1
port 933 nsew ground bidirectional
rlabel metal4 s 530004 -5624 530604 6000 6 vssa1
port 934 nsew ground bidirectional
rlabel metal4 s 494004 -5624 494604 6000 6 vssa1
port 935 nsew ground bidirectional
rlabel metal4 s 458004 -5624 458604 6000 6 vssa1
port 936 nsew ground bidirectional
rlabel metal4 s 422004 -5624 422604 6000 6 vssa1
port 937 nsew ground bidirectional
rlabel metal4 s 386004 -5624 386604 6000 6 vssa1
port 938 nsew ground bidirectional
rlabel metal4 s 350004 -5624 350604 6000 6 vssa1
port 939 nsew ground bidirectional
rlabel metal4 s 314004 -5624 314604 6000 6 vssa1
port 940 nsew ground bidirectional
rlabel metal4 s 278004 -5624 278604 6000 6 vssa1
port 941 nsew ground bidirectional
rlabel metal4 s 242004 -5624 242604 6000 6 vssa1
port 942 nsew ground bidirectional
rlabel metal4 s 206004 -5624 206604 6000 6 vssa1
port 943 nsew ground bidirectional
rlabel metal4 s 170004 -5624 170604 6000 6 vssa1
port 944 nsew ground bidirectional
rlabel metal4 s 134004 -5624 134604 6000 6 vssa1
port 945 nsew ground bidirectional
rlabel metal4 s 98004 -5624 98604 6000 6 vssa1
port 946 nsew ground bidirectional
rlabel metal4 s 62004 -5624 62604 6000 6 vssa1
port 947 nsew ground bidirectional
rlabel metal4 s 26004 -5624 26604 6000 6 vssa1
port 948 nsew ground bidirectional
rlabel metal5 s -6696 708960 590620 709560 6 vssa1
port 949 nsew ground bidirectional
rlabel metal5 s -6696 675076 590620 675676 6 vssa1
port 950 nsew ground bidirectional
rlabel metal5 s -6696 639076 590620 639676 6 vssa1
port 951 nsew ground bidirectional
rlabel metal5 s -6696 603076 590620 603676 6 vssa1
port 952 nsew ground bidirectional
rlabel metal5 s -6696 567076 590620 567676 6 vssa1
port 953 nsew ground bidirectional
rlabel metal5 s -6696 531076 590620 531676 6 vssa1
port 954 nsew ground bidirectional
rlabel metal5 s -6696 495076 590620 495676 6 vssa1
port 955 nsew ground bidirectional
rlabel metal5 s -6696 459076 590620 459676 6 vssa1
port 956 nsew ground bidirectional
rlabel metal5 s -6696 423076 590620 423676 6 vssa1
port 957 nsew ground bidirectional
rlabel metal5 s -6696 387076 590620 387676 6 vssa1
port 958 nsew ground bidirectional
rlabel metal5 s -6696 351076 590620 351676 6 vssa1
port 959 nsew ground bidirectional
rlabel metal5 s -6696 315076 590620 315676 6 vssa1
port 960 nsew ground bidirectional
rlabel metal5 s -6696 279076 590620 279676 6 vssa1
port 961 nsew ground bidirectional
rlabel metal5 s -6696 243076 590620 243676 6 vssa1
port 962 nsew ground bidirectional
rlabel metal5 s -6696 207076 590620 207676 6 vssa1
port 963 nsew ground bidirectional
rlabel metal5 s -6696 171076 590620 171676 6 vssa1
port 964 nsew ground bidirectional
rlabel metal5 s -6696 135076 590620 135676 6 vssa1
port 965 nsew ground bidirectional
rlabel metal5 s -6696 99076 590620 99676 6 vssa1
port 966 nsew ground bidirectional
rlabel metal5 s -6696 63076 590620 63676 6 vssa1
port 967 nsew ground bidirectional
rlabel metal5 s -6696 27076 590620 27676 6 vssa1
port 968 nsew ground bidirectional
rlabel metal5 s -6696 -5624 590620 -5024 8 vssa1
port 969 nsew ground bidirectional
rlabel metal4 s 551604 698000 552204 711440 6 vdda2
port 970 nsew power bidirectional
rlabel metal4 s 515604 698000 516204 711440 6 vdda2
port 971 nsew power bidirectional
rlabel metal4 s 479604 698000 480204 711440 6 vdda2
port 972 nsew power bidirectional
rlabel metal4 s 443604 698000 444204 711440 6 vdda2
port 973 nsew power bidirectional
rlabel metal4 s 407604 698000 408204 711440 6 vdda2
port 974 nsew power bidirectional
rlabel metal4 s 371604 698000 372204 711440 6 vdda2
port 975 nsew power bidirectional
rlabel metal4 s 335604 698000 336204 711440 6 vdda2
port 976 nsew power bidirectional
rlabel metal4 s 299604 698000 300204 711440 6 vdda2
port 977 nsew power bidirectional
rlabel metal4 s 263604 698000 264204 711440 6 vdda2
port 978 nsew power bidirectional
rlabel metal4 s 227604 698000 228204 711440 6 vdda2
port 979 nsew power bidirectional
rlabel metal4 s 191604 698000 192204 711440 6 vdda2
port 980 nsew power bidirectional
rlabel metal4 s 155604 698000 156204 711440 6 vdda2
port 981 nsew power bidirectional
rlabel metal4 s 119604 698000 120204 711440 6 vdda2
port 982 nsew power bidirectional
rlabel metal4 s 83604 698000 84204 711440 6 vdda2
port 983 nsew power bidirectional
rlabel metal4 s 47604 698000 48204 711440 6 vdda2
port 984 nsew power bidirectional
rlabel metal4 s 11604 698000 12204 711440 6 vdda2
port 985 nsew power bidirectional
rlabel metal4 s 590960 -6564 591560 710500 6 vdda2
port 986 nsew power bidirectional
rlabel metal4 s -7636 -6564 -7036 710500 4 vdda2
port 987 nsew power bidirectional
rlabel metal4 s 551604 -7504 552204 6000 8 vdda2
port 988 nsew power bidirectional
rlabel metal4 s 515604 -7504 516204 6000 8 vdda2
port 989 nsew power bidirectional
rlabel metal4 s 479604 -7504 480204 6000 8 vdda2
port 990 nsew power bidirectional
rlabel metal4 s 443604 -7504 444204 6000 8 vdda2
port 991 nsew power bidirectional
rlabel metal4 s 407604 -7504 408204 6000 8 vdda2
port 992 nsew power bidirectional
rlabel metal4 s 371604 -7504 372204 6000 8 vdda2
port 993 nsew power bidirectional
rlabel metal4 s 335604 -7504 336204 6000 8 vdda2
port 994 nsew power bidirectional
rlabel metal4 s 299604 -7504 300204 6000 8 vdda2
port 995 nsew power bidirectional
rlabel metal4 s 263604 -7504 264204 6000 8 vdda2
port 996 nsew power bidirectional
rlabel metal4 s 227604 -7504 228204 6000 8 vdda2
port 997 nsew power bidirectional
rlabel metal4 s 191604 -7504 192204 6000 8 vdda2
port 998 nsew power bidirectional
rlabel metal4 s 155604 -7504 156204 6000 8 vdda2
port 999 nsew power bidirectional
rlabel metal4 s 119604 -7504 120204 6000 8 vdda2
port 1000 nsew power bidirectional
rlabel metal4 s 83604 -7504 84204 6000 8 vdda2
port 1001 nsew power bidirectional
rlabel metal4 s 47604 -7504 48204 6000 8 vdda2
port 1002 nsew power bidirectional
rlabel metal4 s 11604 -7504 12204 6000 8 vdda2
port 1003 nsew power bidirectional
rlabel metal5 s -7636 709900 591560 710500 6 vdda2
port 1004 nsew power bidirectional
rlabel metal5 s -8576 696676 592500 697276 6 vdda2
port 1005 nsew power bidirectional
rlabel metal5 s -8576 660676 592500 661276 6 vdda2
port 1006 nsew power bidirectional
rlabel metal5 s -8576 624676 592500 625276 6 vdda2
port 1007 nsew power bidirectional
rlabel metal5 s -8576 588676 592500 589276 6 vdda2
port 1008 nsew power bidirectional
rlabel metal5 s -8576 552676 592500 553276 6 vdda2
port 1009 nsew power bidirectional
rlabel metal5 s -8576 516676 592500 517276 6 vdda2
port 1010 nsew power bidirectional
rlabel metal5 s -8576 480676 592500 481276 6 vdda2
port 1011 nsew power bidirectional
rlabel metal5 s -8576 444676 592500 445276 6 vdda2
port 1012 nsew power bidirectional
rlabel metal5 s -8576 408676 592500 409276 6 vdda2
port 1013 nsew power bidirectional
rlabel metal5 s -8576 372676 592500 373276 6 vdda2
port 1014 nsew power bidirectional
rlabel metal5 s -8576 336676 592500 337276 6 vdda2
port 1015 nsew power bidirectional
rlabel metal5 s -8576 300676 592500 301276 6 vdda2
port 1016 nsew power bidirectional
rlabel metal5 s -8576 264676 592500 265276 6 vdda2
port 1017 nsew power bidirectional
rlabel metal5 s -8576 228676 592500 229276 6 vdda2
port 1018 nsew power bidirectional
rlabel metal5 s -8576 192676 592500 193276 6 vdda2
port 1019 nsew power bidirectional
rlabel metal5 s -8576 156676 592500 157276 6 vdda2
port 1020 nsew power bidirectional
rlabel metal5 s -8576 120676 592500 121276 6 vdda2
port 1021 nsew power bidirectional
rlabel metal5 s -8576 84676 592500 85276 6 vdda2
port 1022 nsew power bidirectional
rlabel metal5 s -8576 48676 592500 49276 6 vdda2
port 1023 nsew power bidirectional
rlabel metal5 s -8576 12676 592500 13276 6 vdda2
port 1024 nsew power bidirectional
rlabel metal5 s -7636 -6564 591560 -5964 8 vdda2
port 1025 nsew power bidirectional
rlabel metal4 s 591900 -7504 592500 711440 6 vssa2
port 1026 nsew ground bidirectional
rlabel metal4 s 569604 698000 570204 711440 6 vssa2
port 1027 nsew ground bidirectional
rlabel metal4 s 533604 698000 534204 711440 6 vssa2
port 1028 nsew ground bidirectional
rlabel metal4 s 497604 698000 498204 711440 6 vssa2
port 1029 nsew ground bidirectional
rlabel metal4 s 461604 698000 462204 711440 6 vssa2
port 1030 nsew ground bidirectional
rlabel metal4 s 425604 698000 426204 711440 6 vssa2
port 1031 nsew ground bidirectional
rlabel metal4 s 389604 698000 390204 711440 6 vssa2
port 1032 nsew ground bidirectional
rlabel metal4 s 353604 698000 354204 711440 6 vssa2
port 1033 nsew ground bidirectional
rlabel metal4 s 317604 698000 318204 711440 6 vssa2
port 1034 nsew ground bidirectional
rlabel metal4 s 281604 698000 282204 711440 6 vssa2
port 1035 nsew ground bidirectional
rlabel metal4 s 245604 698000 246204 711440 6 vssa2
port 1036 nsew ground bidirectional
rlabel metal4 s 209604 698000 210204 711440 6 vssa2
port 1037 nsew ground bidirectional
rlabel metal4 s 173604 698000 174204 711440 6 vssa2
port 1038 nsew ground bidirectional
rlabel metal4 s 137604 698000 138204 711440 6 vssa2
port 1039 nsew ground bidirectional
rlabel metal4 s 101604 698000 102204 711440 6 vssa2
port 1040 nsew ground bidirectional
rlabel metal4 s 65604 698000 66204 711440 6 vssa2
port 1041 nsew ground bidirectional
rlabel metal4 s 29604 698000 30204 711440 6 vssa2
port 1042 nsew ground bidirectional
rlabel metal4 s -8576 -7504 -7976 711440 4 vssa2
port 1043 nsew ground bidirectional
rlabel metal4 s 569604 -7504 570204 6000 8 vssa2
port 1044 nsew ground bidirectional
rlabel metal4 s 533604 -7504 534204 6000 8 vssa2
port 1045 nsew ground bidirectional
rlabel metal4 s 497604 -7504 498204 6000 8 vssa2
port 1046 nsew ground bidirectional
rlabel metal4 s 461604 -7504 462204 6000 8 vssa2
port 1047 nsew ground bidirectional
rlabel metal4 s 425604 -7504 426204 6000 8 vssa2
port 1048 nsew ground bidirectional
rlabel metal4 s 389604 -7504 390204 6000 8 vssa2
port 1049 nsew ground bidirectional
rlabel metal4 s 353604 -7504 354204 6000 8 vssa2
port 1050 nsew ground bidirectional
rlabel metal4 s 317604 -7504 318204 6000 8 vssa2
port 1051 nsew ground bidirectional
rlabel metal4 s 281604 -7504 282204 6000 8 vssa2
port 1052 nsew ground bidirectional
rlabel metal4 s 245604 -7504 246204 6000 8 vssa2
port 1053 nsew ground bidirectional
rlabel metal4 s 209604 -7504 210204 6000 8 vssa2
port 1054 nsew ground bidirectional
rlabel metal4 s 173604 -7504 174204 6000 8 vssa2
port 1055 nsew ground bidirectional
rlabel metal4 s 137604 -7504 138204 6000 8 vssa2
port 1056 nsew ground bidirectional
rlabel metal4 s 101604 -7504 102204 6000 8 vssa2
port 1057 nsew ground bidirectional
rlabel metal4 s 65604 -7504 66204 6000 8 vssa2
port 1058 nsew ground bidirectional
rlabel metal4 s 29604 -7504 30204 6000 8 vssa2
port 1059 nsew ground bidirectional
rlabel metal5 s -8576 710840 592500 711440 6 vssa2
port 1060 nsew ground bidirectional
rlabel metal5 s -8576 678676 592500 679276 6 vssa2
port 1061 nsew ground bidirectional
rlabel metal5 s -8576 642676 592500 643276 6 vssa2
port 1062 nsew ground bidirectional
rlabel metal5 s -8576 606676 592500 607276 6 vssa2
port 1063 nsew ground bidirectional
rlabel metal5 s -8576 570676 592500 571276 6 vssa2
port 1064 nsew ground bidirectional
rlabel metal5 s -8576 534676 592500 535276 6 vssa2
port 1065 nsew ground bidirectional
rlabel metal5 s -8576 498676 592500 499276 6 vssa2
port 1066 nsew ground bidirectional
rlabel metal5 s -8576 462676 592500 463276 6 vssa2
port 1067 nsew ground bidirectional
rlabel metal5 s -8576 426676 592500 427276 6 vssa2
port 1068 nsew ground bidirectional
rlabel metal5 s -8576 390676 592500 391276 6 vssa2
port 1069 nsew ground bidirectional
rlabel metal5 s -8576 354676 592500 355276 6 vssa2
port 1070 nsew ground bidirectional
rlabel metal5 s -8576 318676 592500 319276 6 vssa2
port 1071 nsew ground bidirectional
rlabel metal5 s -8576 282676 592500 283276 6 vssa2
port 1072 nsew ground bidirectional
rlabel metal5 s -8576 246676 592500 247276 6 vssa2
port 1073 nsew ground bidirectional
rlabel metal5 s -8576 210676 592500 211276 6 vssa2
port 1074 nsew ground bidirectional
rlabel metal5 s -8576 174676 592500 175276 6 vssa2
port 1075 nsew ground bidirectional
rlabel metal5 s -8576 138676 592500 139276 6 vssa2
port 1076 nsew ground bidirectional
rlabel metal5 s -8576 102676 592500 103276 6 vssa2
port 1077 nsew ground bidirectional
rlabel metal5 s -8576 66676 592500 67276 6 vssa2
port 1078 nsew ground bidirectional
rlabel metal5 s -8576 30676 592500 31276 6 vssa2
port 1079 nsew ground bidirectional
rlabel metal5 s -8576 -7504 592500 -6904 8 vssa2
port 1080 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1608194264
<< obsli1 >>
rect 1104 2159 562856 681649
<< obsm1 >>
rect 566 1164 562856 681680
<< metal2 >>
rect 2318 683200 2374 684000
rect 6918 683200 6974 684000
rect 11610 683200 11666 684000
rect 16210 683200 16266 684000
rect 20902 683200 20958 684000
rect 25594 683200 25650 684000
rect 30194 683200 30250 684000
rect 34886 683200 34942 684000
rect 39578 683200 39634 684000
rect 44178 683200 44234 684000
rect 48870 683200 48926 684000
rect 53562 683200 53618 684000
rect 58162 683200 58218 684000
rect 62854 683200 62910 684000
rect 67546 683200 67602 684000
rect 72146 683200 72202 684000
rect 76838 683200 76894 684000
rect 81530 683200 81586 684000
rect 86130 683200 86186 684000
rect 90822 683200 90878 684000
rect 95514 683200 95570 684000
rect 100114 683200 100170 684000
rect 104806 683200 104862 684000
rect 109498 683200 109554 684000
rect 114098 683200 114154 684000
rect 118790 683200 118846 684000
rect 123482 683200 123538 684000
rect 128082 683200 128138 684000
rect 132774 683200 132830 684000
rect 137466 683200 137522 684000
rect 142066 683200 142122 684000
rect 146758 683200 146814 684000
rect 151450 683200 151506 684000
rect 156050 683200 156106 684000
rect 160742 683200 160798 684000
rect 165434 683200 165490 684000
rect 170034 683200 170090 684000
rect 174726 683200 174782 684000
rect 179418 683200 179474 684000
rect 184018 683200 184074 684000
rect 188710 683200 188766 684000
rect 193402 683200 193458 684000
rect 198002 683200 198058 684000
rect 202694 683200 202750 684000
rect 207386 683200 207442 684000
rect 211986 683200 212042 684000
rect 216678 683200 216734 684000
rect 221370 683200 221426 684000
rect 225970 683200 226026 684000
rect 230662 683200 230718 684000
rect 235354 683200 235410 684000
rect 239954 683200 240010 684000
rect 244646 683200 244702 684000
rect 249338 683200 249394 684000
rect 253938 683200 253994 684000
rect 258630 683200 258686 684000
rect 263322 683200 263378 684000
rect 267922 683200 267978 684000
rect 272614 683200 272670 684000
rect 277306 683200 277362 684000
rect 281906 683200 281962 684000
rect 286598 683200 286654 684000
rect 291198 683200 291254 684000
rect 295890 683200 295946 684000
rect 300582 683200 300638 684000
rect 305182 683200 305238 684000
rect 309874 683200 309930 684000
rect 314566 683200 314622 684000
rect 319166 683200 319222 684000
rect 323858 683200 323914 684000
rect 328550 683200 328606 684000
rect 333150 683200 333206 684000
rect 337842 683200 337898 684000
rect 342534 683200 342590 684000
rect 347134 683200 347190 684000
rect 351826 683200 351882 684000
rect 356518 683200 356574 684000
rect 361118 683200 361174 684000
rect 365810 683200 365866 684000
rect 370502 683200 370558 684000
rect 375102 683200 375158 684000
rect 379794 683200 379850 684000
rect 384486 683200 384542 684000
rect 389086 683200 389142 684000
rect 393778 683200 393834 684000
rect 398470 683200 398526 684000
rect 403070 683200 403126 684000
rect 407762 683200 407818 684000
rect 412454 683200 412510 684000
rect 417054 683200 417110 684000
rect 421746 683200 421802 684000
rect 426438 683200 426494 684000
rect 431038 683200 431094 684000
rect 435730 683200 435786 684000
rect 440422 683200 440478 684000
rect 445022 683200 445078 684000
rect 449714 683200 449770 684000
rect 454406 683200 454462 684000
rect 459006 683200 459062 684000
rect 463698 683200 463754 684000
rect 468390 683200 468446 684000
rect 472990 683200 473046 684000
rect 477682 683200 477738 684000
rect 482374 683200 482430 684000
rect 486974 683200 487030 684000
rect 491666 683200 491722 684000
rect 496358 683200 496414 684000
rect 500958 683200 501014 684000
rect 505650 683200 505706 684000
rect 510342 683200 510398 684000
rect 514942 683200 514998 684000
rect 519634 683200 519690 684000
rect 524326 683200 524382 684000
rect 528926 683200 528982 684000
rect 533618 683200 533674 684000
rect 538310 683200 538366 684000
rect 542910 683200 542966 684000
rect 547602 683200 547658 684000
rect 552294 683200 552350 684000
rect 556894 683200 556950 684000
rect 561586 683200 561642 684000
rect 570 0 626 800
rect 1674 0 1730 800
rect 2778 0 2834 800
rect 3882 0 3938 800
rect 4986 0 5042 800
rect 6090 0 6146 800
rect 7194 0 7250 800
rect 8390 0 8446 800
rect 9494 0 9550 800
rect 10598 0 10654 800
rect 11702 0 11758 800
rect 12806 0 12862 800
rect 13910 0 13966 800
rect 15106 0 15162 800
rect 16210 0 16266 800
rect 17314 0 17370 800
rect 18418 0 18474 800
rect 19522 0 19578 800
rect 20626 0 20682 800
rect 21822 0 21878 800
rect 22926 0 22982 800
rect 24030 0 24086 800
rect 25134 0 25190 800
rect 26238 0 26294 800
rect 27342 0 27398 800
rect 28538 0 28594 800
rect 29642 0 29698 800
rect 30746 0 30802 800
rect 31850 0 31906 800
rect 32954 0 33010 800
rect 34058 0 34114 800
rect 35254 0 35310 800
rect 36358 0 36414 800
rect 37462 0 37518 800
rect 38566 0 38622 800
rect 39670 0 39726 800
rect 40774 0 40830 800
rect 41970 0 42026 800
rect 43074 0 43130 800
rect 44178 0 44234 800
rect 45282 0 45338 800
rect 46386 0 46442 800
rect 47490 0 47546 800
rect 48594 0 48650 800
rect 49790 0 49846 800
rect 50894 0 50950 800
rect 51998 0 52054 800
rect 53102 0 53158 800
rect 54206 0 54262 800
rect 55310 0 55366 800
rect 56506 0 56562 800
rect 57610 0 57666 800
rect 58714 0 58770 800
rect 59818 0 59874 800
rect 60922 0 60978 800
rect 62026 0 62082 800
rect 63222 0 63278 800
rect 64326 0 64382 800
rect 65430 0 65486 800
rect 66534 0 66590 800
rect 67638 0 67694 800
rect 68742 0 68798 800
rect 69938 0 69994 800
rect 71042 0 71098 800
rect 72146 0 72202 800
rect 73250 0 73306 800
rect 74354 0 74410 800
rect 75458 0 75514 800
rect 76654 0 76710 800
rect 77758 0 77814 800
rect 78862 0 78918 800
rect 79966 0 80022 800
rect 81070 0 81126 800
rect 82174 0 82230 800
rect 83370 0 83426 800
rect 84474 0 84530 800
rect 85578 0 85634 800
rect 86682 0 86738 800
rect 87786 0 87842 800
rect 88890 0 88946 800
rect 90086 0 90142 800
rect 91190 0 91246 800
rect 92294 0 92350 800
rect 93398 0 93454 800
rect 94502 0 94558 800
rect 95606 0 95662 800
rect 96710 0 96766 800
rect 97906 0 97962 800
rect 99010 0 99066 800
rect 100114 0 100170 800
rect 101218 0 101274 800
rect 102322 0 102378 800
rect 103426 0 103482 800
rect 104622 0 104678 800
rect 105726 0 105782 800
rect 106830 0 106886 800
rect 107934 0 107990 800
rect 109038 0 109094 800
rect 110142 0 110198 800
rect 111338 0 111394 800
rect 112442 0 112498 800
rect 113546 0 113602 800
rect 114650 0 114706 800
rect 115754 0 115810 800
rect 116858 0 116914 800
rect 118054 0 118110 800
rect 119158 0 119214 800
rect 120262 0 120318 800
rect 121366 0 121422 800
rect 122470 0 122526 800
rect 123574 0 123630 800
rect 124770 0 124826 800
rect 125874 0 125930 800
rect 126978 0 127034 800
rect 128082 0 128138 800
rect 129186 0 129242 800
rect 130290 0 130346 800
rect 131486 0 131542 800
rect 132590 0 132646 800
rect 133694 0 133750 800
rect 134798 0 134854 800
rect 135902 0 135958 800
rect 137006 0 137062 800
rect 138202 0 138258 800
rect 139306 0 139362 800
rect 140410 0 140466 800
rect 141514 0 141570 800
rect 142618 0 142674 800
rect 143722 0 143778 800
rect 144826 0 144882 800
rect 146022 0 146078 800
rect 147126 0 147182 800
rect 148230 0 148286 800
rect 149334 0 149390 800
rect 150438 0 150494 800
rect 151542 0 151598 800
rect 152738 0 152794 800
rect 153842 0 153898 800
rect 154946 0 155002 800
rect 156050 0 156106 800
rect 157154 0 157210 800
rect 158258 0 158314 800
rect 159454 0 159510 800
rect 160558 0 160614 800
rect 161662 0 161718 800
rect 162766 0 162822 800
rect 163870 0 163926 800
rect 164974 0 165030 800
rect 166170 0 166226 800
rect 167274 0 167330 800
rect 168378 0 168434 800
rect 169482 0 169538 800
rect 170586 0 170642 800
rect 171690 0 171746 800
rect 172886 0 172942 800
rect 173990 0 174046 800
rect 175094 0 175150 800
rect 176198 0 176254 800
rect 177302 0 177358 800
rect 178406 0 178462 800
rect 179602 0 179658 800
rect 180706 0 180762 800
rect 181810 0 181866 800
rect 182914 0 182970 800
rect 184018 0 184074 800
rect 185122 0 185178 800
rect 186318 0 186374 800
rect 187422 0 187478 800
rect 188526 0 188582 800
rect 189630 0 189686 800
rect 190734 0 190790 800
rect 191838 0 191894 800
rect 192942 0 192998 800
rect 194138 0 194194 800
rect 195242 0 195298 800
rect 196346 0 196402 800
rect 197450 0 197506 800
rect 198554 0 198610 800
rect 199658 0 199714 800
rect 200854 0 200910 800
rect 201958 0 202014 800
rect 203062 0 203118 800
rect 204166 0 204222 800
rect 205270 0 205326 800
rect 206374 0 206430 800
rect 207570 0 207626 800
rect 208674 0 208730 800
rect 209778 0 209834 800
rect 210882 0 210938 800
rect 211986 0 212042 800
rect 213090 0 213146 800
rect 214286 0 214342 800
rect 215390 0 215446 800
rect 216494 0 216550 800
rect 217598 0 217654 800
rect 218702 0 218758 800
rect 219806 0 219862 800
rect 221002 0 221058 800
rect 222106 0 222162 800
rect 223210 0 223266 800
rect 224314 0 224370 800
rect 225418 0 225474 800
rect 226522 0 226578 800
rect 227718 0 227774 800
rect 228822 0 228878 800
rect 229926 0 229982 800
rect 231030 0 231086 800
rect 232134 0 232190 800
rect 233238 0 233294 800
rect 234434 0 234490 800
rect 235538 0 235594 800
rect 236642 0 236698 800
rect 237746 0 237802 800
rect 238850 0 238906 800
rect 239954 0 240010 800
rect 241058 0 241114 800
rect 242254 0 242310 800
rect 243358 0 243414 800
rect 244462 0 244518 800
rect 245566 0 245622 800
rect 246670 0 246726 800
rect 247774 0 247830 800
rect 248970 0 249026 800
rect 250074 0 250130 800
rect 251178 0 251234 800
rect 252282 0 252338 800
rect 253386 0 253442 800
rect 254490 0 254546 800
rect 255686 0 255742 800
rect 256790 0 256846 800
rect 257894 0 257950 800
rect 258998 0 259054 800
rect 260102 0 260158 800
rect 261206 0 261262 800
rect 262402 0 262458 800
rect 263506 0 263562 800
rect 264610 0 264666 800
rect 265714 0 265770 800
rect 266818 0 266874 800
rect 267922 0 267978 800
rect 269118 0 269174 800
rect 270222 0 270278 800
rect 271326 0 271382 800
rect 272430 0 272486 800
rect 273534 0 273590 800
rect 274638 0 274694 800
rect 275834 0 275890 800
rect 276938 0 276994 800
rect 278042 0 278098 800
rect 279146 0 279202 800
rect 280250 0 280306 800
rect 281354 0 281410 800
rect 282550 0 282606 800
rect 283654 0 283710 800
rect 284758 0 284814 800
rect 285862 0 285918 800
rect 286966 0 287022 800
rect 288070 0 288126 800
rect 289174 0 289230 800
rect 290370 0 290426 800
rect 291474 0 291530 800
rect 292578 0 292634 800
rect 293682 0 293738 800
rect 294786 0 294842 800
rect 295890 0 295946 800
rect 297086 0 297142 800
rect 298190 0 298246 800
rect 299294 0 299350 800
rect 300398 0 300454 800
rect 301502 0 301558 800
rect 302606 0 302662 800
rect 303802 0 303858 800
rect 304906 0 304962 800
rect 306010 0 306066 800
rect 307114 0 307170 800
rect 308218 0 308274 800
rect 309322 0 309378 800
rect 310518 0 310574 800
rect 311622 0 311678 800
rect 312726 0 312782 800
rect 313830 0 313886 800
rect 314934 0 314990 800
rect 316038 0 316094 800
rect 317234 0 317290 800
rect 318338 0 318394 800
rect 319442 0 319498 800
rect 320546 0 320602 800
rect 321650 0 321706 800
rect 322754 0 322810 800
rect 323950 0 324006 800
rect 325054 0 325110 800
rect 326158 0 326214 800
rect 327262 0 327318 800
rect 328366 0 328422 800
rect 329470 0 329526 800
rect 330574 0 330630 800
rect 331770 0 331826 800
rect 332874 0 332930 800
rect 333978 0 334034 800
rect 335082 0 335138 800
rect 336186 0 336242 800
rect 337290 0 337346 800
rect 338486 0 338542 800
rect 339590 0 339646 800
rect 340694 0 340750 800
rect 341798 0 341854 800
rect 342902 0 342958 800
rect 344006 0 344062 800
rect 345202 0 345258 800
rect 346306 0 346362 800
rect 347410 0 347466 800
rect 348514 0 348570 800
rect 349618 0 349674 800
rect 350722 0 350778 800
rect 351918 0 351974 800
rect 353022 0 353078 800
rect 354126 0 354182 800
rect 355230 0 355286 800
rect 356334 0 356390 800
rect 357438 0 357494 800
rect 358634 0 358690 800
rect 359738 0 359794 800
rect 360842 0 360898 800
rect 361946 0 362002 800
rect 363050 0 363106 800
rect 364154 0 364210 800
rect 365350 0 365406 800
rect 366454 0 366510 800
rect 367558 0 367614 800
rect 368662 0 368718 800
rect 369766 0 369822 800
rect 370870 0 370926 800
rect 372066 0 372122 800
rect 373170 0 373226 800
rect 374274 0 374330 800
rect 375378 0 375434 800
rect 376482 0 376538 800
rect 377586 0 377642 800
rect 378690 0 378746 800
rect 379886 0 379942 800
rect 380990 0 381046 800
rect 382094 0 382150 800
rect 383198 0 383254 800
rect 384302 0 384358 800
rect 385406 0 385462 800
rect 386602 0 386658 800
rect 387706 0 387762 800
rect 388810 0 388866 800
rect 389914 0 389970 800
rect 391018 0 391074 800
rect 392122 0 392178 800
rect 393318 0 393374 800
rect 394422 0 394478 800
rect 395526 0 395582 800
rect 396630 0 396686 800
rect 397734 0 397790 800
rect 398838 0 398894 800
rect 400034 0 400090 800
rect 401138 0 401194 800
rect 402242 0 402298 800
rect 403346 0 403402 800
rect 404450 0 404506 800
rect 405554 0 405610 800
rect 406750 0 406806 800
rect 407854 0 407910 800
rect 408958 0 409014 800
rect 410062 0 410118 800
rect 411166 0 411222 800
rect 412270 0 412326 800
rect 413466 0 413522 800
rect 414570 0 414626 800
rect 415674 0 415730 800
rect 416778 0 416834 800
rect 417882 0 417938 800
rect 418986 0 419042 800
rect 420182 0 420238 800
rect 421286 0 421342 800
rect 422390 0 422446 800
rect 423494 0 423550 800
rect 424598 0 424654 800
rect 425702 0 425758 800
rect 426806 0 426862 800
rect 428002 0 428058 800
rect 429106 0 429162 800
rect 430210 0 430266 800
rect 431314 0 431370 800
rect 432418 0 432474 800
rect 433522 0 433578 800
rect 434718 0 434774 800
rect 435822 0 435878 800
rect 436926 0 436982 800
rect 438030 0 438086 800
rect 439134 0 439190 800
rect 440238 0 440294 800
rect 441434 0 441490 800
rect 442538 0 442594 800
rect 443642 0 443698 800
rect 444746 0 444802 800
rect 445850 0 445906 800
rect 446954 0 447010 800
rect 448150 0 448206 800
rect 449254 0 449310 800
rect 450358 0 450414 800
rect 451462 0 451518 800
rect 452566 0 452622 800
rect 453670 0 453726 800
rect 454866 0 454922 800
rect 455970 0 456026 800
rect 457074 0 457130 800
rect 458178 0 458234 800
rect 459282 0 459338 800
rect 460386 0 460442 800
rect 461582 0 461638 800
rect 462686 0 462742 800
rect 463790 0 463846 800
rect 464894 0 464950 800
rect 465998 0 466054 800
rect 467102 0 467158 800
rect 468298 0 468354 800
rect 469402 0 469458 800
rect 470506 0 470562 800
rect 471610 0 471666 800
rect 472714 0 472770 800
rect 473818 0 473874 800
rect 474922 0 474978 800
rect 476118 0 476174 800
rect 477222 0 477278 800
rect 478326 0 478382 800
rect 479430 0 479486 800
rect 480534 0 480590 800
rect 481638 0 481694 800
rect 482834 0 482890 800
rect 483938 0 483994 800
rect 485042 0 485098 800
rect 486146 0 486202 800
rect 487250 0 487306 800
rect 488354 0 488410 800
rect 489550 0 489606 800
rect 490654 0 490710 800
rect 491758 0 491814 800
rect 492862 0 492918 800
rect 493966 0 494022 800
rect 495070 0 495126 800
rect 496266 0 496322 800
rect 497370 0 497426 800
rect 498474 0 498530 800
rect 499578 0 499634 800
rect 500682 0 500738 800
rect 501786 0 501842 800
rect 502982 0 503038 800
rect 504086 0 504142 800
rect 505190 0 505246 800
rect 506294 0 506350 800
rect 507398 0 507454 800
rect 508502 0 508558 800
rect 509698 0 509754 800
rect 510802 0 510858 800
rect 511906 0 511962 800
rect 513010 0 513066 800
rect 514114 0 514170 800
rect 515218 0 515274 800
rect 516414 0 516470 800
rect 517518 0 517574 800
rect 518622 0 518678 800
rect 519726 0 519782 800
rect 520830 0 520886 800
rect 521934 0 521990 800
rect 523038 0 523094 800
rect 524234 0 524290 800
rect 525338 0 525394 800
rect 526442 0 526498 800
rect 527546 0 527602 800
rect 528650 0 528706 800
rect 529754 0 529810 800
rect 530950 0 531006 800
rect 532054 0 532110 800
rect 533158 0 533214 800
rect 534262 0 534318 800
rect 535366 0 535422 800
rect 536470 0 536526 800
rect 537666 0 537722 800
rect 538770 0 538826 800
rect 539874 0 539930 800
rect 540978 0 541034 800
rect 542082 0 542138 800
rect 543186 0 543242 800
rect 544382 0 544438 800
rect 545486 0 545542 800
rect 546590 0 546646 800
rect 547694 0 547750 800
rect 548798 0 548854 800
rect 549902 0 549958 800
rect 551098 0 551154 800
rect 552202 0 552258 800
rect 553306 0 553362 800
rect 554410 0 554466 800
rect 555514 0 555570 800
rect 556618 0 556674 800
rect 557814 0 557870 800
rect 558918 0 558974 800
rect 560022 0 560078 800
rect 561126 0 561182 800
rect 562230 0 562286 800
rect 563334 0 563390 800
<< obsm2 >>
rect 572 683144 2262 683200
rect 2430 683144 6862 683200
rect 7030 683144 11554 683200
rect 11722 683144 16154 683200
rect 16322 683144 20846 683200
rect 21014 683144 25538 683200
rect 25706 683144 30138 683200
rect 30306 683144 34830 683200
rect 34998 683144 39522 683200
rect 39690 683144 44122 683200
rect 44290 683144 48814 683200
rect 48982 683144 53506 683200
rect 53674 683144 58106 683200
rect 58274 683144 62798 683200
rect 62966 683144 67490 683200
rect 67658 683144 72090 683200
rect 72258 683144 76782 683200
rect 76950 683144 81474 683200
rect 81642 683144 86074 683200
rect 86242 683144 90766 683200
rect 90934 683144 95458 683200
rect 95626 683144 100058 683200
rect 100226 683144 104750 683200
rect 104918 683144 109442 683200
rect 109610 683144 114042 683200
rect 114210 683144 118734 683200
rect 118902 683144 123426 683200
rect 123594 683144 128026 683200
rect 128194 683144 132718 683200
rect 132886 683144 137410 683200
rect 137578 683144 142010 683200
rect 142178 683144 146702 683200
rect 146870 683144 151394 683200
rect 151562 683144 155994 683200
rect 156162 683144 160686 683200
rect 160854 683144 165378 683200
rect 165546 683144 169978 683200
rect 170146 683144 174670 683200
rect 174838 683144 179362 683200
rect 179530 683144 183962 683200
rect 184130 683144 188654 683200
rect 188822 683144 193346 683200
rect 193514 683144 197946 683200
rect 198114 683144 202638 683200
rect 202806 683144 207330 683200
rect 207498 683144 211930 683200
rect 212098 683144 216622 683200
rect 216790 683144 221314 683200
rect 221482 683144 225914 683200
rect 226082 683144 230606 683200
rect 230774 683144 235298 683200
rect 235466 683144 239898 683200
rect 240066 683144 244590 683200
rect 244758 683144 249282 683200
rect 249450 683144 253882 683200
rect 254050 683144 258574 683200
rect 258742 683144 263266 683200
rect 263434 683144 267866 683200
rect 268034 683144 272558 683200
rect 272726 683144 277250 683200
rect 277418 683144 281850 683200
rect 282018 683144 286542 683200
rect 286710 683144 291142 683200
rect 291310 683144 295834 683200
rect 296002 683144 300526 683200
rect 300694 683144 305126 683200
rect 305294 683144 309818 683200
rect 309986 683144 314510 683200
rect 314678 683144 319110 683200
rect 319278 683144 323802 683200
rect 323970 683144 328494 683200
rect 328662 683144 333094 683200
rect 333262 683144 337786 683200
rect 337954 683144 342478 683200
rect 342646 683144 347078 683200
rect 347246 683144 351770 683200
rect 351938 683144 356462 683200
rect 356630 683144 361062 683200
rect 361230 683144 365754 683200
rect 365922 683144 370446 683200
rect 370614 683144 375046 683200
rect 375214 683144 379738 683200
rect 379906 683144 384430 683200
rect 384598 683144 389030 683200
rect 389198 683144 393722 683200
rect 393890 683144 398414 683200
rect 398582 683144 403014 683200
rect 403182 683144 407706 683200
rect 407874 683144 412398 683200
rect 412566 683144 416998 683200
rect 417166 683144 421690 683200
rect 421858 683144 426382 683200
rect 426550 683144 430982 683200
rect 431150 683144 435674 683200
rect 435842 683144 440366 683200
rect 440534 683144 444966 683200
rect 445134 683144 449658 683200
rect 449826 683144 454350 683200
rect 454518 683144 458950 683200
rect 459118 683144 463642 683200
rect 463810 683144 468334 683200
rect 468502 683144 472934 683200
rect 473102 683144 477626 683200
rect 477794 683144 482318 683200
rect 482486 683144 486918 683200
rect 487086 683144 491610 683200
rect 491778 683144 496302 683200
rect 496470 683144 500902 683200
rect 501070 683144 505594 683200
rect 505762 683144 510286 683200
rect 510454 683144 514886 683200
rect 515054 683144 519578 683200
rect 519746 683144 524270 683200
rect 524438 683144 528870 683200
rect 529038 683144 533562 683200
rect 533730 683144 538254 683200
rect 538422 683144 542854 683200
rect 543022 683144 547546 683200
rect 547714 683144 552238 683200
rect 552406 683144 556838 683200
rect 557006 683144 557476 683200
rect 572 856 557476 683144
rect 682 800 1618 856
rect 1786 800 2722 856
rect 2890 800 3826 856
rect 3994 800 4930 856
rect 5098 800 6034 856
rect 6202 800 7138 856
rect 7306 800 8334 856
rect 8502 800 9438 856
rect 9606 800 10542 856
rect 10710 800 11646 856
rect 11814 800 12750 856
rect 12918 800 13854 856
rect 14022 800 15050 856
rect 15218 800 16154 856
rect 16322 800 17258 856
rect 17426 800 18362 856
rect 18530 800 19466 856
rect 19634 800 20570 856
rect 20738 800 21766 856
rect 21934 800 22870 856
rect 23038 800 23974 856
rect 24142 800 25078 856
rect 25246 800 26182 856
rect 26350 800 27286 856
rect 27454 800 28482 856
rect 28650 800 29586 856
rect 29754 800 30690 856
rect 30858 800 31794 856
rect 31962 800 32898 856
rect 33066 800 34002 856
rect 34170 800 35198 856
rect 35366 800 36302 856
rect 36470 800 37406 856
rect 37574 800 38510 856
rect 38678 800 39614 856
rect 39782 800 40718 856
rect 40886 800 41914 856
rect 42082 800 43018 856
rect 43186 800 44122 856
rect 44290 800 45226 856
rect 45394 800 46330 856
rect 46498 800 47434 856
rect 47602 800 48538 856
rect 48706 800 49734 856
rect 49902 800 50838 856
rect 51006 800 51942 856
rect 52110 800 53046 856
rect 53214 800 54150 856
rect 54318 800 55254 856
rect 55422 800 56450 856
rect 56618 800 57554 856
rect 57722 800 58658 856
rect 58826 800 59762 856
rect 59930 800 60866 856
rect 61034 800 61970 856
rect 62138 800 63166 856
rect 63334 800 64270 856
rect 64438 800 65374 856
rect 65542 800 66478 856
rect 66646 800 67582 856
rect 67750 800 68686 856
rect 68854 800 69882 856
rect 70050 800 70986 856
rect 71154 800 72090 856
rect 72258 800 73194 856
rect 73362 800 74298 856
rect 74466 800 75402 856
rect 75570 800 76598 856
rect 76766 800 77702 856
rect 77870 800 78806 856
rect 78974 800 79910 856
rect 80078 800 81014 856
rect 81182 800 82118 856
rect 82286 800 83314 856
rect 83482 800 84418 856
rect 84586 800 85522 856
rect 85690 800 86626 856
rect 86794 800 87730 856
rect 87898 800 88834 856
rect 89002 800 90030 856
rect 90198 800 91134 856
rect 91302 800 92238 856
rect 92406 800 93342 856
rect 93510 800 94446 856
rect 94614 800 95550 856
rect 95718 800 96654 856
rect 96822 800 97850 856
rect 98018 800 98954 856
rect 99122 800 100058 856
rect 100226 800 101162 856
rect 101330 800 102266 856
rect 102434 800 103370 856
rect 103538 800 104566 856
rect 104734 800 105670 856
rect 105838 800 106774 856
rect 106942 800 107878 856
rect 108046 800 108982 856
rect 109150 800 110086 856
rect 110254 800 111282 856
rect 111450 800 112386 856
rect 112554 800 113490 856
rect 113658 800 114594 856
rect 114762 800 115698 856
rect 115866 800 116802 856
rect 116970 800 117998 856
rect 118166 800 119102 856
rect 119270 800 120206 856
rect 120374 800 121310 856
rect 121478 800 122414 856
rect 122582 800 123518 856
rect 123686 800 124714 856
rect 124882 800 125818 856
rect 125986 800 126922 856
rect 127090 800 128026 856
rect 128194 800 129130 856
rect 129298 800 130234 856
rect 130402 800 131430 856
rect 131598 800 132534 856
rect 132702 800 133638 856
rect 133806 800 134742 856
rect 134910 800 135846 856
rect 136014 800 136950 856
rect 137118 800 138146 856
rect 138314 800 139250 856
rect 139418 800 140354 856
rect 140522 800 141458 856
rect 141626 800 142562 856
rect 142730 800 143666 856
rect 143834 800 144770 856
rect 144938 800 145966 856
rect 146134 800 147070 856
rect 147238 800 148174 856
rect 148342 800 149278 856
rect 149446 800 150382 856
rect 150550 800 151486 856
rect 151654 800 152682 856
rect 152850 800 153786 856
rect 153954 800 154890 856
rect 155058 800 155994 856
rect 156162 800 157098 856
rect 157266 800 158202 856
rect 158370 800 159398 856
rect 159566 800 160502 856
rect 160670 800 161606 856
rect 161774 800 162710 856
rect 162878 800 163814 856
rect 163982 800 164918 856
rect 165086 800 166114 856
rect 166282 800 167218 856
rect 167386 800 168322 856
rect 168490 800 169426 856
rect 169594 800 170530 856
rect 170698 800 171634 856
rect 171802 800 172830 856
rect 172998 800 173934 856
rect 174102 800 175038 856
rect 175206 800 176142 856
rect 176310 800 177246 856
rect 177414 800 178350 856
rect 178518 800 179546 856
rect 179714 800 180650 856
rect 180818 800 181754 856
rect 181922 800 182858 856
rect 183026 800 183962 856
rect 184130 800 185066 856
rect 185234 800 186262 856
rect 186430 800 187366 856
rect 187534 800 188470 856
rect 188638 800 189574 856
rect 189742 800 190678 856
rect 190846 800 191782 856
rect 191950 800 192886 856
rect 193054 800 194082 856
rect 194250 800 195186 856
rect 195354 800 196290 856
rect 196458 800 197394 856
rect 197562 800 198498 856
rect 198666 800 199602 856
rect 199770 800 200798 856
rect 200966 800 201902 856
rect 202070 800 203006 856
rect 203174 800 204110 856
rect 204278 800 205214 856
rect 205382 800 206318 856
rect 206486 800 207514 856
rect 207682 800 208618 856
rect 208786 800 209722 856
rect 209890 800 210826 856
rect 210994 800 211930 856
rect 212098 800 213034 856
rect 213202 800 214230 856
rect 214398 800 215334 856
rect 215502 800 216438 856
rect 216606 800 217542 856
rect 217710 800 218646 856
rect 218814 800 219750 856
rect 219918 800 220946 856
rect 221114 800 222050 856
rect 222218 800 223154 856
rect 223322 800 224258 856
rect 224426 800 225362 856
rect 225530 800 226466 856
rect 226634 800 227662 856
rect 227830 800 228766 856
rect 228934 800 229870 856
rect 230038 800 230974 856
rect 231142 800 232078 856
rect 232246 800 233182 856
rect 233350 800 234378 856
rect 234546 800 235482 856
rect 235650 800 236586 856
rect 236754 800 237690 856
rect 237858 800 238794 856
rect 238962 800 239898 856
rect 240066 800 241002 856
rect 241170 800 242198 856
rect 242366 800 243302 856
rect 243470 800 244406 856
rect 244574 800 245510 856
rect 245678 800 246614 856
rect 246782 800 247718 856
rect 247886 800 248914 856
rect 249082 800 250018 856
rect 250186 800 251122 856
rect 251290 800 252226 856
rect 252394 800 253330 856
rect 253498 800 254434 856
rect 254602 800 255630 856
rect 255798 800 256734 856
rect 256902 800 257838 856
rect 258006 800 258942 856
rect 259110 800 260046 856
rect 260214 800 261150 856
rect 261318 800 262346 856
rect 262514 800 263450 856
rect 263618 800 264554 856
rect 264722 800 265658 856
rect 265826 800 266762 856
rect 266930 800 267866 856
rect 268034 800 269062 856
rect 269230 800 270166 856
rect 270334 800 271270 856
rect 271438 800 272374 856
rect 272542 800 273478 856
rect 273646 800 274582 856
rect 274750 800 275778 856
rect 275946 800 276882 856
rect 277050 800 277986 856
rect 278154 800 279090 856
rect 279258 800 280194 856
rect 280362 800 281298 856
rect 281466 800 282494 856
rect 282662 800 283598 856
rect 283766 800 284702 856
rect 284870 800 285806 856
rect 285974 800 286910 856
rect 287078 800 288014 856
rect 288182 800 289118 856
rect 289286 800 290314 856
rect 290482 800 291418 856
rect 291586 800 292522 856
rect 292690 800 293626 856
rect 293794 800 294730 856
rect 294898 800 295834 856
rect 296002 800 297030 856
rect 297198 800 298134 856
rect 298302 800 299238 856
rect 299406 800 300342 856
rect 300510 800 301446 856
rect 301614 800 302550 856
rect 302718 800 303746 856
rect 303914 800 304850 856
rect 305018 800 305954 856
rect 306122 800 307058 856
rect 307226 800 308162 856
rect 308330 800 309266 856
rect 309434 800 310462 856
rect 310630 800 311566 856
rect 311734 800 312670 856
rect 312838 800 313774 856
rect 313942 800 314878 856
rect 315046 800 315982 856
rect 316150 800 317178 856
rect 317346 800 318282 856
rect 318450 800 319386 856
rect 319554 800 320490 856
rect 320658 800 321594 856
rect 321762 800 322698 856
rect 322866 800 323894 856
rect 324062 800 324998 856
rect 325166 800 326102 856
rect 326270 800 327206 856
rect 327374 800 328310 856
rect 328478 800 329414 856
rect 329582 800 330518 856
rect 330686 800 331714 856
rect 331882 800 332818 856
rect 332986 800 333922 856
rect 334090 800 335026 856
rect 335194 800 336130 856
rect 336298 800 337234 856
rect 337402 800 338430 856
rect 338598 800 339534 856
rect 339702 800 340638 856
rect 340806 800 341742 856
rect 341910 800 342846 856
rect 343014 800 343950 856
rect 344118 800 345146 856
rect 345314 800 346250 856
rect 346418 800 347354 856
rect 347522 800 348458 856
rect 348626 800 349562 856
rect 349730 800 350666 856
rect 350834 800 351862 856
rect 352030 800 352966 856
rect 353134 800 354070 856
rect 354238 800 355174 856
rect 355342 800 356278 856
rect 356446 800 357382 856
rect 357550 800 358578 856
rect 358746 800 359682 856
rect 359850 800 360786 856
rect 360954 800 361890 856
rect 362058 800 362994 856
rect 363162 800 364098 856
rect 364266 800 365294 856
rect 365462 800 366398 856
rect 366566 800 367502 856
rect 367670 800 368606 856
rect 368774 800 369710 856
rect 369878 800 370814 856
rect 370982 800 372010 856
rect 372178 800 373114 856
rect 373282 800 374218 856
rect 374386 800 375322 856
rect 375490 800 376426 856
rect 376594 800 377530 856
rect 377698 800 378634 856
rect 378802 800 379830 856
rect 379998 800 380934 856
rect 381102 800 382038 856
rect 382206 800 383142 856
rect 383310 800 384246 856
rect 384414 800 385350 856
rect 385518 800 386546 856
rect 386714 800 387650 856
rect 387818 800 388754 856
rect 388922 800 389858 856
rect 390026 800 390962 856
rect 391130 800 392066 856
rect 392234 800 393262 856
rect 393430 800 394366 856
rect 394534 800 395470 856
rect 395638 800 396574 856
rect 396742 800 397678 856
rect 397846 800 398782 856
rect 398950 800 399978 856
rect 400146 800 401082 856
rect 401250 800 402186 856
rect 402354 800 403290 856
rect 403458 800 404394 856
rect 404562 800 405498 856
rect 405666 800 406694 856
rect 406862 800 407798 856
rect 407966 800 408902 856
rect 409070 800 410006 856
rect 410174 800 411110 856
rect 411278 800 412214 856
rect 412382 800 413410 856
rect 413578 800 414514 856
rect 414682 800 415618 856
rect 415786 800 416722 856
rect 416890 800 417826 856
rect 417994 800 418930 856
rect 419098 800 420126 856
rect 420294 800 421230 856
rect 421398 800 422334 856
rect 422502 800 423438 856
rect 423606 800 424542 856
rect 424710 800 425646 856
rect 425814 800 426750 856
rect 426918 800 427946 856
rect 428114 800 429050 856
rect 429218 800 430154 856
rect 430322 800 431258 856
rect 431426 800 432362 856
rect 432530 800 433466 856
rect 433634 800 434662 856
rect 434830 800 435766 856
rect 435934 800 436870 856
rect 437038 800 437974 856
rect 438142 800 439078 856
rect 439246 800 440182 856
rect 440350 800 441378 856
rect 441546 800 442482 856
rect 442650 800 443586 856
rect 443754 800 444690 856
rect 444858 800 445794 856
rect 445962 800 446898 856
rect 447066 800 448094 856
rect 448262 800 449198 856
rect 449366 800 450302 856
rect 450470 800 451406 856
rect 451574 800 452510 856
rect 452678 800 453614 856
rect 453782 800 454810 856
rect 454978 800 455914 856
rect 456082 800 457018 856
rect 457186 800 458122 856
rect 458290 800 459226 856
rect 459394 800 460330 856
rect 460498 800 461526 856
rect 461694 800 462630 856
rect 462798 800 463734 856
rect 463902 800 464838 856
rect 465006 800 465942 856
rect 466110 800 467046 856
rect 467214 800 468242 856
rect 468410 800 469346 856
rect 469514 800 470450 856
rect 470618 800 471554 856
rect 471722 800 472658 856
rect 472826 800 473762 856
rect 473930 800 474866 856
rect 475034 800 476062 856
rect 476230 800 477166 856
rect 477334 800 478270 856
rect 478438 800 479374 856
rect 479542 800 480478 856
rect 480646 800 481582 856
rect 481750 800 482778 856
rect 482946 800 483882 856
rect 484050 800 484986 856
rect 485154 800 486090 856
rect 486258 800 487194 856
rect 487362 800 488298 856
rect 488466 800 489494 856
rect 489662 800 490598 856
rect 490766 800 491702 856
rect 491870 800 492806 856
rect 492974 800 493910 856
rect 494078 800 495014 856
rect 495182 800 496210 856
rect 496378 800 497314 856
rect 497482 800 498418 856
rect 498586 800 499522 856
rect 499690 800 500626 856
rect 500794 800 501730 856
rect 501898 800 502926 856
rect 503094 800 504030 856
rect 504198 800 505134 856
rect 505302 800 506238 856
rect 506406 800 507342 856
rect 507510 800 508446 856
rect 508614 800 509642 856
rect 509810 800 510746 856
rect 510914 800 511850 856
rect 512018 800 512954 856
rect 513122 800 514058 856
rect 514226 800 515162 856
rect 515330 800 516358 856
rect 516526 800 517462 856
rect 517630 800 518566 856
rect 518734 800 519670 856
rect 519838 800 520774 856
rect 520942 800 521878 856
rect 522046 800 522982 856
rect 523150 800 524178 856
rect 524346 800 525282 856
rect 525450 800 526386 856
rect 526554 800 527490 856
rect 527658 800 528594 856
rect 528762 800 529698 856
rect 529866 800 530894 856
rect 531062 800 531998 856
rect 532166 800 533102 856
rect 533270 800 534206 856
rect 534374 800 535310 856
rect 535478 800 536414 856
rect 536582 800 537610 856
rect 537778 800 538714 856
rect 538882 800 539818 856
rect 539986 800 540922 856
rect 541090 800 542026 856
rect 542194 800 543130 856
rect 543298 800 544326 856
rect 544494 800 545430 856
rect 545598 800 546534 856
rect 546702 800 547638 856
rect 547806 800 548742 856
rect 548910 800 549846 856
rect 550014 800 551042 856
rect 551210 800 552146 856
rect 552314 800 553250 856
rect 553418 800 554354 856
rect 554522 800 555458 856
rect 555626 800 556562 856
rect 556730 800 557476 856
<< metal3 >>
rect 0 626832 800 626952
rect 0 512864 800 512984
rect 0 398896 800 399016
rect 0 284928 800 285048
rect 0 170960 800 171080
rect 0 56992 800 57112
rect 563200 615408 564000 615528
rect 563200 478592 564000 478712
rect 563200 341776 564000 341896
rect 563200 204960 564000 205080
rect 563200 68280 564000 68400
<< obsm3 >>
rect 4208 2143 557488 681665
<< metal4 >>
rect 4208 2128 4528 681680
rect 19568 2128 19888 681680
rect 34928 2128 35248 681680
rect 50288 2128 50608 681680
rect 65648 2128 65968 681680
rect 81008 2128 81328 681680
rect 96368 2128 96688 681680
rect 111728 2128 112048 681680
rect 127088 2128 127408 681680
rect 142448 2128 142768 681680
rect 157808 2128 158128 681680
rect 173168 2128 173488 681680
rect 188528 2128 188848 681680
rect 203888 2128 204208 681680
rect 219248 2128 219568 681680
rect 234608 2128 234928 681680
rect 249968 2128 250288 681680
rect 265328 2128 265648 681680
rect 280688 2128 281008 681680
rect 296048 2128 296368 681680
rect 311408 2128 311728 681680
rect 326768 2128 327088 681680
rect 342128 2128 342448 681680
rect 357488 2128 357808 681680
rect 372848 2128 373168 681680
rect 388208 2128 388528 681680
rect 403568 2128 403888 681680
rect 418928 2128 419248 681680
rect 434288 2128 434608 681680
rect 449648 2128 449968 681680
rect 465008 2128 465328 681680
rect 480368 2128 480688 681680
rect 495728 2128 496048 681680
rect 511088 2128 511408 681680
rect 526448 2128 526768 681680
rect 541808 2128 542128 681680
rect 557168 2128 557488 681680
<< obsm4 >>
rect 18459 3571 19488 677653
rect 19968 3571 34848 677653
rect 35328 3571 50208 677653
rect 50688 3571 65568 677653
rect 66048 3571 80928 677653
rect 81408 3571 96288 677653
rect 96768 3571 111648 677653
rect 112128 3571 127008 677653
rect 127488 3571 142368 677653
rect 142848 3571 157728 677653
rect 158208 3571 173088 677653
rect 173568 3571 188448 677653
rect 188928 3571 203808 677653
rect 204288 3571 219168 677653
rect 219648 3571 234528 677653
rect 235008 3571 249888 677653
rect 250368 3571 265248 677653
rect 265728 3571 280608 677653
rect 281088 3571 295968 677653
rect 296448 3571 311328 677653
rect 311808 3571 326688 677653
rect 327168 3571 342048 677653
rect 342528 3571 357408 677653
rect 357888 3571 372768 677653
rect 373248 3571 388128 677653
rect 388608 3571 403488 677653
rect 403968 3571 418848 677653
rect 419328 3571 434208 677653
rect 434688 3571 449568 677653
rect 450048 3571 464928 677653
rect 465408 3571 480288 677653
rect 480768 3571 495648 677653
rect 496128 3571 511008 677653
rect 511488 3571 526368 677653
rect 526848 3571 533541 677653
<< labels >>
rlabel metal3 s 0 56992 800 57112 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal3 s 0 284928 800 285048 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal3 s 0 398896 800 399016 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal3 s 0 512864 800 512984 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 547602 683200 547658 684000 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 552294 683200 552350 684000 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 554410 0 554466 800 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 556894 683200 556950 684000 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal2 s 555514 0 555570 800 6 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal2 s 556618 0 556674 800 6 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s 563200 204960 564000 205080 6 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 0 170960 800 171080 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal2 s 557814 0 557870 800 6 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal2 s 558918 0 558974 800 6 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal2 s 560022 0 560078 800 6 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal2 s 561586 683200 561642 684000 6 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s 563200 341776 564000 341896 6 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal2 s 561126 0 561182 800 6 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s 0 626832 800 626952 6 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s 563200 478592 564000 478712 6 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal2 s 562230 0 562286 800 6 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 563200 615408 564000 615528 6 analog_io[29]
port 22 nsew signal bidirectional
rlabel metal2 s 549902 0 549958 800 6 analog_io[2]
port 23 nsew signal bidirectional
rlabel metal2 s 563334 0 563390 800 6 analog_io[30]
port 24 nsew signal bidirectional
rlabel metal2 s 533618 683200 533674 684000 6 analog_io[3]
port 25 nsew signal bidirectional
rlabel metal2 s 538310 683200 538366 684000 6 analog_io[4]
port 26 nsew signal bidirectional
rlabel metal3 s 563200 68280 564000 68400 6 analog_io[5]
port 27 nsew signal bidirectional
rlabel metal2 s 551098 0 551154 800 6 analog_io[6]
port 28 nsew signal bidirectional
rlabel metal2 s 552202 0 552258 800 6 analog_io[7]
port 29 nsew signal bidirectional
rlabel metal2 s 553306 0 553362 800 6 analog_io[8]
port 30 nsew signal bidirectional
rlabel metal2 s 542910 683200 542966 684000 6 analog_io[9]
port 31 nsew signal bidirectional
rlabel metal2 s 2318 683200 2374 684000 6 io_in[0]
port 32 nsew signal input
rlabel metal2 s 142066 683200 142122 684000 6 io_in[10]
port 33 nsew signal input
rlabel metal2 s 156050 683200 156106 684000 6 io_in[11]
port 34 nsew signal input
rlabel metal2 s 170034 683200 170090 684000 6 io_in[12]
port 35 nsew signal input
rlabel metal2 s 184018 683200 184074 684000 6 io_in[13]
port 36 nsew signal input
rlabel metal2 s 198002 683200 198058 684000 6 io_in[14]
port 37 nsew signal input
rlabel metal2 s 211986 683200 212042 684000 6 io_in[15]
port 38 nsew signal input
rlabel metal2 s 225970 683200 226026 684000 6 io_in[16]
port 39 nsew signal input
rlabel metal2 s 239954 683200 240010 684000 6 io_in[17]
port 40 nsew signal input
rlabel metal2 s 253938 683200 253994 684000 6 io_in[18]
port 41 nsew signal input
rlabel metal2 s 267922 683200 267978 684000 6 io_in[19]
port 42 nsew signal input
rlabel metal2 s 16210 683200 16266 684000 6 io_in[1]
port 43 nsew signal input
rlabel metal2 s 281906 683200 281962 684000 6 io_in[20]
port 44 nsew signal input
rlabel metal2 s 295890 683200 295946 684000 6 io_in[21]
port 45 nsew signal input
rlabel metal2 s 309874 683200 309930 684000 6 io_in[22]
port 46 nsew signal input
rlabel metal2 s 323858 683200 323914 684000 6 io_in[23]
port 47 nsew signal input
rlabel metal2 s 337842 683200 337898 684000 6 io_in[24]
port 48 nsew signal input
rlabel metal2 s 351826 683200 351882 684000 6 io_in[25]
port 49 nsew signal input
rlabel metal2 s 365810 683200 365866 684000 6 io_in[26]
port 50 nsew signal input
rlabel metal2 s 379794 683200 379850 684000 6 io_in[27]
port 51 nsew signal input
rlabel metal2 s 393778 683200 393834 684000 6 io_in[28]
port 52 nsew signal input
rlabel metal2 s 407762 683200 407818 684000 6 io_in[29]
port 53 nsew signal input
rlabel metal2 s 30194 683200 30250 684000 6 io_in[2]
port 54 nsew signal input
rlabel metal2 s 421746 683200 421802 684000 6 io_in[30]
port 55 nsew signal input
rlabel metal2 s 435730 683200 435786 684000 6 io_in[31]
port 56 nsew signal input
rlabel metal2 s 449714 683200 449770 684000 6 io_in[32]
port 57 nsew signal input
rlabel metal2 s 463698 683200 463754 684000 6 io_in[33]
port 58 nsew signal input
rlabel metal2 s 477682 683200 477738 684000 6 io_in[34]
port 59 nsew signal input
rlabel metal2 s 491666 683200 491722 684000 6 io_in[35]
port 60 nsew signal input
rlabel metal2 s 505650 683200 505706 684000 6 io_in[36]
port 61 nsew signal input
rlabel metal2 s 519634 683200 519690 684000 6 io_in[37]
port 62 nsew signal input
rlabel metal2 s 44178 683200 44234 684000 6 io_in[3]
port 63 nsew signal input
rlabel metal2 s 58162 683200 58218 684000 6 io_in[4]
port 64 nsew signal input
rlabel metal2 s 72146 683200 72202 684000 6 io_in[5]
port 65 nsew signal input
rlabel metal2 s 86130 683200 86186 684000 6 io_in[6]
port 66 nsew signal input
rlabel metal2 s 100114 683200 100170 684000 6 io_in[7]
port 67 nsew signal input
rlabel metal2 s 114098 683200 114154 684000 6 io_in[8]
port 68 nsew signal input
rlabel metal2 s 128082 683200 128138 684000 6 io_in[9]
port 69 nsew signal input
rlabel metal2 s 6918 683200 6974 684000 6 io_oeb[0]
port 70 nsew signal output
rlabel metal2 s 146758 683200 146814 684000 6 io_oeb[10]
port 71 nsew signal output
rlabel metal2 s 160742 683200 160798 684000 6 io_oeb[11]
port 72 nsew signal output
rlabel metal2 s 174726 683200 174782 684000 6 io_oeb[12]
port 73 nsew signal output
rlabel metal2 s 188710 683200 188766 684000 6 io_oeb[13]
port 74 nsew signal output
rlabel metal2 s 202694 683200 202750 684000 6 io_oeb[14]
port 75 nsew signal output
rlabel metal2 s 216678 683200 216734 684000 6 io_oeb[15]
port 76 nsew signal output
rlabel metal2 s 230662 683200 230718 684000 6 io_oeb[16]
port 77 nsew signal output
rlabel metal2 s 244646 683200 244702 684000 6 io_oeb[17]
port 78 nsew signal output
rlabel metal2 s 258630 683200 258686 684000 6 io_oeb[18]
port 79 nsew signal output
rlabel metal2 s 272614 683200 272670 684000 6 io_oeb[19]
port 80 nsew signal output
rlabel metal2 s 20902 683200 20958 684000 6 io_oeb[1]
port 81 nsew signal output
rlabel metal2 s 286598 683200 286654 684000 6 io_oeb[20]
port 82 nsew signal output
rlabel metal2 s 300582 683200 300638 684000 6 io_oeb[21]
port 83 nsew signal output
rlabel metal2 s 314566 683200 314622 684000 6 io_oeb[22]
port 84 nsew signal output
rlabel metal2 s 328550 683200 328606 684000 6 io_oeb[23]
port 85 nsew signal output
rlabel metal2 s 342534 683200 342590 684000 6 io_oeb[24]
port 86 nsew signal output
rlabel metal2 s 356518 683200 356574 684000 6 io_oeb[25]
port 87 nsew signal output
rlabel metal2 s 370502 683200 370558 684000 6 io_oeb[26]
port 88 nsew signal output
rlabel metal2 s 384486 683200 384542 684000 6 io_oeb[27]
port 89 nsew signal output
rlabel metal2 s 398470 683200 398526 684000 6 io_oeb[28]
port 90 nsew signal output
rlabel metal2 s 412454 683200 412510 684000 6 io_oeb[29]
port 91 nsew signal output
rlabel metal2 s 34886 683200 34942 684000 6 io_oeb[2]
port 92 nsew signal output
rlabel metal2 s 426438 683200 426494 684000 6 io_oeb[30]
port 93 nsew signal output
rlabel metal2 s 440422 683200 440478 684000 6 io_oeb[31]
port 94 nsew signal output
rlabel metal2 s 454406 683200 454462 684000 6 io_oeb[32]
port 95 nsew signal output
rlabel metal2 s 468390 683200 468446 684000 6 io_oeb[33]
port 96 nsew signal output
rlabel metal2 s 482374 683200 482430 684000 6 io_oeb[34]
port 97 nsew signal output
rlabel metal2 s 496358 683200 496414 684000 6 io_oeb[35]
port 98 nsew signal output
rlabel metal2 s 510342 683200 510398 684000 6 io_oeb[36]
port 99 nsew signal output
rlabel metal2 s 524326 683200 524382 684000 6 io_oeb[37]
port 100 nsew signal output
rlabel metal2 s 48870 683200 48926 684000 6 io_oeb[3]
port 101 nsew signal output
rlabel metal2 s 62854 683200 62910 684000 6 io_oeb[4]
port 102 nsew signal output
rlabel metal2 s 76838 683200 76894 684000 6 io_oeb[5]
port 103 nsew signal output
rlabel metal2 s 90822 683200 90878 684000 6 io_oeb[6]
port 104 nsew signal output
rlabel metal2 s 104806 683200 104862 684000 6 io_oeb[7]
port 105 nsew signal output
rlabel metal2 s 118790 683200 118846 684000 6 io_oeb[8]
port 106 nsew signal output
rlabel metal2 s 132774 683200 132830 684000 6 io_oeb[9]
port 107 nsew signal output
rlabel metal2 s 11610 683200 11666 684000 6 io_out[0]
port 108 nsew signal output
rlabel metal2 s 151450 683200 151506 684000 6 io_out[10]
port 109 nsew signal output
rlabel metal2 s 165434 683200 165490 684000 6 io_out[11]
port 110 nsew signal output
rlabel metal2 s 179418 683200 179474 684000 6 io_out[12]
port 111 nsew signal output
rlabel metal2 s 193402 683200 193458 684000 6 io_out[13]
port 112 nsew signal output
rlabel metal2 s 207386 683200 207442 684000 6 io_out[14]
port 113 nsew signal output
rlabel metal2 s 221370 683200 221426 684000 6 io_out[15]
port 114 nsew signal output
rlabel metal2 s 235354 683200 235410 684000 6 io_out[16]
port 115 nsew signal output
rlabel metal2 s 249338 683200 249394 684000 6 io_out[17]
port 116 nsew signal output
rlabel metal2 s 263322 683200 263378 684000 6 io_out[18]
port 117 nsew signal output
rlabel metal2 s 277306 683200 277362 684000 6 io_out[19]
port 118 nsew signal output
rlabel metal2 s 25594 683200 25650 684000 6 io_out[1]
port 119 nsew signal output
rlabel metal2 s 291198 683200 291254 684000 6 io_out[20]
port 120 nsew signal output
rlabel metal2 s 305182 683200 305238 684000 6 io_out[21]
port 121 nsew signal output
rlabel metal2 s 319166 683200 319222 684000 6 io_out[22]
port 122 nsew signal output
rlabel metal2 s 333150 683200 333206 684000 6 io_out[23]
port 123 nsew signal output
rlabel metal2 s 347134 683200 347190 684000 6 io_out[24]
port 124 nsew signal output
rlabel metal2 s 361118 683200 361174 684000 6 io_out[25]
port 125 nsew signal output
rlabel metal2 s 375102 683200 375158 684000 6 io_out[26]
port 126 nsew signal output
rlabel metal2 s 389086 683200 389142 684000 6 io_out[27]
port 127 nsew signal output
rlabel metal2 s 403070 683200 403126 684000 6 io_out[28]
port 128 nsew signal output
rlabel metal2 s 417054 683200 417110 684000 6 io_out[29]
port 129 nsew signal output
rlabel metal2 s 39578 683200 39634 684000 6 io_out[2]
port 130 nsew signal output
rlabel metal2 s 431038 683200 431094 684000 6 io_out[30]
port 131 nsew signal output
rlabel metal2 s 445022 683200 445078 684000 6 io_out[31]
port 132 nsew signal output
rlabel metal2 s 459006 683200 459062 684000 6 io_out[32]
port 133 nsew signal output
rlabel metal2 s 472990 683200 473046 684000 6 io_out[33]
port 134 nsew signal output
rlabel metal2 s 486974 683200 487030 684000 6 io_out[34]
port 135 nsew signal output
rlabel metal2 s 500958 683200 501014 684000 6 io_out[35]
port 136 nsew signal output
rlabel metal2 s 514942 683200 514998 684000 6 io_out[36]
port 137 nsew signal output
rlabel metal2 s 528926 683200 528982 684000 6 io_out[37]
port 138 nsew signal output
rlabel metal2 s 53562 683200 53618 684000 6 io_out[3]
port 139 nsew signal output
rlabel metal2 s 67546 683200 67602 684000 6 io_out[4]
port 140 nsew signal output
rlabel metal2 s 81530 683200 81586 684000 6 io_out[5]
port 141 nsew signal output
rlabel metal2 s 95514 683200 95570 684000 6 io_out[6]
port 142 nsew signal output
rlabel metal2 s 109498 683200 109554 684000 6 io_out[7]
port 143 nsew signal output
rlabel metal2 s 123482 683200 123538 684000 6 io_out[8]
port 144 nsew signal output
rlabel metal2 s 137466 683200 137522 684000 6 io_out[9]
port 145 nsew signal output
rlabel metal2 s 119158 0 119214 800 6 la_data_in[0]
port 146 nsew signal input
rlabel metal2 s 454866 0 454922 800 6 la_data_in[100]
port 147 nsew signal input
rlabel metal2 s 458178 0 458234 800 6 la_data_in[101]
port 148 nsew signal input
rlabel metal2 s 461582 0 461638 800 6 la_data_in[102]
port 149 nsew signal input
rlabel metal2 s 464894 0 464950 800 6 la_data_in[103]
port 150 nsew signal input
rlabel metal2 s 468298 0 468354 800 6 la_data_in[104]
port 151 nsew signal input
rlabel metal2 s 471610 0 471666 800 6 la_data_in[105]
port 152 nsew signal input
rlabel metal2 s 474922 0 474978 800 6 la_data_in[106]
port 153 nsew signal input
rlabel metal2 s 478326 0 478382 800 6 la_data_in[107]
port 154 nsew signal input
rlabel metal2 s 481638 0 481694 800 6 la_data_in[108]
port 155 nsew signal input
rlabel metal2 s 485042 0 485098 800 6 la_data_in[109]
port 156 nsew signal input
rlabel metal2 s 152738 0 152794 800 6 la_data_in[10]
port 157 nsew signal input
rlabel metal2 s 488354 0 488410 800 6 la_data_in[110]
port 158 nsew signal input
rlabel metal2 s 491758 0 491814 800 6 la_data_in[111]
port 159 nsew signal input
rlabel metal2 s 495070 0 495126 800 6 la_data_in[112]
port 160 nsew signal input
rlabel metal2 s 498474 0 498530 800 6 la_data_in[113]
port 161 nsew signal input
rlabel metal2 s 501786 0 501842 800 6 la_data_in[114]
port 162 nsew signal input
rlabel metal2 s 505190 0 505246 800 6 la_data_in[115]
port 163 nsew signal input
rlabel metal2 s 508502 0 508558 800 6 la_data_in[116]
port 164 nsew signal input
rlabel metal2 s 511906 0 511962 800 6 la_data_in[117]
port 165 nsew signal input
rlabel metal2 s 515218 0 515274 800 6 la_data_in[118]
port 166 nsew signal input
rlabel metal2 s 518622 0 518678 800 6 la_data_in[119]
port 167 nsew signal input
rlabel metal2 s 156050 0 156106 800 6 la_data_in[11]
port 168 nsew signal input
rlabel metal2 s 521934 0 521990 800 6 la_data_in[120]
port 169 nsew signal input
rlabel metal2 s 525338 0 525394 800 6 la_data_in[121]
port 170 nsew signal input
rlabel metal2 s 528650 0 528706 800 6 la_data_in[122]
port 171 nsew signal input
rlabel metal2 s 532054 0 532110 800 6 la_data_in[123]
port 172 nsew signal input
rlabel metal2 s 535366 0 535422 800 6 la_data_in[124]
port 173 nsew signal input
rlabel metal2 s 538770 0 538826 800 6 la_data_in[125]
port 174 nsew signal input
rlabel metal2 s 542082 0 542138 800 6 la_data_in[126]
port 175 nsew signal input
rlabel metal2 s 545486 0 545542 800 6 la_data_in[127]
port 176 nsew signal input
rlabel metal2 s 159454 0 159510 800 6 la_data_in[12]
port 177 nsew signal input
rlabel metal2 s 162766 0 162822 800 6 la_data_in[13]
port 178 nsew signal input
rlabel metal2 s 166170 0 166226 800 6 la_data_in[14]
port 179 nsew signal input
rlabel metal2 s 169482 0 169538 800 6 la_data_in[15]
port 180 nsew signal input
rlabel metal2 s 172886 0 172942 800 6 la_data_in[16]
port 181 nsew signal input
rlabel metal2 s 176198 0 176254 800 6 la_data_in[17]
port 182 nsew signal input
rlabel metal2 s 179602 0 179658 800 6 la_data_in[18]
port 183 nsew signal input
rlabel metal2 s 182914 0 182970 800 6 la_data_in[19]
port 184 nsew signal input
rlabel metal2 s 122470 0 122526 800 6 la_data_in[1]
port 185 nsew signal input
rlabel metal2 s 186318 0 186374 800 6 la_data_in[20]
port 186 nsew signal input
rlabel metal2 s 189630 0 189686 800 6 la_data_in[21]
port 187 nsew signal input
rlabel metal2 s 192942 0 192998 800 6 la_data_in[22]
port 188 nsew signal input
rlabel metal2 s 196346 0 196402 800 6 la_data_in[23]
port 189 nsew signal input
rlabel metal2 s 199658 0 199714 800 6 la_data_in[24]
port 190 nsew signal input
rlabel metal2 s 203062 0 203118 800 6 la_data_in[25]
port 191 nsew signal input
rlabel metal2 s 206374 0 206430 800 6 la_data_in[26]
port 192 nsew signal input
rlabel metal2 s 209778 0 209834 800 6 la_data_in[27]
port 193 nsew signal input
rlabel metal2 s 213090 0 213146 800 6 la_data_in[28]
port 194 nsew signal input
rlabel metal2 s 216494 0 216550 800 6 la_data_in[29]
port 195 nsew signal input
rlabel metal2 s 125874 0 125930 800 6 la_data_in[2]
port 196 nsew signal input
rlabel metal2 s 219806 0 219862 800 6 la_data_in[30]
port 197 nsew signal input
rlabel metal2 s 223210 0 223266 800 6 la_data_in[31]
port 198 nsew signal input
rlabel metal2 s 226522 0 226578 800 6 la_data_in[32]
port 199 nsew signal input
rlabel metal2 s 229926 0 229982 800 6 la_data_in[33]
port 200 nsew signal input
rlabel metal2 s 233238 0 233294 800 6 la_data_in[34]
port 201 nsew signal input
rlabel metal2 s 236642 0 236698 800 6 la_data_in[35]
port 202 nsew signal input
rlabel metal2 s 239954 0 240010 800 6 la_data_in[36]
port 203 nsew signal input
rlabel metal2 s 243358 0 243414 800 6 la_data_in[37]
port 204 nsew signal input
rlabel metal2 s 246670 0 246726 800 6 la_data_in[38]
port 205 nsew signal input
rlabel metal2 s 250074 0 250130 800 6 la_data_in[39]
port 206 nsew signal input
rlabel metal2 s 129186 0 129242 800 6 la_data_in[3]
port 207 nsew signal input
rlabel metal2 s 253386 0 253442 800 6 la_data_in[40]
port 208 nsew signal input
rlabel metal2 s 256790 0 256846 800 6 la_data_in[41]
port 209 nsew signal input
rlabel metal2 s 260102 0 260158 800 6 la_data_in[42]
port 210 nsew signal input
rlabel metal2 s 263506 0 263562 800 6 la_data_in[43]
port 211 nsew signal input
rlabel metal2 s 266818 0 266874 800 6 la_data_in[44]
port 212 nsew signal input
rlabel metal2 s 270222 0 270278 800 6 la_data_in[45]
port 213 nsew signal input
rlabel metal2 s 273534 0 273590 800 6 la_data_in[46]
port 214 nsew signal input
rlabel metal2 s 276938 0 276994 800 6 la_data_in[47]
port 215 nsew signal input
rlabel metal2 s 280250 0 280306 800 6 la_data_in[48]
port 216 nsew signal input
rlabel metal2 s 283654 0 283710 800 6 la_data_in[49]
port 217 nsew signal input
rlabel metal2 s 132590 0 132646 800 6 la_data_in[4]
port 218 nsew signal input
rlabel metal2 s 286966 0 287022 800 6 la_data_in[50]
port 219 nsew signal input
rlabel metal2 s 290370 0 290426 800 6 la_data_in[51]
port 220 nsew signal input
rlabel metal2 s 293682 0 293738 800 6 la_data_in[52]
port 221 nsew signal input
rlabel metal2 s 297086 0 297142 800 6 la_data_in[53]
port 222 nsew signal input
rlabel metal2 s 300398 0 300454 800 6 la_data_in[54]
port 223 nsew signal input
rlabel metal2 s 303802 0 303858 800 6 la_data_in[55]
port 224 nsew signal input
rlabel metal2 s 307114 0 307170 800 6 la_data_in[56]
port 225 nsew signal input
rlabel metal2 s 310518 0 310574 800 6 la_data_in[57]
port 226 nsew signal input
rlabel metal2 s 313830 0 313886 800 6 la_data_in[58]
port 227 nsew signal input
rlabel metal2 s 317234 0 317290 800 6 la_data_in[59]
port 228 nsew signal input
rlabel metal2 s 135902 0 135958 800 6 la_data_in[5]
port 229 nsew signal input
rlabel metal2 s 320546 0 320602 800 6 la_data_in[60]
port 230 nsew signal input
rlabel metal2 s 323950 0 324006 800 6 la_data_in[61]
port 231 nsew signal input
rlabel metal2 s 327262 0 327318 800 6 la_data_in[62]
port 232 nsew signal input
rlabel metal2 s 330574 0 330630 800 6 la_data_in[63]
port 233 nsew signal input
rlabel metal2 s 333978 0 334034 800 6 la_data_in[64]
port 234 nsew signal input
rlabel metal2 s 337290 0 337346 800 6 la_data_in[65]
port 235 nsew signal input
rlabel metal2 s 340694 0 340750 800 6 la_data_in[66]
port 236 nsew signal input
rlabel metal2 s 344006 0 344062 800 6 la_data_in[67]
port 237 nsew signal input
rlabel metal2 s 347410 0 347466 800 6 la_data_in[68]
port 238 nsew signal input
rlabel metal2 s 350722 0 350778 800 6 la_data_in[69]
port 239 nsew signal input
rlabel metal2 s 139306 0 139362 800 6 la_data_in[6]
port 240 nsew signal input
rlabel metal2 s 354126 0 354182 800 6 la_data_in[70]
port 241 nsew signal input
rlabel metal2 s 357438 0 357494 800 6 la_data_in[71]
port 242 nsew signal input
rlabel metal2 s 360842 0 360898 800 6 la_data_in[72]
port 243 nsew signal input
rlabel metal2 s 364154 0 364210 800 6 la_data_in[73]
port 244 nsew signal input
rlabel metal2 s 367558 0 367614 800 6 la_data_in[74]
port 245 nsew signal input
rlabel metal2 s 370870 0 370926 800 6 la_data_in[75]
port 246 nsew signal input
rlabel metal2 s 374274 0 374330 800 6 la_data_in[76]
port 247 nsew signal input
rlabel metal2 s 377586 0 377642 800 6 la_data_in[77]
port 248 nsew signal input
rlabel metal2 s 380990 0 381046 800 6 la_data_in[78]
port 249 nsew signal input
rlabel metal2 s 384302 0 384358 800 6 la_data_in[79]
port 250 nsew signal input
rlabel metal2 s 142618 0 142674 800 6 la_data_in[7]
port 251 nsew signal input
rlabel metal2 s 387706 0 387762 800 6 la_data_in[80]
port 252 nsew signal input
rlabel metal2 s 391018 0 391074 800 6 la_data_in[81]
port 253 nsew signal input
rlabel metal2 s 394422 0 394478 800 6 la_data_in[82]
port 254 nsew signal input
rlabel metal2 s 397734 0 397790 800 6 la_data_in[83]
port 255 nsew signal input
rlabel metal2 s 401138 0 401194 800 6 la_data_in[84]
port 256 nsew signal input
rlabel metal2 s 404450 0 404506 800 6 la_data_in[85]
port 257 nsew signal input
rlabel metal2 s 407854 0 407910 800 6 la_data_in[86]
port 258 nsew signal input
rlabel metal2 s 411166 0 411222 800 6 la_data_in[87]
port 259 nsew signal input
rlabel metal2 s 414570 0 414626 800 6 la_data_in[88]
port 260 nsew signal input
rlabel metal2 s 417882 0 417938 800 6 la_data_in[89]
port 261 nsew signal input
rlabel metal2 s 146022 0 146078 800 6 la_data_in[8]
port 262 nsew signal input
rlabel metal2 s 421286 0 421342 800 6 la_data_in[90]
port 263 nsew signal input
rlabel metal2 s 424598 0 424654 800 6 la_data_in[91]
port 264 nsew signal input
rlabel metal2 s 428002 0 428058 800 6 la_data_in[92]
port 265 nsew signal input
rlabel metal2 s 431314 0 431370 800 6 la_data_in[93]
port 266 nsew signal input
rlabel metal2 s 434718 0 434774 800 6 la_data_in[94]
port 267 nsew signal input
rlabel metal2 s 438030 0 438086 800 6 la_data_in[95]
port 268 nsew signal input
rlabel metal2 s 441434 0 441490 800 6 la_data_in[96]
port 269 nsew signal input
rlabel metal2 s 444746 0 444802 800 6 la_data_in[97]
port 270 nsew signal input
rlabel metal2 s 448150 0 448206 800 6 la_data_in[98]
port 271 nsew signal input
rlabel metal2 s 451462 0 451518 800 6 la_data_in[99]
port 272 nsew signal input
rlabel metal2 s 149334 0 149390 800 6 la_data_in[9]
port 273 nsew signal input
rlabel metal2 s 120262 0 120318 800 6 la_data_out[0]
port 274 nsew signal output
rlabel metal2 s 455970 0 456026 800 6 la_data_out[100]
port 275 nsew signal output
rlabel metal2 s 459282 0 459338 800 6 la_data_out[101]
port 276 nsew signal output
rlabel metal2 s 462686 0 462742 800 6 la_data_out[102]
port 277 nsew signal output
rlabel metal2 s 465998 0 466054 800 6 la_data_out[103]
port 278 nsew signal output
rlabel metal2 s 469402 0 469458 800 6 la_data_out[104]
port 279 nsew signal output
rlabel metal2 s 472714 0 472770 800 6 la_data_out[105]
port 280 nsew signal output
rlabel metal2 s 476118 0 476174 800 6 la_data_out[106]
port 281 nsew signal output
rlabel metal2 s 479430 0 479486 800 6 la_data_out[107]
port 282 nsew signal output
rlabel metal2 s 482834 0 482890 800 6 la_data_out[108]
port 283 nsew signal output
rlabel metal2 s 486146 0 486202 800 6 la_data_out[109]
port 284 nsew signal output
rlabel metal2 s 153842 0 153898 800 6 la_data_out[10]
port 285 nsew signal output
rlabel metal2 s 489550 0 489606 800 6 la_data_out[110]
port 286 nsew signal output
rlabel metal2 s 492862 0 492918 800 6 la_data_out[111]
port 287 nsew signal output
rlabel metal2 s 496266 0 496322 800 6 la_data_out[112]
port 288 nsew signal output
rlabel metal2 s 499578 0 499634 800 6 la_data_out[113]
port 289 nsew signal output
rlabel metal2 s 502982 0 503038 800 6 la_data_out[114]
port 290 nsew signal output
rlabel metal2 s 506294 0 506350 800 6 la_data_out[115]
port 291 nsew signal output
rlabel metal2 s 509698 0 509754 800 6 la_data_out[116]
port 292 nsew signal output
rlabel metal2 s 513010 0 513066 800 6 la_data_out[117]
port 293 nsew signal output
rlabel metal2 s 516414 0 516470 800 6 la_data_out[118]
port 294 nsew signal output
rlabel metal2 s 519726 0 519782 800 6 la_data_out[119]
port 295 nsew signal output
rlabel metal2 s 157154 0 157210 800 6 la_data_out[11]
port 296 nsew signal output
rlabel metal2 s 523038 0 523094 800 6 la_data_out[120]
port 297 nsew signal output
rlabel metal2 s 526442 0 526498 800 6 la_data_out[121]
port 298 nsew signal output
rlabel metal2 s 529754 0 529810 800 6 la_data_out[122]
port 299 nsew signal output
rlabel metal2 s 533158 0 533214 800 6 la_data_out[123]
port 300 nsew signal output
rlabel metal2 s 536470 0 536526 800 6 la_data_out[124]
port 301 nsew signal output
rlabel metal2 s 539874 0 539930 800 6 la_data_out[125]
port 302 nsew signal output
rlabel metal2 s 543186 0 543242 800 6 la_data_out[126]
port 303 nsew signal output
rlabel metal2 s 546590 0 546646 800 6 la_data_out[127]
port 304 nsew signal output
rlabel metal2 s 160558 0 160614 800 6 la_data_out[12]
port 305 nsew signal output
rlabel metal2 s 163870 0 163926 800 6 la_data_out[13]
port 306 nsew signal output
rlabel metal2 s 167274 0 167330 800 6 la_data_out[14]
port 307 nsew signal output
rlabel metal2 s 170586 0 170642 800 6 la_data_out[15]
port 308 nsew signal output
rlabel metal2 s 173990 0 174046 800 6 la_data_out[16]
port 309 nsew signal output
rlabel metal2 s 177302 0 177358 800 6 la_data_out[17]
port 310 nsew signal output
rlabel metal2 s 180706 0 180762 800 6 la_data_out[18]
port 311 nsew signal output
rlabel metal2 s 184018 0 184074 800 6 la_data_out[19]
port 312 nsew signal output
rlabel metal2 s 123574 0 123630 800 6 la_data_out[1]
port 313 nsew signal output
rlabel metal2 s 187422 0 187478 800 6 la_data_out[20]
port 314 nsew signal output
rlabel metal2 s 190734 0 190790 800 6 la_data_out[21]
port 315 nsew signal output
rlabel metal2 s 194138 0 194194 800 6 la_data_out[22]
port 316 nsew signal output
rlabel metal2 s 197450 0 197506 800 6 la_data_out[23]
port 317 nsew signal output
rlabel metal2 s 200854 0 200910 800 6 la_data_out[24]
port 318 nsew signal output
rlabel metal2 s 204166 0 204222 800 6 la_data_out[25]
port 319 nsew signal output
rlabel metal2 s 207570 0 207626 800 6 la_data_out[26]
port 320 nsew signal output
rlabel metal2 s 210882 0 210938 800 6 la_data_out[27]
port 321 nsew signal output
rlabel metal2 s 214286 0 214342 800 6 la_data_out[28]
port 322 nsew signal output
rlabel metal2 s 217598 0 217654 800 6 la_data_out[29]
port 323 nsew signal output
rlabel metal2 s 126978 0 127034 800 6 la_data_out[2]
port 324 nsew signal output
rlabel metal2 s 221002 0 221058 800 6 la_data_out[30]
port 325 nsew signal output
rlabel metal2 s 224314 0 224370 800 6 la_data_out[31]
port 326 nsew signal output
rlabel metal2 s 227718 0 227774 800 6 la_data_out[32]
port 327 nsew signal output
rlabel metal2 s 231030 0 231086 800 6 la_data_out[33]
port 328 nsew signal output
rlabel metal2 s 234434 0 234490 800 6 la_data_out[34]
port 329 nsew signal output
rlabel metal2 s 237746 0 237802 800 6 la_data_out[35]
port 330 nsew signal output
rlabel metal2 s 241058 0 241114 800 6 la_data_out[36]
port 331 nsew signal output
rlabel metal2 s 244462 0 244518 800 6 la_data_out[37]
port 332 nsew signal output
rlabel metal2 s 247774 0 247830 800 6 la_data_out[38]
port 333 nsew signal output
rlabel metal2 s 251178 0 251234 800 6 la_data_out[39]
port 334 nsew signal output
rlabel metal2 s 130290 0 130346 800 6 la_data_out[3]
port 335 nsew signal output
rlabel metal2 s 254490 0 254546 800 6 la_data_out[40]
port 336 nsew signal output
rlabel metal2 s 257894 0 257950 800 6 la_data_out[41]
port 337 nsew signal output
rlabel metal2 s 261206 0 261262 800 6 la_data_out[42]
port 338 nsew signal output
rlabel metal2 s 264610 0 264666 800 6 la_data_out[43]
port 339 nsew signal output
rlabel metal2 s 267922 0 267978 800 6 la_data_out[44]
port 340 nsew signal output
rlabel metal2 s 271326 0 271382 800 6 la_data_out[45]
port 341 nsew signal output
rlabel metal2 s 274638 0 274694 800 6 la_data_out[46]
port 342 nsew signal output
rlabel metal2 s 278042 0 278098 800 6 la_data_out[47]
port 343 nsew signal output
rlabel metal2 s 281354 0 281410 800 6 la_data_out[48]
port 344 nsew signal output
rlabel metal2 s 284758 0 284814 800 6 la_data_out[49]
port 345 nsew signal output
rlabel metal2 s 133694 0 133750 800 6 la_data_out[4]
port 346 nsew signal output
rlabel metal2 s 288070 0 288126 800 6 la_data_out[50]
port 347 nsew signal output
rlabel metal2 s 291474 0 291530 800 6 la_data_out[51]
port 348 nsew signal output
rlabel metal2 s 294786 0 294842 800 6 la_data_out[52]
port 349 nsew signal output
rlabel metal2 s 298190 0 298246 800 6 la_data_out[53]
port 350 nsew signal output
rlabel metal2 s 301502 0 301558 800 6 la_data_out[54]
port 351 nsew signal output
rlabel metal2 s 304906 0 304962 800 6 la_data_out[55]
port 352 nsew signal output
rlabel metal2 s 308218 0 308274 800 6 la_data_out[56]
port 353 nsew signal output
rlabel metal2 s 311622 0 311678 800 6 la_data_out[57]
port 354 nsew signal output
rlabel metal2 s 314934 0 314990 800 6 la_data_out[58]
port 355 nsew signal output
rlabel metal2 s 318338 0 318394 800 6 la_data_out[59]
port 356 nsew signal output
rlabel metal2 s 137006 0 137062 800 6 la_data_out[5]
port 357 nsew signal output
rlabel metal2 s 321650 0 321706 800 6 la_data_out[60]
port 358 nsew signal output
rlabel metal2 s 325054 0 325110 800 6 la_data_out[61]
port 359 nsew signal output
rlabel metal2 s 328366 0 328422 800 6 la_data_out[62]
port 360 nsew signal output
rlabel metal2 s 331770 0 331826 800 6 la_data_out[63]
port 361 nsew signal output
rlabel metal2 s 335082 0 335138 800 6 la_data_out[64]
port 362 nsew signal output
rlabel metal2 s 338486 0 338542 800 6 la_data_out[65]
port 363 nsew signal output
rlabel metal2 s 341798 0 341854 800 6 la_data_out[66]
port 364 nsew signal output
rlabel metal2 s 345202 0 345258 800 6 la_data_out[67]
port 365 nsew signal output
rlabel metal2 s 348514 0 348570 800 6 la_data_out[68]
port 366 nsew signal output
rlabel metal2 s 351918 0 351974 800 6 la_data_out[69]
port 367 nsew signal output
rlabel metal2 s 140410 0 140466 800 6 la_data_out[6]
port 368 nsew signal output
rlabel metal2 s 355230 0 355286 800 6 la_data_out[70]
port 369 nsew signal output
rlabel metal2 s 358634 0 358690 800 6 la_data_out[71]
port 370 nsew signal output
rlabel metal2 s 361946 0 362002 800 6 la_data_out[72]
port 371 nsew signal output
rlabel metal2 s 365350 0 365406 800 6 la_data_out[73]
port 372 nsew signal output
rlabel metal2 s 368662 0 368718 800 6 la_data_out[74]
port 373 nsew signal output
rlabel metal2 s 372066 0 372122 800 6 la_data_out[75]
port 374 nsew signal output
rlabel metal2 s 375378 0 375434 800 6 la_data_out[76]
port 375 nsew signal output
rlabel metal2 s 378690 0 378746 800 6 la_data_out[77]
port 376 nsew signal output
rlabel metal2 s 382094 0 382150 800 6 la_data_out[78]
port 377 nsew signal output
rlabel metal2 s 385406 0 385462 800 6 la_data_out[79]
port 378 nsew signal output
rlabel metal2 s 143722 0 143778 800 6 la_data_out[7]
port 379 nsew signal output
rlabel metal2 s 388810 0 388866 800 6 la_data_out[80]
port 380 nsew signal output
rlabel metal2 s 392122 0 392178 800 6 la_data_out[81]
port 381 nsew signal output
rlabel metal2 s 395526 0 395582 800 6 la_data_out[82]
port 382 nsew signal output
rlabel metal2 s 398838 0 398894 800 6 la_data_out[83]
port 383 nsew signal output
rlabel metal2 s 402242 0 402298 800 6 la_data_out[84]
port 384 nsew signal output
rlabel metal2 s 405554 0 405610 800 6 la_data_out[85]
port 385 nsew signal output
rlabel metal2 s 408958 0 409014 800 6 la_data_out[86]
port 386 nsew signal output
rlabel metal2 s 412270 0 412326 800 6 la_data_out[87]
port 387 nsew signal output
rlabel metal2 s 415674 0 415730 800 6 la_data_out[88]
port 388 nsew signal output
rlabel metal2 s 418986 0 419042 800 6 la_data_out[89]
port 389 nsew signal output
rlabel metal2 s 147126 0 147182 800 6 la_data_out[8]
port 390 nsew signal output
rlabel metal2 s 422390 0 422446 800 6 la_data_out[90]
port 391 nsew signal output
rlabel metal2 s 425702 0 425758 800 6 la_data_out[91]
port 392 nsew signal output
rlabel metal2 s 429106 0 429162 800 6 la_data_out[92]
port 393 nsew signal output
rlabel metal2 s 432418 0 432474 800 6 la_data_out[93]
port 394 nsew signal output
rlabel metal2 s 435822 0 435878 800 6 la_data_out[94]
port 395 nsew signal output
rlabel metal2 s 439134 0 439190 800 6 la_data_out[95]
port 396 nsew signal output
rlabel metal2 s 442538 0 442594 800 6 la_data_out[96]
port 397 nsew signal output
rlabel metal2 s 445850 0 445906 800 6 la_data_out[97]
port 398 nsew signal output
rlabel metal2 s 449254 0 449310 800 6 la_data_out[98]
port 399 nsew signal output
rlabel metal2 s 452566 0 452622 800 6 la_data_out[99]
port 400 nsew signal output
rlabel metal2 s 150438 0 150494 800 6 la_data_out[9]
port 401 nsew signal output
rlabel metal2 s 121366 0 121422 800 6 la_oen[0]
port 402 nsew signal input
rlabel metal2 s 457074 0 457130 800 6 la_oen[100]
port 403 nsew signal input
rlabel metal2 s 460386 0 460442 800 6 la_oen[101]
port 404 nsew signal input
rlabel metal2 s 463790 0 463846 800 6 la_oen[102]
port 405 nsew signal input
rlabel metal2 s 467102 0 467158 800 6 la_oen[103]
port 406 nsew signal input
rlabel metal2 s 470506 0 470562 800 6 la_oen[104]
port 407 nsew signal input
rlabel metal2 s 473818 0 473874 800 6 la_oen[105]
port 408 nsew signal input
rlabel metal2 s 477222 0 477278 800 6 la_oen[106]
port 409 nsew signal input
rlabel metal2 s 480534 0 480590 800 6 la_oen[107]
port 410 nsew signal input
rlabel metal2 s 483938 0 483994 800 6 la_oen[108]
port 411 nsew signal input
rlabel metal2 s 487250 0 487306 800 6 la_oen[109]
port 412 nsew signal input
rlabel metal2 s 154946 0 155002 800 6 la_oen[10]
port 413 nsew signal input
rlabel metal2 s 490654 0 490710 800 6 la_oen[110]
port 414 nsew signal input
rlabel metal2 s 493966 0 494022 800 6 la_oen[111]
port 415 nsew signal input
rlabel metal2 s 497370 0 497426 800 6 la_oen[112]
port 416 nsew signal input
rlabel metal2 s 500682 0 500738 800 6 la_oen[113]
port 417 nsew signal input
rlabel metal2 s 504086 0 504142 800 6 la_oen[114]
port 418 nsew signal input
rlabel metal2 s 507398 0 507454 800 6 la_oen[115]
port 419 nsew signal input
rlabel metal2 s 510802 0 510858 800 6 la_oen[116]
port 420 nsew signal input
rlabel metal2 s 514114 0 514170 800 6 la_oen[117]
port 421 nsew signal input
rlabel metal2 s 517518 0 517574 800 6 la_oen[118]
port 422 nsew signal input
rlabel metal2 s 520830 0 520886 800 6 la_oen[119]
port 423 nsew signal input
rlabel metal2 s 158258 0 158314 800 6 la_oen[11]
port 424 nsew signal input
rlabel metal2 s 524234 0 524290 800 6 la_oen[120]
port 425 nsew signal input
rlabel metal2 s 527546 0 527602 800 6 la_oen[121]
port 426 nsew signal input
rlabel metal2 s 530950 0 531006 800 6 la_oen[122]
port 427 nsew signal input
rlabel metal2 s 534262 0 534318 800 6 la_oen[123]
port 428 nsew signal input
rlabel metal2 s 537666 0 537722 800 6 la_oen[124]
port 429 nsew signal input
rlabel metal2 s 540978 0 541034 800 6 la_oen[125]
port 430 nsew signal input
rlabel metal2 s 544382 0 544438 800 6 la_oen[126]
port 431 nsew signal input
rlabel metal2 s 547694 0 547750 800 6 la_oen[127]
port 432 nsew signal input
rlabel metal2 s 161662 0 161718 800 6 la_oen[12]
port 433 nsew signal input
rlabel metal2 s 164974 0 165030 800 6 la_oen[13]
port 434 nsew signal input
rlabel metal2 s 168378 0 168434 800 6 la_oen[14]
port 435 nsew signal input
rlabel metal2 s 171690 0 171746 800 6 la_oen[15]
port 436 nsew signal input
rlabel metal2 s 175094 0 175150 800 6 la_oen[16]
port 437 nsew signal input
rlabel metal2 s 178406 0 178462 800 6 la_oen[17]
port 438 nsew signal input
rlabel metal2 s 181810 0 181866 800 6 la_oen[18]
port 439 nsew signal input
rlabel metal2 s 185122 0 185178 800 6 la_oen[19]
port 440 nsew signal input
rlabel metal2 s 124770 0 124826 800 6 la_oen[1]
port 441 nsew signal input
rlabel metal2 s 188526 0 188582 800 6 la_oen[20]
port 442 nsew signal input
rlabel metal2 s 191838 0 191894 800 6 la_oen[21]
port 443 nsew signal input
rlabel metal2 s 195242 0 195298 800 6 la_oen[22]
port 444 nsew signal input
rlabel metal2 s 198554 0 198610 800 6 la_oen[23]
port 445 nsew signal input
rlabel metal2 s 201958 0 202014 800 6 la_oen[24]
port 446 nsew signal input
rlabel metal2 s 205270 0 205326 800 6 la_oen[25]
port 447 nsew signal input
rlabel metal2 s 208674 0 208730 800 6 la_oen[26]
port 448 nsew signal input
rlabel metal2 s 211986 0 212042 800 6 la_oen[27]
port 449 nsew signal input
rlabel metal2 s 215390 0 215446 800 6 la_oen[28]
port 450 nsew signal input
rlabel metal2 s 218702 0 218758 800 6 la_oen[29]
port 451 nsew signal input
rlabel metal2 s 128082 0 128138 800 6 la_oen[2]
port 452 nsew signal input
rlabel metal2 s 222106 0 222162 800 6 la_oen[30]
port 453 nsew signal input
rlabel metal2 s 225418 0 225474 800 6 la_oen[31]
port 454 nsew signal input
rlabel metal2 s 228822 0 228878 800 6 la_oen[32]
port 455 nsew signal input
rlabel metal2 s 232134 0 232190 800 6 la_oen[33]
port 456 nsew signal input
rlabel metal2 s 235538 0 235594 800 6 la_oen[34]
port 457 nsew signal input
rlabel metal2 s 238850 0 238906 800 6 la_oen[35]
port 458 nsew signal input
rlabel metal2 s 242254 0 242310 800 6 la_oen[36]
port 459 nsew signal input
rlabel metal2 s 245566 0 245622 800 6 la_oen[37]
port 460 nsew signal input
rlabel metal2 s 248970 0 249026 800 6 la_oen[38]
port 461 nsew signal input
rlabel metal2 s 252282 0 252338 800 6 la_oen[39]
port 462 nsew signal input
rlabel metal2 s 131486 0 131542 800 6 la_oen[3]
port 463 nsew signal input
rlabel metal2 s 255686 0 255742 800 6 la_oen[40]
port 464 nsew signal input
rlabel metal2 s 258998 0 259054 800 6 la_oen[41]
port 465 nsew signal input
rlabel metal2 s 262402 0 262458 800 6 la_oen[42]
port 466 nsew signal input
rlabel metal2 s 265714 0 265770 800 6 la_oen[43]
port 467 nsew signal input
rlabel metal2 s 269118 0 269174 800 6 la_oen[44]
port 468 nsew signal input
rlabel metal2 s 272430 0 272486 800 6 la_oen[45]
port 469 nsew signal input
rlabel metal2 s 275834 0 275890 800 6 la_oen[46]
port 470 nsew signal input
rlabel metal2 s 279146 0 279202 800 6 la_oen[47]
port 471 nsew signal input
rlabel metal2 s 282550 0 282606 800 6 la_oen[48]
port 472 nsew signal input
rlabel metal2 s 285862 0 285918 800 6 la_oen[49]
port 473 nsew signal input
rlabel metal2 s 134798 0 134854 800 6 la_oen[4]
port 474 nsew signal input
rlabel metal2 s 289174 0 289230 800 6 la_oen[50]
port 475 nsew signal input
rlabel metal2 s 292578 0 292634 800 6 la_oen[51]
port 476 nsew signal input
rlabel metal2 s 295890 0 295946 800 6 la_oen[52]
port 477 nsew signal input
rlabel metal2 s 299294 0 299350 800 6 la_oen[53]
port 478 nsew signal input
rlabel metal2 s 302606 0 302662 800 6 la_oen[54]
port 479 nsew signal input
rlabel metal2 s 306010 0 306066 800 6 la_oen[55]
port 480 nsew signal input
rlabel metal2 s 309322 0 309378 800 6 la_oen[56]
port 481 nsew signal input
rlabel metal2 s 312726 0 312782 800 6 la_oen[57]
port 482 nsew signal input
rlabel metal2 s 316038 0 316094 800 6 la_oen[58]
port 483 nsew signal input
rlabel metal2 s 319442 0 319498 800 6 la_oen[59]
port 484 nsew signal input
rlabel metal2 s 138202 0 138258 800 6 la_oen[5]
port 485 nsew signal input
rlabel metal2 s 322754 0 322810 800 6 la_oen[60]
port 486 nsew signal input
rlabel metal2 s 326158 0 326214 800 6 la_oen[61]
port 487 nsew signal input
rlabel metal2 s 329470 0 329526 800 6 la_oen[62]
port 488 nsew signal input
rlabel metal2 s 332874 0 332930 800 6 la_oen[63]
port 489 nsew signal input
rlabel metal2 s 336186 0 336242 800 6 la_oen[64]
port 490 nsew signal input
rlabel metal2 s 339590 0 339646 800 6 la_oen[65]
port 491 nsew signal input
rlabel metal2 s 342902 0 342958 800 6 la_oen[66]
port 492 nsew signal input
rlabel metal2 s 346306 0 346362 800 6 la_oen[67]
port 493 nsew signal input
rlabel metal2 s 349618 0 349674 800 6 la_oen[68]
port 494 nsew signal input
rlabel metal2 s 353022 0 353078 800 6 la_oen[69]
port 495 nsew signal input
rlabel metal2 s 141514 0 141570 800 6 la_oen[6]
port 496 nsew signal input
rlabel metal2 s 356334 0 356390 800 6 la_oen[70]
port 497 nsew signal input
rlabel metal2 s 359738 0 359794 800 6 la_oen[71]
port 498 nsew signal input
rlabel metal2 s 363050 0 363106 800 6 la_oen[72]
port 499 nsew signal input
rlabel metal2 s 366454 0 366510 800 6 la_oen[73]
port 500 nsew signal input
rlabel metal2 s 369766 0 369822 800 6 la_oen[74]
port 501 nsew signal input
rlabel metal2 s 373170 0 373226 800 6 la_oen[75]
port 502 nsew signal input
rlabel metal2 s 376482 0 376538 800 6 la_oen[76]
port 503 nsew signal input
rlabel metal2 s 379886 0 379942 800 6 la_oen[77]
port 504 nsew signal input
rlabel metal2 s 383198 0 383254 800 6 la_oen[78]
port 505 nsew signal input
rlabel metal2 s 386602 0 386658 800 6 la_oen[79]
port 506 nsew signal input
rlabel metal2 s 144826 0 144882 800 6 la_oen[7]
port 507 nsew signal input
rlabel metal2 s 389914 0 389970 800 6 la_oen[80]
port 508 nsew signal input
rlabel metal2 s 393318 0 393374 800 6 la_oen[81]
port 509 nsew signal input
rlabel metal2 s 396630 0 396686 800 6 la_oen[82]
port 510 nsew signal input
rlabel metal2 s 400034 0 400090 800 6 la_oen[83]
port 511 nsew signal input
rlabel metal2 s 403346 0 403402 800 6 la_oen[84]
port 512 nsew signal input
rlabel metal2 s 406750 0 406806 800 6 la_oen[85]
port 513 nsew signal input
rlabel metal2 s 410062 0 410118 800 6 la_oen[86]
port 514 nsew signal input
rlabel metal2 s 413466 0 413522 800 6 la_oen[87]
port 515 nsew signal input
rlabel metal2 s 416778 0 416834 800 6 la_oen[88]
port 516 nsew signal input
rlabel metal2 s 420182 0 420238 800 6 la_oen[89]
port 517 nsew signal input
rlabel metal2 s 148230 0 148286 800 6 la_oen[8]
port 518 nsew signal input
rlabel metal2 s 423494 0 423550 800 6 la_oen[90]
port 519 nsew signal input
rlabel metal2 s 426806 0 426862 800 6 la_oen[91]
port 520 nsew signal input
rlabel metal2 s 430210 0 430266 800 6 la_oen[92]
port 521 nsew signal input
rlabel metal2 s 433522 0 433578 800 6 la_oen[93]
port 522 nsew signal input
rlabel metal2 s 436926 0 436982 800 6 la_oen[94]
port 523 nsew signal input
rlabel metal2 s 440238 0 440294 800 6 la_oen[95]
port 524 nsew signal input
rlabel metal2 s 443642 0 443698 800 6 la_oen[96]
port 525 nsew signal input
rlabel metal2 s 446954 0 447010 800 6 la_oen[97]
port 526 nsew signal input
rlabel metal2 s 450358 0 450414 800 6 la_oen[98]
port 527 nsew signal input
rlabel metal2 s 453670 0 453726 800 6 la_oen[99]
port 528 nsew signal input
rlabel metal2 s 151542 0 151598 800 6 la_oen[9]
port 529 nsew signal input
rlabel metal2 s 548798 0 548854 800 6 user_clock2
port 530 nsew signal input
rlabel metal2 s 570 0 626 800 6 wb_clk_i
port 531 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wb_rst_i
port 532 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 wbs_ack_o
port 533 nsew signal output
rlabel metal2 s 7194 0 7250 800 6 wbs_adr_i[0]
port 534 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 wbs_adr_i[10]
port 535 nsew signal input
rlabel metal2 s 48594 0 48650 800 6 wbs_adr_i[11]
port 536 nsew signal input
rlabel metal2 s 51998 0 52054 800 6 wbs_adr_i[12]
port 537 nsew signal input
rlabel metal2 s 55310 0 55366 800 6 wbs_adr_i[13]
port 538 nsew signal input
rlabel metal2 s 58714 0 58770 800 6 wbs_adr_i[14]
port 539 nsew signal input
rlabel metal2 s 62026 0 62082 800 6 wbs_adr_i[15]
port 540 nsew signal input
rlabel metal2 s 65430 0 65486 800 6 wbs_adr_i[16]
port 541 nsew signal input
rlabel metal2 s 68742 0 68798 800 6 wbs_adr_i[17]
port 542 nsew signal input
rlabel metal2 s 72146 0 72202 800 6 wbs_adr_i[18]
port 543 nsew signal input
rlabel metal2 s 75458 0 75514 800 6 wbs_adr_i[19]
port 544 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 wbs_adr_i[1]
port 545 nsew signal input
rlabel metal2 s 78862 0 78918 800 6 wbs_adr_i[20]
port 546 nsew signal input
rlabel metal2 s 82174 0 82230 800 6 wbs_adr_i[21]
port 547 nsew signal input
rlabel metal2 s 85578 0 85634 800 6 wbs_adr_i[22]
port 548 nsew signal input
rlabel metal2 s 88890 0 88946 800 6 wbs_adr_i[23]
port 549 nsew signal input
rlabel metal2 s 92294 0 92350 800 6 wbs_adr_i[24]
port 550 nsew signal input
rlabel metal2 s 95606 0 95662 800 6 wbs_adr_i[25]
port 551 nsew signal input
rlabel metal2 s 99010 0 99066 800 6 wbs_adr_i[26]
port 552 nsew signal input
rlabel metal2 s 102322 0 102378 800 6 wbs_adr_i[27]
port 553 nsew signal input
rlabel metal2 s 105726 0 105782 800 6 wbs_adr_i[28]
port 554 nsew signal input
rlabel metal2 s 109038 0 109094 800 6 wbs_adr_i[29]
port 555 nsew signal input
rlabel metal2 s 16210 0 16266 800 6 wbs_adr_i[2]
port 556 nsew signal input
rlabel metal2 s 112442 0 112498 800 6 wbs_adr_i[30]
port 557 nsew signal input
rlabel metal2 s 115754 0 115810 800 6 wbs_adr_i[31]
port 558 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 wbs_adr_i[3]
port 559 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 wbs_adr_i[4]
port 560 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 wbs_adr_i[5]
port 561 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 wbs_adr_i[6]
port 562 nsew signal input
rlabel metal2 s 35254 0 35310 800 6 wbs_adr_i[7]
port 563 nsew signal input
rlabel metal2 s 38566 0 38622 800 6 wbs_adr_i[8]
port 564 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 wbs_adr_i[9]
port 565 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 wbs_cyc_i
port 566 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 wbs_dat_i[0]
port 567 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 wbs_dat_i[10]
port 568 nsew signal input
rlabel metal2 s 49790 0 49846 800 6 wbs_dat_i[11]
port 569 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 wbs_dat_i[12]
port 570 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 wbs_dat_i[13]
port 571 nsew signal input
rlabel metal2 s 59818 0 59874 800 6 wbs_dat_i[14]
port 572 nsew signal input
rlabel metal2 s 63222 0 63278 800 6 wbs_dat_i[15]
port 573 nsew signal input
rlabel metal2 s 66534 0 66590 800 6 wbs_dat_i[16]
port 574 nsew signal input
rlabel metal2 s 69938 0 69994 800 6 wbs_dat_i[17]
port 575 nsew signal input
rlabel metal2 s 73250 0 73306 800 6 wbs_dat_i[18]
port 576 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 wbs_dat_i[19]
port 577 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 wbs_dat_i[1]
port 578 nsew signal input
rlabel metal2 s 79966 0 80022 800 6 wbs_dat_i[20]
port 579 nsew signal input
rlabel metal2 s 83370 0 83426 800 6 wbs_dat_i[21]
port 580 nsew signal input
rlabel metal2 s 86682 0 86738 800 6 wbs_dat_i[22]
port 581 nsew signal input
rlabel metal2 s 90086 0 90142 800 6 wbs_dat_i[23]
port 582 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 wbs_dat_i[24]
port 583 nsew signal input
rlabel metal2 s 96710 0 96766 800 6 wbs_dat_i[25]
port 584 nsew signal input
rlabel metal2 s 100114 0 100170 800 6 wbs_dat_i[26]
port 585 nsew signal input
rlabel metal2 s 103426 0 103482 800 6 wbs_dat_i[27]
port 586 nsew signal input
rlabel metal2 s 106830 0 106886 800 6 wbs_dat_i[28]
port 587 nsew signal input
rlabel metal2 s 110142 0 110198 800 6 wbs_dat_i[29]
port 588 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 wbs_dat_i[2]
port 589 nsew signal input
rlabel metal2 s 113546 0 113602 800 6 wbs_dat_i[30]
port 590 nsew signal input
rlabel metal2 s 116858 0 116914 800 6 wbs_dat_i[31]
port 591 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 wbs_dat_i[3]
port 592 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 wbs_dat_i[4]
port 593 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 wbs_dat_i[5]
port 594 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 wbs_dat_i[6]
port 595 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 wbs_dat_i[7]
port 596 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 wbs_dat_i[8]
port 597 nsew signal input
rlabel metal2 s 43074 0 43130 800 6 wbs_dat_i[9]
port 598 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 wbs_dat_o[0]
port 599 nsew signal output
rlabel metal2 s 47490 0 47546 800 6 wbs_dat_o[10]
port 600 nsew signal output
rlabel metal2 s 50894 0 50950 800 6 wbs_dat_o[11]
port 601 nsew signal output
rlabel metal2 s 54206 0 54262 800 6 wbs_dat_o[12]
port 602 nsew signal output
rlabel metal2 s 57610 0 57666 800 6 wbs_dat_o[13]
port 603 nsew signal output
rlabel metal2 s 60922 0 60978 800 6 wbs_dat_o[14]
port 604 nsew signal output
rlabel metal2 s 64326 0 64382 800 6 wbs_dat_o[15]
port 605 nsew signal output
rlabel metal2 s 67638 0 67694 800 6 wbs_dat_o[16]
port 606 nsew signal output
rlabel metal2 s 71042 0 71098 800 6 wbs_dat_o[17]
port 607 nsew signal output
rlabel metal2 s 74354 0 74410 800 6 wbs_dat_o[18]
port 608 nsew signal output
rlabel metal2 s 77758 0 77814 800 6 wbs_dat_o[19]
port 609 nsew signal output
rlabel metal2 s 13910 0 13966 800 6 wbs_dat_o[1]
port 610 nsew signal output
rlabel metal2 s 81070 0 81126 800 6 wbs_dat_o[20]
port 611 nsew signal output
rlabel metal2 s 84474 0 84530 800 6 wbs_dat_o[21]
port 612 nsew signal output
rlabel metal2 s 87786 0 87842 800 6 wbs_dat_o[22]
port 613 nsew signal output
rlabel metal2 s 91190 0 91246 800 6 wbs_dat_o[23]
port 614 nsew signal output
rlabel metal2 s 94502 0 94558 800 6 wbs_dat_o[24]
port 615 nsew signal output
rlabel metal2 s 97906 0 97962 800 6 wbs_dat_o[25]
port 616 nsew signal output
rlabel metal2 s 101218 0 101274 800 6 wbs_dat_o[26]
port 617 nsew signal output
rlabel metal2 s 104622 0 104678 800 6 wbs_dat_o[27]
port 618 nsew signal output
rlabel metal2 s 107934 0 107990 800 6 wbs_dat_o[28]
port 619 nsew signal output
rlabel metal2 s 111338 0 111394 800 6 wbs_dat_o[29]
port 620 nsew signal output
rlabel metal2 s 18418 0 18474 800 6 wbs_dat_o[2]
port 621 nsew signal output
rlabel metal2 s 114650 0 114706 800 6 wbs_dat_o[30]
port 622 nsew signal output
rlabel metal2 s 118054 0 118110 800 6 wbs_dat_o[31]
port 623 nsew signal output
rlabel metal2 s 22926 0 22982 800 6 wbs_dat_o[3]
port 624 nsew signal output
rlabel metal2 s 27342 0 27398 800 6 wbs_dat_o[4]
port 625 nsew signal output
rlabel metal2 s 30746 0 30802 800 6 wbs_dat_o[5]
port 626 nsew signal output
rlabel metal2 s 34058 0 34114 800 6 wbs_dat_o[6]
port 627 nsew signal output
rlabel metal2 s 37462 0 37518 800 6 wbs_dat_o[7]
port 628 nsew signal output
rlabel metal2 s 40774 0 40830 800 6 wbs_dat_o[8]
port 629 nsew signal output
rlabel metal2 s 44178 0 44234 800 6 wbs_dat_o[9]
port 630 nsew signal output
rlabel metal2 s 10598 0 10654 800 6 wbs_sel_i[0]
port 631 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 wbs_sel_i[1]
port 632 nsew signal input
rlabel metal2 s 19522 0 19578 800 6 wbs_sel_i[2]
port 633 nsew signal input
rlabel metal2 s 24030 0 24086 800 6 wbs_sel_i[3]
port 634 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 wbs_stb_i
port 635 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 wbs_we_i
port 636 nsew signal input
rlabel metal4 s 557168 2128 557488 681680 6 VPWR
port 637 nsew power bidirectional
rlabel metal4 s 526448 2128 526768 681680 6 VPWR
port 638 nsew power bidirectional
rlabel metal4 s 495728 2128 496048 681680 6 VPWR
port 639 nsew power bidirectional
rlabel metal4 s 465008 2128 465328 681680 6 VPWR
port 640 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 681680 6 VPWR
port 641 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 681680 6 VPWR
port 642 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 681680 6 VPWR
port 643 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 681680 6 VPWR
port 644 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 681680 6 VPWR
port 645 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 681680 6 VPWR
port 646 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 681680 6 VPWR
port 647 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 681680 6 VPWR
port 648 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 681680 6 VPWR
port 649 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 681680 6 VPWR
port 650 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 681680 6 VPWR
port 651 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 681680 6 VPWR
port 652 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 681680 6 VPWR
port 653 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 681680 6 VPWR
port 654 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 681680 6 VPWR
port 655 nsew power bidirectional
rlabel metal4 s 541808 2128 542128 681680 6 VGND
port 656 nsew ground bidirectional
rlabel metal4 s 511088 2128 511408 681680 6 VGND
port 657 nsew ground bidirectional
rlabel metal4 s 480368 2128 480688 681680 6 VGND
port 658 nsew ground bidirectional
rlabel metal4 s 449648 2128 449968 681680 6 VGND
port 659 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 681680 6 VGND
port 660 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 681680 6 VGND
port 661 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 681680 6 VGND
port 662 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 681680 6 VGND
port 663 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 681680 6 VGND
port 664 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 681680 6 VGND
port 665 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 681680 6 VGND
port 666 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 681680 6 VGND
port 667 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 681680 6 VGND
port 668 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 681680 6 VGND
port 669 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 681680 6 VGND
port 670 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 681680 6 VGND
port 671 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 681680 6 VGND
port 672 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 681680 6 VGND
port 673 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 564000 684000
string LEFview TRUE
<< end >>

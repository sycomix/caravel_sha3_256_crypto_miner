magic
tech sky130A
magscale 1 2
timestamp 1608366604
<< obsli1 >>
rect 1104 2159 562856 681649
<< obsm1 >>
rect 566 1844 562856 681680
<< metal2 >>
rect 2226 683200 2282 684000
rect 6642 683200 6698 684000
rect 11058 683200 11114 684000
rect 15474 683200 15530 684000
rect 19982 683200 20038 684000
rect 24398 683200 24454 684000
rect 28814 683200 28870 684000
rect 33230 683200 33286 684000
rect 37738 683200 37794 684000
rect 42154 683200 42210 684000
rect 46570 683200 46626 684000
rect 50986 683200 51042 684000
rect 55494 683200 55550 684000
rect 59910 683200 59966 684000
rect 64326 683200 64382 684000
rect 68834 683200 68890 684000
rect 73250 683200 73306 684000
rect 77666 683200 77722 684000
rect 82082 683200 82138 684000
rect 86590 683200 86646 684000
rect 91006 683200 91062 684000
rect 95422 683200 95478 684000
rect 99838 683200 99894 684000
rect 104346 683200 104402 684000
rect 108762 683200 108818 684000
rect 113178 683200 113234 684000
rect 117594 683200 117650 684000
rect 122102 683200 122158 684000
rect 126518 683200 126574 684000
rect 130934 683200 130990 684000
rect 135442 683200 135498 684000
rect 139858 683200 139914 684000
rect 144274 683200 144330 684000
rect 148690 683200 148746 684000
rect 153198 683200 153254 684000
rect 157614 683200 157670 684000
rect 162030 683200 162086 684000
rect 166446 683200 166502 684000
rect 170954 683200 171010 684000
rect 175370 683200 175426 684000
rect 179786 683200 179842 684000
rect 184202 683200 184258 684000
rect 188710 683200 188766 684000
rect 193126 683200 193182 684000
rect 197542 683200 197598 684000
rect 202050 683200 202106 684000
rect 206466 683200 206522 684000
rect 210882 683200 210938 684000
rect 215298 683200 215354 684000
rect 219806 683200 219862 684000
rect 224222 683200 224278 684000
rect 228638 683200 228694 684000
rect 233054 683200 233110 684000
rect 237562 683200 237618 684000
rect 241978 683200 242034 684000
rect 246394 683200 246450 684000
rect 250810 683200 250866 684000
rect 255318 683200 255374 684000
rect 259734 683200 259790 684000
rect 264150 683200 264206 684000
rect 268658 683200 268714 684000
rect 273074 683200 273130 684000
rect 277490 683200 277546 684000
rect 281906 683200 281962 684000
rect 286414 683200 286470 684000
rect 290830 683200 290886 684000
rect 295246 683200 295302 684000
rect 299662 683200 299718 684000
rect 304170 683200 304226 684000
rect 308586 683200 308642 684000
rect 313002 683200 313058 684000
rect 317510 683200 317566 684000
rect 321926 683200 321982 684000
rect 326342 683200 326398 684000
rect 330758 683200 330814 684000
rect 335266 683200 335322 684000
rect 339682 683200 339738 684000
rect 344098 683200 344154 684000
rect 348514 683200 348570 684000
rect 353022 683200 353078 684000
rect 357438 683200 357494 684000
rect 361854 683200 361910 684000
rect 366270 683200 366326 684000
rect 370778 683200 370834 684000
rect 375194 683200 375250 684000
rect 379610 683200 379666 684000
rect 384118 683200 384174 684000
rect 388534 683200 388590 684000
rect 392950 683200 393006 684000
rect 397366 683200 397422 684000
rect 401874 683200 401930 684000
rect 406290 683200 406346 684000
rect 410706 683200 410762 684000
rect 415122 683200 415178 684000
rect 419630 683200 419686 684000
rect 424046 683200 424102 684000
rect 428462 683200 428518 684000
rect 432878 683200 432934 684000
rect 437386 683200 437442 684000
rect 441802 683200 441858 684000
rect 446218 683200 446274 684000
rect 450726 683200 450782 684000
rect 455142 683200 455198 684000
rect 459558 683200 459614 684000
rect 463974 683200 464030 684000
rect 468482 683200 468538 684000
rect 472898 683200 472954 684000
rect 477314 683200 477370 684000
rect 481730 683200 481786 684000
rect 486238 683200 486294 684000
rect 490654 683200 490710 684000
rect 495070 683200 495126 684000
rect 499486 683200 499542 684000
rect 503994 683200 504050 684000
rect 508410 683200 508466 684000
rect 512826 683200 512882 684000
rect 517334 683200 517390 684000
rect 521750 683200 521806 684000
rect 526166 683200 526222 684000
rect 530582 683200 530638 684000
rect 535090 683200 535146 684000
rect 539506 683200 539562 684000
rect 543922 683200 543978 684000
rect 548338 683200 548394 684000
rect 552846 683200 552902 684000
rect 557262 683200 557318 684000
rect 561678 683200 561734 684000
rect 570 0 626 800
rect 1674 0 1730 800
rect 2778 0 2834 800
rect 3974 0 4030 800
rect 5078 0 5134 800
rect 6182 0 6238 800
rect 7378 0 7434 800
rect 8482 0 8538 800
rect 9586 0 9642 800
rect 10782 0 10838 800
rect 11886 0 11942 800
rect 12990 0 13046 800
rect 14186 0 14242 800
rect 15290 0 15346 800
rect 16394 0 16450 800
rect 17590 0 17646 800
rect 18694 0 18750 800
rect 19798 0 19854 800
rect 20994 0 21050 800
rect 22098 0 22154 800
rect 23202 0 23258 800
rect 24398 0 24454 800
rect 25502 0 25558 800
rect 26606 0 26662 800
rect 27802 0 27858 800
rect 28906 0 28962 800
rect 30010 0 30066 800
rect 31206 0 31262 800
rect 32310 0 32366 800
rect 33414 0 33470 800
rect 34610 0 34666 800
rect 35714 0 35770 800
rect 36818 0 36874 800
rect 38014 0 38070 800
rect 39118 0 39174 800
rect 40222 0 40278 800
rect 41418 0 41474 800
rect 42522 0 42578 800
rect 43626 0 43682 800
rect 44822 0 44878 800
rect 45926 0 45982 800
rect 47030 0 47086 800
rect 48226 0 48282 800
rect 49330 0 49386 800
rect 50434 0 50490 800
rect 51630 0 51686 800
rect 52734 0 52790 800
rect 53838 0 53894 800
rect 55034 0 55090 800
rect 56138 0 56194 800
rect 57242 0 57298 800
rect 58438 0 58494 800
rect 59542 0 59598 800
rect 60646 0 60702 800
rect 61842 0 61898 800
rect 62946 0 63002 800
rect 64050 0 64106 800
rect 65246 0 65302 800
rect 66350 0 66406 800
rect 67454 0 67510 800
rect 68650 0 68706 800
rect 69754 0 69810 800
rect 70858 0 70914 800
rect 72054 0 72110 800
rect 73158 0 73214 800
rect 74262 0 74318 800
rect 75458 0 75514 800
rect 76562 0 76618 800
rect 77666 0 77722 800
rect 78862 0 78918 800
rect 79966 0 80022 800
rect 81070 0 81126 800
rect 82266 0 82322 800
rect 83370 0 83426 800
rect 84474 0 84530 800
rect 85670 0 85726 800
rect 86774 0 86830 800
rect 87878 0 87934 800
rect 89074 0 89130 800
rect 90178 0 90234 800
rect 91282 0 91338 800
rect 92478 0 92534 800
rect 93582 0 93638 800
rect 94686 0 94742 800
rect 95882 0 95938 800
rect 96986 0 97042 800
rect 98090 0 98146 800
rect 99286 0 99342 800
rect 100390 0 100446 800
rect 101494 0 101550 800
rect 102690 0 102746 800
rect 103794 0 103850 800
rect 104898 0 104954 800
rect 106094 0 106150 800
rect 107198 0 107254 800
rect 108302 0 108358 800
rect 109498 0 109554 800
rect 110602 0 110658 800
rect 111706 0 111762 800
rect 112902 0 112958 800
rect 114006 0 114062 800
rect 115110 0 115166 800
rect 116306 0 116362 800
rect 117410 0 117466 800
rect 118514 0 118570 800
rect 119710 0 119766 800
rect 120814 0 120870 800
rect 121918 0 121974 800
rect 123114 0 123170 800
rect 124218 0 124274 800
rect 125322 0 125378 800
rect 126518 0 126574 800
rect 127622 0 127678 800
rect 128726 0 128782 800
rect 129922 0 129978 800
rect 131026 0 131082 800
rect 132130 0 132186 800
rect 133326 0 133382 800
rect 134430 0 134486 800
rect 135534 0 135590 800
rect 136730 0 136786 800
rect 137834 0 137890 800
rect 138938 0 138994 800
rect 140134 0 140190 800
rect 141238 0 141294 800
rect 142342 0 142398 800
rect 143538 0 143594 800
rect 144642 0 144698 800
rect 145746 0 145802 800
rect 146942 0 146998 800
rect 148046 0 148102 800
rect 149150 0 149206 800
rect 150346 0 150402 800
rect 151450 0 151506 800
rect 152554 0 152610 800
rect 153750 0 153806 800
rect 154854 0 154910 800
rect 155958 0 156014 800
rect 157154 0 157210 800
rect 158258 0 158314 800
rect 159362 0 159418 800
rect 160558 0 160614 800
rect 161662 0 161718 800
rect 162766 0 162822 800
rect 163962 0 164018 800
rect 165066 0 165122 800
rect 166170 0 166226 800
rect 167366 0 167422 800
rect 168470 0 168526 800
rect 169574 0 169630 800
rect 170770 0 170826 800
rect 171874 0 171930 800
rect 172978 0 173034 800
rect 174174 0 174230 800
rect 175278 0 175334 800
rect 176382 0 176438 800
rect 177578 0 177634 800
rect 178682 0 178738 800
rect 179786 0 179842 800
rect 180982 0 181038 800
rect 182086 0 182142 800
rect 183190 0 183246 800
rect 184386 0 184442 800
rect 185490 0 185546 800
rect 186594 0 186650 800
rect 187790 0 187846 800
rect 188894 0 188950 800
rect 189998 0 190054 800
rect 191194 0 191250 800
rect 192298 0 192354 800
rect 193402 0 193458 800
rect 194598 0 194654 800
rect 195702 0 195758 800
rect 196806 0 196862 800
rect 198002 0 198058 800
rect 199106 0 199162 800
rect 200210 0 200266 800
rect 201406 0 201462 800
rect 202510 0 202566 800
rect 203614 0 203670 800
rect 204810 0 204866 800
rect 205914 0 205970 800
rect 207018 0 207074 800
rect 208214 0 208270 800
rect 209318 0 209374 800
rect 210422 0 210478 800
rect 211618 0 211674 800
rect 212722 0 212778 800
rect 213826 0 213882 800
rect 215022 0 215078 800
rect 216126 0 216182 800
rect 217230 0 217286 800
rect 218426 0 218482 800
rect 219530 0 219586 800
rect 220634 0 220690 800
rect 221830 0 221886 800
rect 222934 0 222990 800
rect 224038 0 224094 800
rect 225234 0 225290 800
rect 226338 0 226394 800
rect 227442 0 227498 800
rect 228638 0 228694 800
rect 229742 0 229798 800
rect 230846 0 230902 800
rect 232042 0 232098 800
rect 233146 0 233202 800
rect 234250 0 234306 800
rect 235446 0 235502 800
rect 236550 0 236606 800
rect 237654 0 237710 800
rect 238850 0 238906 800
rect 239954 0 240010 800
rect 241058 0 241114 800
rect 242254 0 242310 800
rect 243358 0 243414 800
rect 244462 0 244518 800
rect 245658 0 245714 800
rect 246762 0 246818 800
rect 247866 0 247922 800
rect 249062 0 249118 800
rect 250166 0 250222 800
rect 251270 0 251326 800
rect 252466 0 252522 800
rect 253570 0 253626 800
rect 254674 0 254730 800
rect 255870 0 255926 800
rect 256974 0 257030 800
rect 258078 0 258134 800
rect 259274 0 259330 800
rect 260378 0 260434 800
rect 261482 0 261538 800
rect 262678 0 262734 800
rect 263782 0 263838 800
rect 264886 0 264942 800
rect 266082 0 266138 800
rect 267186 0 267242 800
rect 268290 0 268346 800
rect 269486 0 269542 800
rect 270590 0 270646 800
rect 271694 0 271750 800
rect 272890 0 272946 800
rect 273994 0 274050 800
rect 275098 0 275154 800
rect 276294 0 276350 800
rect 277398 0 277454 800
rect 278502 0 278558 800
rect 279698 0 279754 800
rect 280802 0 280858 800
rect 281906 0 281962 800
rect 283102 0 283158 800
rect 284206 0 284262 800
rect 285310 0 285366 800
rect 286506 0 286562 800
rect 287610 0 287666 800
rect 288714 0 288770 800
rect 289910 0 289966 800
rect 291014 0 291070 800
rect 292118 0 292174 800
rect 293314 0 293370 800
rect 294418 0 294474 800
rect 295522 0 295578 800
rect 296718 0 296774 800
rect 297822 0 297878 800
rect 298926 0 298982 800
rect 300122 0 300178 800
rect 301226 0 301282 800
rect 302330 0 302386 800
rect 303526 0 303582 800
rect 304630 0 304686 800
rect 305734 0 305790 800
rect 306930 0 306986 800
rect 308034 0 308090 800
rect 309138 0 309194 800
rect 310334 0 310390 800
rect 311438 0 311494 800
rect 312542 0 312598 800
rect 313738 0 313794 800
rect 314842 0 314898 800
rect 315946 0 316002 800
rect 317142 0 317198 800
rect 318246 0 318302 800
rect 319350 0 319406 800
rect 320546 0 320602 800
rect 321650 0 321706 800
rect 322754 0 322810 800
rect 323950 0 324006 800
rect 325054 0 325110 800
rect 326158 0 326214 800
rect 327354 0 327410 800
rect 328458 0 328514 800
rect 329562 0 329618 800
rect 330758 0 330814 800
rect 331862 0 331918 800
rect 332966 0 333022 800
rect 334162 0 334218 800
rect 335266 0 335322 800
rect 336370 0 336426 800
rect 337566 0 337622 800
rect 338670 0 338726 800
rect 339774 0 339830 800
rect 340970 0 341026 800
rect 342074 0 342130 800
rect 343178 0 343234 800
rect 344374 0 344430 800
rect 345478 0 345534 800
rect 346582 0 346638 800
rect 347778 0 347834 800
rect 348882 0 348938 800
rect 349986 0 350042 800
rect 351182 0 351238 800
rect 352286 0 352342 800
rect 353390 0 353446 800
rect 354586 0 354642 800
rect 355690 0 355746 800
rect 356794 0 356850 800
rect 357990 0 358046 800
rect 359094 0 359150 800
rect 360198 0 360254 800
rect 361394 0 361450 800
rect 362498 0 362554 800
rect 363602 0 363658 800
rect 364798 0 364854 800
rect 365902 0 365958 800
rect 367006 0 367062 800
rect 368202 0 368258 800
rect 369306 0 369362 800
rect 370410 0 370466 800
rect 371606 0 371662 800
rect 372710 0 372766 800
rect 373814 0 373870 800
rect 375010 0 375066 800
rect 376114 0 376170 800
rect 377218 0 377274 800
rect 378414 0 378470 800
rect 379518 0 379574 800
rect 380622 0 380678 800
rect 381818 0 381874 800
rect 382922 0 382978 800
rect 384026 0 384082 800
rect 385222 0 385278 800
rect 386326 0 386382 800
rect 387430 0 387486 800
rect 388626 0 388682 800
rect 389730 0 389786 800
rect 390834 0 390890 800
rect 392030 0 392086 800
rect 393134 0 393190 800
rect 394238 0 394294 800
rect 395434 0 395490 800
rect 396538 0 396594 800
rect 397642 0 397698 800
rect 398838 0 398894 800
rect 399942 0 399998 800
rect 401046 0 401102 800
rect 402242 0 402298 800
rect 403346 0 403402 800
rect 404450 0 404506 800
rect 405646 0 405702 800
rect 406750 0 406806 800
rect 407854 0 407910 800
rect 409050 0 409106 800
rect 410154 0 410210 800
rect 411258 0 411314 800
rect 412454 0 412510 800
rect 413558 0 413614 800
rect 414662 0 414718 800
rect 415858 0 415914 800
rect 416962 0 417018 800
rect 418066 0 418122 800
rect 419262 0 419318 800
rect 420366 0 420422 800
rect 421470 0 421526 800
rect 422666 0 422722 800
rect 423770 0 423826 800
rect 424874 0 424930 800
rect 426070 0 426126 800
rect 427174 0 427230 800
rect 428278 0 428334 800
rect 429474 0 429530 800
rect 430578 0 430634 800
rect 431682 0 431738 800
rect 432878 0 432934 800
rect 433982 0 434038 800
rect 435086 0 435142 800
rect 436282 0 436338 800
rect 437386 0 437442 800
rect 438490 0 438546 800
rect 439686 0 439742 800
rect 440790 0 440846 800
rect 441894 0 441950 800
rect 443090 0 443146 800
rect 444194 0 444250 800
rect 445298 0 445354 800
rect 446494 0 446550 800
rect 447598 0 447654 800
rect 448702 0 448758 800
rect 449898 0 449954 800
rect 451002 0 451058 800
rect 452106 0 452162 800
rect 453302 0 453358 800
rect 454406 0 454462 800
rect 455510 0 455566 800
rect 456706 0 456762 800
rect 457810 0 457866 800
rect 458914 0 458970 800
rect 460110 0 460166 800
rect 461214 0 461270 800
rect 462318 0 462374 800
rect 463514 0 463570 800
rect 464618 0 464674 800
rect 465722 0 465778 800
rect 466918 0 466974 800
rect 468022 0 468078 800
rect 469126 0 469182 800
rect 470322 0 470378 800
rect 471426 0 471482 800
rect 472530 0 472586 800
rect 473726 0 473782 800
rect 474830 0 474886 800
rect 475934 0 475990 800
rect 477130 0 477186 800
rect 478234 0 478290 800
rect 479338 0 479394 800
rect 480534 0 480590 800
rect 481638 0 481694 800
rect 482742 0 482798 800
rect 483938 0 483994 800
rect 485042 0 485098 800
rect 486146 0 486202 800
rect 487342 0 487398 800
rect 488446 0 488502 800
rect 489550 0 489606 800
rect 490746 0 490802 800
rect 491850 0 491906 800
rect 492954 0 493010 800
rect 494150 0 494206 800
rect 495254 0 495310 800
rect 496358 0 496414 800
rect 497554 0 497610 800
rect 498658 0 498714 800
rect 499762 0 499818 800
rect 500958 0 501014 800
rect 502062 0 502118 800
rect 503166 0 503222 800
rect 504362 0 504418 800
rect 505466 0 505522 800
rect 506570 0 506626 800
rect 507766 0 507822 800
rect 508870 0 508926 800
rect 509974 0 510030 800
rect 511170 0 511226 800
rect 512274 0 512330 800
rect 513378 0 513434 800
rect 514574 0 514630 800
rect 515678 0 515734 800
rect 516782 0 516838 800
rect 517978 0 518034 800
rect 519082 0 519138 800
rect 520186 0 520242 800
rect 521382 0 521438 800
rect 522486 0 522542 800
rect 523590 0 523646 800
rect 524786 0 524842 800
rect 525890 0 525946 800
rect 526994 0 527050 800
rect 528190 0 528246 800
rect 529294 0 529350 800
rect 530398 0 530454 800
rect 531594 0 531650 800
rect 532698 0 532754 800
rect 533802 0 533858 800
rect 534998 0 535054 800
rect 536102 0 536158 800
rect 537206 0 537262 800
rect 538402 0 538458 800
rect 539506 0 539562 800
rect 540610 0 540666 800
rect 541806 0 541862 800
rect 542910 0 542966 800
rect 544014 0 544070 800
rect 545210 0 545266 800
rect 546314 0 546370 800
rect 547418 0 547474 800
rect 548614 0 548670 800
rect 549718 0 549774 800
rect 550822 0 550878 800
rect 552018 0 552074 800
rect 553122 0 553178 800
rect 554226 0 554282 800
rect 555422 0 555478 800
rect 556526 0 556582 800
rect 557630 0 557686 800
rect 558826 0 558882 800
rect 559930 0 559986 800
rect 561034 0 561090 800
rect 562230 0 562286 800
rect 563334 0 563390 800
<< obsm2 >>
rect 572 683144 2170 683200
rect 2338 683144 6586 683200
rect 6754 683144 11002 683200
rect 11170 683144 15418 683200
rect 15586 683144 19926 683200
rect 20094 683144 24342 683200
rect 24510 683144 28758 683200
rect 28926 683144 33174 683200
rect 33342 683144 37682 683200
rect 37850 683144 42098 683200
rect 42266 683144 46514 683200
rect 46682 683144 50930 683200
rect 51098 683144 55438 683200
rect 55606 683144 59854 683200
rect 60022 683144 64270 683200
rect 64438 683144 68778 683200
rect 68946 683144 73194 683200
rect 73362 683144 77610 683200
rect 77778 683144 82026 683200
rect 82194 683144 86534 683200
rect 86702 683144 90950 683200
rect 91118 683144 95366 683200
rect 95534 683144 99782 683200
rect 99950 683144 104290 683200
rect 104458 683144 108706 683200
rect 108874 683144 113122 683200
rect 113290 683144 117538 683200
rect 117706 683144 122046 683200
rect 122214 683144 126462 683200
rect 126630 683144 130878 683200
rect 131046 683144 135386 683200
rect 135554 683144 139802 683200
rect 139970 683144 144218 683200
rect 144386 683144 148634 683200
rect 148802 683144 153142 683200
rect 153310 683144 157558 683200
rect 157726 683144 161974 683200
rect 162142 683144 166390 683200
rect 166558 683144 170898 683200
rect 171066 683144 175314 683200
rect 175482 683144 179730 683200
rect 179898 683144 184146 683200
rect 184314 683144 188654 683200
rect 188822 683144 193070 683200
rect 193238 683144 197486 683200
rect 197654 683144 201994 683200
rect 202162 683144 206410 683200
rect 206578 683144 210826 683200
rect 210994 683144 215242 683200
rect 215410 683144 219750 683200
rect 219918 683144 224166 683200
rect 224334 683144 228582 683200
rect 228750 683144 232998 683200
rect 233166 683144 237506 683200
rect 237674 683144 241922 683200
rect 242090 683144 246338 683200
rect 246506 683144 250754 683200
rect 250922 683144 255262 683200
rect 255430 683144 259678 683200
rect 259846 683144 264094 683200
rect 264262 683144 268602 683200
rect 268770 683144 273018 683200
rect 273186 683144 277434 683200
rect 277602 683144 281850 683200
rect 282018 683144 286358 683200
rect 286526 683144 290774 683200
rect 290942 683144 295190 683200
rect 295358 683144 299606 683200
rect 299774 683144 304114 683200
rect 304282 683144 308530 683200
rect 308698 683144 312946 683200
rect 313114 683144 317454 683200
rect 317622 683144 321870 683200
rect 322038 683144 326286 683200
rect 326454 683144 330702 683200
rect 330870 683144 335210 683200
rect 335378 683144 339626 683200
rect 339794 683144 344042 683200
rect 344210 683144 348458 683200
rect 348626 683144 352966 683200
rect 353134 683144 357382 683200
rect 357550 683144 361798 683200
rect 361966 683144 366214 683200
rect 366382 683144 370722 683200
rect 370890 683144 375138 683200
rect 375306 683144 379554 683200
rect 379722 683144 384062 683200
rect 384230 683144 388478 683200
rect 388646 683144 392894 683200
rect 393062 683144 397310 683200
rect 397478 683144 401818 683200
rect 401986 683144 406234 683200
rect 406402 683144 410650 683200
rect 410818 683144 415066 683200
rect 415234 683144 419574 683200
rect 419742 683144 423990 683200
rect 424158 683144 428406 683200
rect 428574 683144 432822 683200
rect 432990 683144 437330 683200
rect 437498 683144 441746 683200
rect 441914 683144 446162 683200
rect 446330 683144 450670 683200
rect 450838 683144 455086 683200
rect 455254 683144 459502 683200
rect 459670 683144 463918 683200
rect 464086 683144 468426 683200
rect 468594 683144 472842 683200
rect 473010 683144 477258 683200
rect 477426 683144 481674 683200
rect 481842 683144 486182 683200
rect 486350 683144 490598 683200
rect 490766 683144 495014 683200
rect 495182 683144 499430 683200
rect 499598 683144 503938 683200
rect 504106 683144 508354 683200
rect 508522 683144 512770 683200
rect 512938 683144 517278 683200
rect 517446 683144 521694 683200
rect 521862 683144 526110 683200
rect 526278 683144 530526 683200
rect 530694 683144 535034 683200
rect 535202 683144 539450 683200
rect 539618 683144 543866 683200
rect 544034 683144 548282 683200
rect 548450 683144 552790 683200
rect 552958 683144 557206 683200
rect 557374 683144 557476 683200
rect 572 856 557476 683144
rect 682 800 1618 856
rect 1786 800 2722 856
rect 2890 800 3918 856
rect 4086 800 5022 856
rect 5190 800 6126 856
rect 6294 800 7322 856
rect 7490 800 8426 856
rect 8594 800 9530 856
rect 9698 800 10726 856
rect 10894 800 11830 856
rect 11998 800 12934 856
rect 13102 800 14130 856
rect 14298 800 15234 856
rect 15402 800 16338 856
rect 16506 800 17534 856
rect 17702 800 18638 856
rect 18806 800 19742 856
rect 19910 800 20938 856
rect 21106 800 22042 856
rect 22210 800 23146 856
rect 23314 800 24342 856
rect 24510 800 25446 856
rect 25614 800 26550 856
rect 26718 800 27746 856
rect 27914 800 28850 856
rect 29018 800 29954 856
rect 30122 800 31150 856
rect 31318 800 32254 856
rect 32422 800 33358 856
rect 33526 800 34554 856
rect 34722 800 35658 856
rect 35826 800 36762 856
rect 36930 800 37958 856
rect 38126 800 39062 856
rect 39230 800 40166 856
rect 40334 800 41362 856
rect 41530 800 42466 856
rect 42634 800 43570 856
rect 43738 800 44766 856
rect 44934 800 45870 856
rect 46038 800 46974 856
rect 47142 800 48170 856
rect 48338 800 49274 856
rect 49442 800 50378 856
rect 50546 800 51574 856
rect 51742 800 52678 856
rect 52846 800 53782 856
rect 53950 800 54978 856
rect 55146 800 56082 856
rect 56250 800 57186 856
rect 57354 800 58382 856
rect 58550 800 59486 856
rect 59654 800 60590 856
rect 60758 800 61786 856
rect 61954 800 62890 856
rect 63058 800 63994 856
rect 64162 800 65190 856
rect 65358 800 66294 856
rect 66462 800 67398 856
rect 67566 800 68594 856
rect 68762 800 69698 856
rect 69866 800 70802 856
rect 70970 800 71998 856
rect 72166 800 73102 856
rect 73270 800 74206 856
rect 74374 800 75402 856
rect 75570 800 76506 856
rect 76674 800 77610 856
rect 77778 800 78806 856
rect 78974 800 79910 856
rect 80078 800 81014 856
rect 81182 800 82210 856
rect 82378 800 83314 856
rect 83482 800 84418 856
rect 84586 800 85614 856
rect 85782 800 86718 856
rect 86886 800 87822 856
rect 87990 800 89018 856
rect 89186 800 90122 856
rect 90290 800 91226 856
rect 91394 800 92422 856
rect 92590 800 93526 856
rect 93694 800 94630 856
rect 94798 800 95826 856
rect 95994 800 96930 856
rect 97098 800 98034 856
rect 98202 800 99230 856
rect 99398 800 100334 856
rect 100502 800 101438 856
rect 101606 800 102634 856
rect 102802 800 103738 856
rect 103906 800 104842 856
rect 105010 800 106038 856
rect 106206 800 107142 856
rect 107310 800 108246 856
rect 108414 800 109442 856
rect 109610 800 110546 856
rect 110714 800 111650 856
rect 111818 800 112846 856
rect 113014 800 113950 856
rect 114118 800 115054 856
rect 115222 800 116250 856
rect 116418 800 117354 856
rect 117522 800 118458 856
rect 118626 800 119654 856
rect 119822 800 120758 856
rect 120926 800 121862 856
rect 122030 800 123058 856
rect 123226 800 124162 856
rect 124330 800 125266 856
rect 125434 800 126462 856
rect 126630 800 127566 856
rect 127734 800 128670 856
rect 128838 800 129866 856
rect 130034 800 130970 856
rect 131138 800 132074 856
rect 132242 800 133270 856
rect 133438 800 134374 856
rect 134542 800 135478 856
rect 135646 800 136674 856
rect 136842 800 137778 856
rect 137946 800 138882 856
rect 139050 800 140078 856
rect 140246 800 141182 856
rect 141350 800 142286 856
rect 142454 800 143482 856
rect 143650 800 144586 856
rect 144754 800 145690 856
rect 145858 800 146886 856
rect 147054 800 147990 856
rect 148158 800 149094 856
rect 149262 800 150290 856
rect 150458 800 151394 856
rect 151562 800 152498 856
rect 152666 800 153694 856
rect 153862 800 154798 856
rect 154966 800 155902 856
rect 156070 800 157098 856
rect 157266 800 158202 856
rect 158370 800 159306 856
rect 159474 800 160502 856
rect 160670 800 161606 856
rect 161774 800 162710 856
rect 162878 800 163906 856
rect 164074 800 165010 856
rect 165178 800 166114 856
rect 166282 800 167310 856
rect 167478 800 168414 856
rect 168582 800 169518 856
rect 169686 800 170714 856
rect 170882 800 171818 856
rect 171986 800 172922 856
rect 173090 800 174118 856
rect 174286 800 175222 856
rect 175390 800 176326 856
rect 176494 800 177522 856
rect 177690 800 178626 856
rect 178794 800 179730 856
rect 179898 800 180926 856
rect 181094 800 182030 856
rect 182198 800 183134 856
rect 183302 800 184330 856
rect 184498 800 185434 856
rect 185602 800 186538 856
rect 186706 800 187734 856
rect 187902 800 188838 856
rect 189006 800 189942 856
rect 190110 800 191138 856
rect 191306 800 192242 856
rect 192410 800 193346 856
rect 193514 800 194542 856
rect 194710 800 195646 856
rect 195814 800 196750 856
rect 196918 800 197946 856
rect 198114 800 199050 856
rect 199218 800 200154 856
rect 200322 800 201350 856
rect 201518 800 202454 856
rect 202622 800 203558 856
rect 203726 800 204754 856
rect 204922 800 205858 856
rect 206026 800 206962 856
rect 207130 800 208158 856
rect 208326 800 209262 856
rect 209430 800 210366 856
rect 210534 800 211562 856
rect 211730 800 212666 856
rect 212834 800 213770 856
rect 213938 800 214966 856
rect 215134 800 216070 856
rect 216238 800 217174 856
rect 217342 800 218370 856
rect 218538 800 219474 856
rect 219642 800 220578 856
rect 220746 800 221774 856
rect 221942 800 222878 856
rect 223046 800 223982 856
rect 224150 800 225178 856
rect 225346 800 226282 856
rect 226450 800 227386 856
rect 227554 800 228582 856
rect 228750 800 229686 856
rect 229854 800 230790 856
rect 230958 800 231986 856
rect 232154 800 233090 856
rect 233258 800 234194 856
rect 234362 800 235390 856
rect 235558 800 236494 856
rect 236662 800 237598 856
rect 237766 800 238794 856
rect 238962 800 239898 856
rect 240066 800 241002 856
rect 241170 800 242198 856
rect 242366 800 243302 856
rect 243470 800 244406 856
rect 244574 800 245602 856
rect 245770 800 246706 856
rect 246874 800 247810 856
rect 247978 800 249006 856
rect 249174 800 250110 856
rect 250278 800 251214 856
rect 251382 800 252410 856
rect 252578 800 253514 856
rect 253682 800 254618 856
rect 254786 800 255814 856
rect 255982 800 256918 856
rect 257086 800 258022 856
rect 258190 800 259218 856
rect 259386 800 260322 856
rect 260490 800 261426 856
rect 261594 800 262622 856
rect 262790 800 263726 856
rect 263894 800 264830 856
rect 264998 800 266026 856
rect 266194 800 267130 856
rect 267298 800 268234 856
rect 268402 800 269430 856
rect 269598 800 270534 856
rect 270702 800 271638 856
rect 271806 800 272834 856
rect 273002 800 273938 856
rect 274106 800 275042 856
rect 275210 800 276238 856
rect 276406 800 277342 856
rect 277510 800 278446 856
rect 278614 800 279642 856
rect 279810 800 280746 856
rect 280914 800 281850 856
rect 282018 800 283046 856
rect 283214 800 284150 856
rect 284318 800 285254 856
rect 285422 800 286450 856
rect 286618 800 287554 856
rect 287722 800 288658 856
rect 288826 800 289854 856
rect 290022 800 290958 856
rect 291126 800 292062 856
rect 292230 800 293258 856
rect 293426 800 294362 856
rect 294530 800 295466 856
rect 295634 800 296662 856
rect 296830 800 297766 856
rect 297934 800 298870 856
rect 299038 800 300066 856
rect 300234 800 301170 856
rect 301338 800 302274 856
rect 302442 800 303470 856
rect 303638 800 304574 856
rect 304742 800 305678 856
rect 305846 800 306874 856
rect 307042 800 307978 856
rect 308146 800 309082 856
rect 309250 800 310278 856
rect 310446 800 311382 856
rect 311550 800 312486 856
rect 312654 800 313682 856
rect 313850 800 314786 856
rect 314954 800 315890 856
rect 316058 800 317086 856
rect 317254 800 318190 856
rect 318358 800 319294 856
rect 319462 800 320490 856
rect 320658 800 321594 856
rect 321762 800 322698 856
rect 322866 800 323894 856
rect 324062 800 324998 856
rect 325166 800 326102 856
rect 326270 800 327298 856
rect 327466 800 328402 856
rect 328570 800 329506 856
rect 329674 800 330702 856
rect 330870 800 331806 856
rect 331974 800 332910 856
rect 333078 800 334106 856
rect 334274 800 335210 856
rect 335378 800 336314 856
rect 336482 800 337510 856
rect 337678 800 338614 856
rect 338782 800 339718 856
rect 339886 800 340914 856
rect 341082 800 342018 856
rect 342186 800 343122 856
rect 343290 800 344318 856
rect 344486 800 345422 856
rect 345590 800 346526 856
rect 346694 800 347722 856
rect 347890 800 348826 856
rect 348994 800 349930 856
rect 350098 800 351126 856
rect 351294 800 352230 856
rect 352398 800 353334 856
rect 353502 800 354530 856
rect 354698 800 355634 856
rect 355802 800 356738 856
rect 356906 800 357934 856
rect 358102 800 359038 856
rect 359206 800 360142 856
rect 360310 800 361338 856
rect 361506 800 362442 856
rect 362610 800 363546 856
rect 363714 800 364742 856
rect 364910 800 365846 856
rect 366014 800 366950 856
rect 367118 800 368146 856
rect 368314 800 369250 856
rect 369418 800 370354 856
rect 370522 800 371550 856
rect 371718 800 372654 856
rect 372822 800 373758 856
rect 373926 800 374954 856
rect 375122 800 376058 856
rect 376226 800 377162 856
rect 377330 800 378358 856
rect 378526 800 379462 856
rect 379630 800 380566 856
rect 380734 800 381762 856
rect 381930 800 382866 856
rect 383034 800 383970 856
rect 384138 800 385166 856
rect 385334 800 386270 856
rect 386438 800 387374 856
rect 387542 800 388570 856
rect 388738 800 389674 856
rect 389842 800 390778 856
rect 390946 800 391974 856
rect 392142 800 393078 856
rect 393246 800 394182 856
rect 394350 800 395378 856
rect 395546 800 396482 856
rect 396650 800 397586 856
rect 397754 800 398782 856
rect 398950 800 399886 856
rect 400054 800 400990 856
rect 401158 800 402186 856
rect 402354 800 403290 856
rect 403458 800 404394 856
rect 404562 800 405590 856
rect 405758 800 406694 856
rect 406862 800 407798 856
rect 407966 800 408994 856
rect 409162 800 410098 856
rect 410266 800 411202 856
rect 411370 800 412398 856
rect 412566 800 413502 856
rect 413670 800 414606 856
rect 414774 800 415802 856
rect 415970 800 416906 856
rect 417074 800 418010 856
rect 418178 800 419206 856
rect 419374 800 420310 856
rect 420478 800 421414 856
rect 421582 800 422610 856
rect 422778 800 423714 856
rect 423882 800 424818 856
rect 424986 800 426014 856
rect 426182 800 427118 856
rect 427286 800 428222 856
rect 428390 800 429418 856
rect 429586 800 430522 856
rect 430690 800 431626 856
rect 431794 800 432822 856
rect 432990 800 433926 856
rect 434094 800 435030 856
rect 435198 800 436226 856
rect 436394 800 437330 856
rect 437498 800 438434 856
rect 438602 800 439630 856
rect 439798 800 440734 856
rect 440902 800 441838 856
rect 442006 800 443034 856
rect 443202 800 444138 856
rect 444306 800 445242 856
rect 445410 800 446438 856
rect 446606 800 447542 856
rect 447710 800 448646 856
rect 448814 800 449842 856
rect 450010 800 450946 856
rect 451114 800 452050 856
rect 452218 800 453246 856
rect 453414 800 454350 856
rect 454518 800 455454 856
rect 455622 800 456650 856
rect 456818 800 457754 856
rect 457922 800 458858 856
rect 459026 800 460054 856
rect 460222 800 461158 856
rect 461326 800 462262 856
rect 462430 800 463458 856
rect 463626 800 464562 856
rect 464730 800 465666 856
rect 465834 800 466862 856
rect 467030 800 467966 856
rect 468134 800 469070 856
rect 469238 800 470266 856
rect 470434 800 471370 856
rect 471538 800 472474 856
rect 472642 800 473670 856
rect 473838 800 474774 856
rect 474942 800 475878 856
rect 476046 800 477074 856
rect 477242 800 478178 856
rect 478346 800 479282 856
rect 479450 800 480478 856
rect 480646 800 481582 856
rect 481750 800 482686 856
rect 482854 800 483882 856
rect 484050 800 484986 856
rect 485154 800 486090 856
rect 486258 800 487286 856
rect 487454 800 488390 856
rect 488558 800 489494 856
rect 489662 800 490690 856
rect 490858 800 491794 856
rect 491962 800 492898 856
rect 493066 800 494094 856
rect 494262 800 495198 856
rect 495366 800 496302 856
rect 496470 800 497498 856
rect 497666 800 498602 856
rect 498770 800 499706 856
rect 499874 800 500902 856
rect 501070 800 502006 856
rect 502174 800 503110 856
rect 503278 800 504306 856
rect 504474 800 505410 856
rect 505578 800 506514 856
rect 506682 800 507710 856
rect 507878 800 508814 856
rect 508982 800 509918 856
rect 510086 800 511114 856
rect 511282 800 512218 856
rect 512386 800 513322 856
rect 513490 800 514518 856
rect 514686 800 515622 856
rect 515790 800 516726 856
rect 516894 800 517922 856
rect 518090 800 519026 856
rect 519194 800 520130 856
rect 520298 800 521326 856
rect 521494 800 522430 856
rect 522598 800 523534 856
rect 523702 800 524730 856
rect 524898 800 525834 856
rect 526002 800 526938 856
rect 527106 800 528134 856
rect 528302 800 529238 856
rect 529406 800 530342 856
rect 530510 800 531538 856
rect 531706 800 532642 856
rect 532810 800 533746 856
rect 533914 800 534942 856
rect 535110 800 536046 856
rect 536214 800 537150 856
rect 537318 800 538346 856
rect 538514 800 539450 856
rect 539618 800 540554 856
rect 540722 800 541750 856
rect 541918 800 542854 856
rect 543022 800 543958 856
rect 544126 800 545154 856
rect 545322 800 546258 856
rect 546426 800 547362 856
rect 547530 800 548558 856
rect 548726 800 549662 856
rect 549830 800 550766 856
rect 550934 800 551962 856
rect 552130 800 553066 856
rect 553234 800 554170 856
rect 554338 800 555366 856
rect 555534 800 556470 856
rect 556638 800 557476 856
<< metal3 >>
rect 0 598272 800 598392
rect 0 427320 800 427440
rect 0 256368 800 256488
rect 0 85416 800 85536
rect 563200 641112 564000 641232
rect 563200 555568 564000 555688
rect 563200 470160 564000 470280
rect 563200 384616 564000 384736
rect 563200 299072 564000 299192
rect 563200 213664 564000 213784
rect 563200 128120 564000 128240
rect 563200 42712 564000 42832
<< obsm3 >>
rect 2681 2143 557488 681665
<< metal4 >>
rect 4208 2128 4528 681680
rect 19568 2128 19888 681680
rect 34928 2128 35248 681680
rect 50288 2128 50608 681680
rect 65648 2128 65968 681680
rect 81008 2128 81328 681680
rect 96368 2128 96688 681680
rect 111728 2128 112048 681680
rect 127088 2128 127408 681680
rect 142448 2128 142768 681680
rect 157808 2128 158128 681680
rect 173168 2128 173488 681680
rect 188528 2128 188848 681680
rect 203888 2128 204208 681680
rect 219248 2128 219568 681680
rect 234608 2128 234928 681680
rect 249968 2128 250288 681680
rect 265328 2128 265648 681680
rect 280688 2128 281008 681680
rect 296048 2128 296368 681680
rect 311408 2128 311728 681680
rect 326768 2128 327088 681680
rect 342128 2128 342448 681680
rect 357488 2128 357808 681680
rect 372848 2128 373168 681680
rect 388208 2128 388528 681680
rect 403568 2128 403888 681680
rect 418928 2128 419248 681680
rect 434288 2128 434608 681680
rect 449648 2128 449968 681680
rect 465008 2128 465328 681680
rect 480368 2128 480688 681680
rect 495728 2128 496048 681680
rect 511088 2128 511408 681680
rect 526448 2128 526768 681680
rect 541808 2128 542128 681680
rect 557168 2128 557488 681680
<< obsm4 >>
rect 2819 9147 4128 675885
rect 4608 9147 19488 675885
rect 19968 9147 34848 675885
rect 35328 9147 50208 675885
rect 50688 9147 65568 675885
rect 66048 9147 80928 675885
rect 81408 9147 96288 675885
rect 96768 9147 111648 675885
rect 112128 9147 127008 675885
rect 127488 9147 142368 675885
rect 142848 9147 157728 675885
rect 158208 9147 173088 675885
rect 173568 9147 188448 675885
rect 188928 9147 203808 675885
rect 204288 9147 219168 675885
rect 219648 9147 234528 675885
rect 235008 9147 249888 675885
rect 250368 9147 265248 675885
rect 265728 9147 280608 675885
rect 281088 9147 295968 675885
rect 296448 9147 311328 675885
rect 311808 9147 326688 675885
rect 327168 9147 342048 675885
rect 342528 9147 357408 675885
rect 357888 9147 372768 675885
rect 373248 9147 388128 675885
rect 388608 9147 403488 675885
rect 403968 9147 418848 675885
rect 419328 9147 434208 675885
rect 434688 9147 449568 675885
rect 450048 9147 464928 675885
rect 465408 9147 480288 675885
rect 480768 9147 495648 675885
rect 496128 9147 511008 675885
rect 511488 9147 526368 675885
rect 526848 9147 541728 675885
rect 542208 9147 545317 675885
<< labels >>
rlabel metal2 s 508410 683200 508466 684000 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal3 s 563200 213664 564000 213784 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal3 s 0 256368 800 256488 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 539506 683200 539562 684000 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal3 s 563200 299072 564000 299192 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 557630 0 557686 800 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal3 s 0 427320 800 427440 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 558826 0 558882 800 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal2 s 543922 683200 543978 684000 6 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal2 s 559930 0 559986 800 6 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal2 s 548338 683200 548394 684000 6 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal2 s 512826 683200 512882 684000 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s 0 598272 800 598392 6 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal2 s 561034 0 561090 800 6 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s 563200 384616 564000 384736 6 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal2 s 562230 0 562286 800 6 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal2 s 552846 683200 552902 684000 6 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s 563200 470160 564000 470280 6 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal2 s 563334 0 563390 800 6 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s 563200 555568 564000 555688 6 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal2 s 557262 683200 557318 684000 6 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 563200 641112 564000 641232 6 analog_io[29]
port 22 nsew signal bidirectional
rlabel metal2 s 517334 683200 517390 684000 6 analog_io[2]
port 23 nsew signal bidirectional
rlabel metal2 s 561678 683200 561734 684000 6 analog_io[30]
port 24 nsew signal bidirectional
rlabel metal3 s 563200 42712 564000 42832 6 analog_io[3]
port 25 nsew signal bidirectional
rlabel metal2 s 521750 683200 521806 684000 6 analog_io[4]
port 26 nsew signal bidirectional
rlabel metal3 s 563200 128120 564000 128240 6 analog_io[5]
port 27 nsew signal bidirectional
rlabel metal3 s 0 85416 800 85536 6 analog_io[6]
port 28 nsew signal bidirectional
rlabel metal2 s 526166 683200 526222 684000 6 analog_io[7]
port 29 nsew signal bidirectional
rlabel metal2 s 530582 683200 530638 684000 6 analog_io[8]
port 30 nsew signal bidirectional
rlabel metal2 s 535090 683200 535146 684000 6 analog_io[9]
port 31 nsew signal bidirectional
rlabel metal2 s 2226 683200 2282 684000 6 io_in[0]
port 32 nsew signal input
rlabel metal2 s 135442 683200 135498 684000 6 io_in[10]
port 33 nsew signal input
rlabel metal2 s 148690 683200 148746 684000 6 io_in[11]
port 34 nsew signal input
rlabel metal2 s 162030 683200 162086 684000 6 io_in[12]
port 35 nsew signal input
rlabel metal2 s 175370 683200 175426 684000 6 io_in[13]
port 36 nsew signal input
rlabel metal2 s 188710 683200 188766 684000 6 io_in[14]
port 37 nsew signal input
rlabel metal2 s 202050 683200 202106 684000 6 io_in[15]
port 38 nsew signal input
rlabel metal2 s 215298 683200 215354 684000 6 io_in[16]
port 39 nsew signal input
rlabel metal2 s 228638 683200 228694 684000 6 io_in[17]
port 40 nsew signal input
rlabel metal2 s 241978 683200 242034 684000 6 io_in[18]
port 41 nsew signal input
rlabel metal2 s 255318 683200 255374 684000 6 io_in[19]
port 42 nsew signal input
rlabel metal2 s 15474 683200 15530 684000 6 io_in[1]
port 43 nsew signal input
rlabel metal2 s 268658 683200 268714 684000 6 io_in[20]
port 44 nsew signal input
rlabel metal2 s 281906 683200 281962 684000 6 io_in[21]
port 45 nsew signal input
rlabel metal2 s 295246 683200 295302 684000 6 io_in[22]
port 46 nsew signal input
rlabel metal2 s 308586 683200 308642 684000 6 io_in[23]
port 47 nsew signal input
rlabel metal2 s 321926 683200 321982 684000 6 io_in[24]
port 48 nsew signal input
rlabel metal2 s 335266 683200 335322 684000 6 io_in[25]
port 49 nsew signal input
rlabel metal2 s 348514 683200 348570 684000 6 io_in[26]
port 50 nsew signal input
rlabel metal2 s 361854 683200 361910 684000 6 io_in[27]
port 51 nsew signal input
rlabel metal2 s 375194 683200 375250 684000 6 io_in[28]
port 52 nsew signal input
rlabel metal2 s 388534 683200 388590 684000 6 io_in[29]
port 53 nsew signal input
rlabel metal2 s 28814 683200 28870 684000 6 io_in[2]
port 54 nsew signal input
rlabel metal2 s 401874 683200 401930 684000 6 io_in[30]
port 55 nsew signal input
rlabel metal2 s 415122 683200 415178 684000 6 io_in[31]
port 56 nsew signal input
rlabel metal2 s 428462 683200 428518 684000 6 io_in[32]
port 57 nsew signal input
rlabel metal2 s 441802 683200 441858 684000 6 io_in[33]
port 58 nsew signal input
rlabel metal2 s 455142 683200 455198 684000 6 io_in[34]
port 59 nsew signal input
rlabel metal2 s 468482 683200 468538 684000 6 io_in[35]
port 60 nsew signal input
rlabel metal2 s 481730 683200 481786 684000 6 io_in[36]
port 61 nsew signal input
rlabel metal2 s 495070 683200 495126 684000 6 io_in[37]
port 62 nsew signal input
rlabel metal2 s 42154 683200 42210 684000 6 io_in[3]
port 63 nsew signal input
rlabel metal2 s 55494 683200 55550 684000 6 io_in[4]
port 64 nsew signal input
rlabel metal2 s 68834 683200 68890 684000 6 io_in[5]
port 65 nsew signal input
rlabel metal2 s 82082 683200 82138 684000 6 io_in[6]
port 66 nsew signal input
rlabel metal2 s 95422 683200 95478 684000 6 io_in[7]
port 67 nsew signal input
rlabel metal2 s 108762 683200 108818 684000 6 io_in[8]
port 68 nsew signal input
rlabel metal2 s 122102 683200 122158 684000 6 io_in[9]
port 69 nsew signal input
rlabel metal2 s 6642 683200 6698 684000 6 io_oeb[0]
port 70 nsew signal output
rlabel metal2 s 139858 683200 139914 684000 6 io_oeb[10]
port 71 nsew signal output
rlabel metal2 s 153198 683200 153254 684000 6 io_oeb[11]
port 72 nsew signal output
rlabel metal2 s 166446 683200 166502 684000 6 io_oeb[12]
port 73 nsew signal output
rlabel metal2 s 179786 683200 179842 684000 6 io_oeb[13]
port 74 nsew signal output
rlabel metal2 s 193126 683200 193182 684000 6 io_oeb[14]
port 75 nsew signal output
rlabel metal2 s 206466 683200 206522 684000 6 io_oeb[15]
port 76 nsew signal output
rlabel metal2 s 219806 683200 219862 684000 6 io_oeb[16]
port 77 nsew signal output
rlabel metal2 s 233054 683200 233110 684000 6 io_oeb[17]
port 78 nsew signal output
rlabel metal2 s 246394 683200 246450 684000 6 io_oeb[18]
port 79 nsew signal output
rlabel metal2 s 259734 683200 259790 684000 6 io_oeb[19]
port 80 nsew signal output
rlabel metal2 s 19982 683200 20038 684000 6 io_oeb[1]
port 81 nsew signal output
rlabel metal2 s 273074 683200 273130 684000 6 io_oeb[20]
port 82 nsew signal output
rlabel metal2 s 286414 683200 286470 684000 6 io_oeb[21]
port 83 nsew signal output
rlabel metal2 s 299662 683200 299718 684000 6 io_oeb[22]
port 84 nsew signal output
rlabel metal2 s 313002 683200 313058 684000 6 io_oeb[23]
port 85 nsew signal output
rlabel metal2 s 326342 683200 326398 684000 6 io_oeb[24]
port 86 nsew signal output
rlabel metal2 s 339682 683200 339738 684000 6 io_oeb[25]
port 87 nsew signal output
rlabel metal2 s 353022 683200 353078 684000 6 io_oeb[26]
port 88 nsew signal output
rlabel metal2 s 366270 683200 366326 684000 6 io_oeb[27]
port 89 nsew signal output
rlabel metal2 s 379610 683200 379666 684000 6 io_oeb[28]
port 90 nsew signal output
rlabel metal2 s 392950 683200 393006 684000 6 io_oeb[29]
port 91 nsew signal output
rlabel metal2 s 33230 683200 33286 684000 6 io_oeb[2]
port 92 nsew signal output
rlabel metal2 s 406290 683200 406346 684000 6 io_oeb[30]
port 93 nsew signal output
rlabel metal2 s 419630 683200 419686 684000 6 io_oeb[31]
port 94 nsew signal output
rlabel metal2 s 432878 683200 432934 684000 6 io_oeb[32]
port 95 nsew signal output
rlabel metal2 s 446218 683200 446274 684000 6 io_oeb[33]
port 96 nsew signal output
rlabel metal2 s 459558 683200 459614 684000 6 io_oeb[34]
port 97 nsew signal output
rlabel metal2 s 472898 683200 472954 684000 6 io_oeb[35]
port 98 nsew signal output
rlabel metal2 s 486238 683200 486294 684000 6 io_oeb[36]
port 99 nsew signal output
rlabel metal2 s 499486 683200 499542 684000 6 io_oeb[37]
port 100 nsew signal output
rlabel metal2 s 46570 683200 46626 684000 6 io_oeb[3]
port 101 nsew signal output
rlabel metal2 s 59910 683200 59966 684000 6 io_oeb[4]
port 102 nsew signal output
rlabel metal2 s 73250 683200 73306 684000 6 io_oeb[5]
port 103 nsew signal output
rlabel metal2 s 86590 683200 86646 684000 6 io_oeb[6]
port 104 nsew signal output
rlabel metal2 s 99838 683200 99894 684000 6 io_oeb[7]
port 105 nsew signal output
rlabel metal2 s 113178 683200 113234 684000 6 io_oeb[8]
port 106 nsew signal output
rlabel metal2 s 126518 683200 126574 684000 6 io_oeb[9]
port 107 nsew signal output
rlabel metal2 s 11058 683200 11114 684000 6 io_out[0]
port 108 nsew signal output
rlabel metal2 s 144274 683200 144330 684000 6 io_out[10]
port 109 nsew signal output
rlabel metal2 s 157614 683200 157670 684000 6 io_out[11]
port 110 nsew signal output
rlabel metal2 s 170954 683200 171010 684000 6 io_out[12]
port 111 nsew signal output
rlabel metal2 s 184202 683200 184258 684000 6 io_out[13]
port 112 nsew signal output
rlabel metal2 s 197542 683200 197598 684000 6 io_out[14]
port 113 nsew signal output
rlabel metal2 s 210882 683200 210938 684000 6 io_out[15]
port 114 nsew signal output
rlabel metal2 s 224222 683200 224278 684000 6 io_out[16]
port 115 nsew signal output
rlabel metal2 s 237562 683200 237618 684000 6 io_out[17]
port 116 nsew signal output
rlabel metal2 s 250810 683200 250866 684000 6 io_out[18]
port 117 nsew signal output
rlabel metal2 s 264150 683200 264206 684000 6 io_out[19]
port 118 nsew signal output
rlabel metal2 s 24398 683200 24454 684000 6 io_out[1]
port 119 nsew signal output
rlabel metal2 s 277490 683200 277546 684000 6 io_out[20]
port 120 nsew signal output
rlabel metal2 s 290830 683200 290886 684000 6 io_out[21]
port 121 nsew signal output
rlabel metal2 s 304170 683200 304226 684000 6 io_out[22]
port 122 nsew signal output
rlabel metal2 s 317510 683200 317566 684000 6 io_out[23]
port 123 nsew signal output
rlabel metal2 s 330758 683200 330814 684000 6 io_out[24]
port 124 nsew signal output
rlabel metal2 s 344098 683200 344154 684000 6 io_out[25]
port 125 nsew signal output
rlabel metal2 s 357438 683200 357494 684000 6 io_out[26]
port 126 nsew signal output
rlabel metal2 s 370778 683200 370834 684000 6 io_out[27]
port 127 nsew signal output
rlabel metal2 s 384118 683200 384174 684000 6 io_out[28]
port 128 nsew signal output
rlabel metal2 s 397366 683200 397422 684000 6 io_out[29]
port 129 nsew signal output
rlabel metal2 s 37738 683200 37794 684000 6 io_out[2]
port 130 nsew signal output
rlabel metal2 s 410706 683200 410762 684000 6 io_out[30]
port 131 nsew signal output
rlabel metal2 s 424046 683200 424102 684000 6 io_out[31]
port 132 nsew signal output
rlabel metal2 s 437386 683200 437442 684000 6 io_out[32]
port 133 nsew signal output
rlabel metal2 s 450726 683200 450782 684000 6 io_out[33]
port 134 nsew signal output
rlabel metal2 s 463974 683200 464030 684000 6 io_out[34]
port 135 nsew signal output
rlabel metal2 s 477314 683200 477370 684000 6 io_out[35]
port 136 nsew signal output
rlabel metal2 s 490654 683200 490710 684000 6 io_out[36]
port 137 nsew signal output
rlabel metal2 s 503994 683200 504050 684000 6 io_out[37]
port 138 nsew signal output
rlabel metal2 s 50986 683200 51042 684000 6 io_out[3]
port 139 nsew signal output
rlabel metal2 s 64326 683200 64382 684000 6 io_out[4]
port 140 nsew signal output
rlabel metal2 s 77666 683200 77722 684000 6 io_out[5]
port 141 nsew signal output
rlabel metal2 s 91006 683200 91062 684000 6 io_out[6]
port 142 nsew signal output
rlabel metal2 s 104346 683200 104402 684000 6 io_out[7]
port 143 nsew signal output
rlabel metal2 s 117594 683200 117650 684000 6 io_out[8]
port 144 nsew signal output
rlabel metal2 s 130934 683200 130990 684000 6 io_out[9]
port 145 nsew signal output
rlabel metal2 s 120814 0 120870 800 6 la_data_in[0]
port 146 nsew signal input
rlabel metal2 s 461214 0 461270 800 6 la_data_in[100]
port 147 nsew signal input
rlabel metal2 s 464618 0 464674 800 6 la_data_in[101]
port 148 nsew signal input
rlabel metal2 s 468022 0 468078 800 6 la_data_in[102]
port 149 nsew signal input
rlabel metal2 s 471426 0 471482 800 6 la_data_in[103]
port 150 nsew signal input
rlabel metal2 s 474830 0 474886 800 6 la_data_in[104]
port 151 nsew signal input
rlabel metal2 s 478234 0 478290 800 6 la_data_in[105]
port 152 nsew signal input
rlabel metal2 s 481638 0 481694 800 6 la_data_in[106]
port 153 nsew signal input
rlabel metal2 s 485042 0 485098 800 6 la_data_in[107]
port 154 nsew signal input
rlabel metal2 s 488446 0 488502 800 6 la_data_in[108]
port 155 nsew signal input
rlabel metal2 s 491850 0 491906 800 6 la_data_in[109]
port 156 nsew signal input
rlabel metal2 s 154854 0 154910 800 6 la_data_in[10]
port 157 nsew signal input
rlabel metal2 s 495254 0 495310 800 6 la_data_in[110]
port 158 nsew signal input
rlabel metal2 s 498658 0 498714 800 6 la_data_in[111]
port 159 nsew signal input
rlabel metal2 s 502062 0 502118 800 6 la_data_in[112]
port 160 nsew signal input
rlabel metal2 s 505466 0 505522 800 6 la_data_in[113]
port 161 nsew signal input
rlabel metal2 s 508870 0 508926 800 6 la_data_in[114]
port 162 nsew signal input
rlabel metal2 s 512274 0 512330 800 6 la_data_in[115]
port 163 nsew signal input
rlabel metal2 s 515678 0 515734 800 6 la_data_in[116]
port 164 nsew signal input
rlabel metal2 s 519082 0 519138 800 6 la_data_in[117]
port 165 nsew signal input
rlabel metal2 s 522486 0 522542 800 6 la_data_in[118]
port 166 nsew signal input
rlabel metal2 s 525890 0 525946 800 6 la_data_in[119]
port 167 nsew signal input
rlabel metal2 s 158258 0 158314 800 6 la_data_in[11]
port 168 nsew signal input
rlabel metal2 s 529294 0 529350 800 6 la_data_in[120]
port 169 nsew signal input
rlabel metal2 s 532698 0 532754 800 6 la_data_in[121]
port 170 nsew signal input
rlabel metal2 s 536102 0 536158 800 6 la_data_in[122]
port 171 nsew signal input
rlabel metal2 s 539506 0 539562 800 6 la_data_in[123]
port 172 nsew signal input
rlabel metal2 s 542910 0 542966 800 6 la_data_in[124]
port 173 nsew signal input
rlabel metal2 s 546314 0 546370 800 6 la_data_in[125]
port 174 nsew signal input
rlabel metal2 s 549718 0 549774 800 6 la_data_in[126]
port 175 nsew signal input
rlabel metal2 s 553122 0 553178 800 6 la_data_in[127]
port 176 nsew signal input
rlabel metal2 s 161662 0 161718 800 6 la_data_in[12]
port 177 nsew signal input
rlabel metal2 s 165066 0 165122 800 6 la_data_in[13]
port 178 nsew signal input
rlabel metal2 s 168470 0 168526 800 6 la_data_in[14]
port 179 nsew signal input
rlabel metal2 s 171874 0 171930 800 6 la_data_in[15]
port 180 nsew signal input
rlabel metal2 s 175278 0 175334 800 6 la_data_in[16]
port 181 nsew signal input
rlabel metal2 s 178682 0 178738 800 6 la_data_in[17]
port 182 nsew signal input
rlabel metal2 s 182086 0 182142 800 6 la_data_in[18]
port 183 nsew signal input
rlabel metal2 s 185490 0 185546 800 6 la_data_in[19]
port 184 nsew signal input
rlabel metal2 s 124218 0 124274 800 6 la_data_in[1]
port 185 nsew signal input
rlabel metal2 s 188894 0 188950 800 6 la_data_in[20]
port 186 nsew signal input
rlabel metal2 s 192298 0 192354 800 6 la_data_in[21]
port 187 nsew signal input
rlabel metal2 s 195702 0 195758 800 6 la_data_in[22]
port 188 nsew signal input
rlabel metal2 s 199106 0 199162 800 6 la_data_in[23]
port 189 nsew signal input
rlabel metal2 s 202510 0 202566 800 6 la_data_in[24]
port 190 nsew signal input
rlabel metal2 s 205914 0 205970 800 6 la_data_in[25]
port 191 nsew signal input
rlabel metal2 s 209318 0 209374 800 6 la_data_in[26]
port 192 nsew signal input
rlabel metal2 s 212722 0 212778 800 6 la_data_in[27]
port 193 nsew signal input
rlabel metal2 s 216126 0 216182 800 6 la_data_in[28]
port 194 nsew signal input
rlabel metal2 s 219530 0 219586 800 6 la_data_in[29]
port 195 nsew signal input
rlabel metal2 s 127622 0 127678 800 6 la_data_in[2]
port 196 nsew signal input
rlabel metal2 s 222934 0 222990 800 6 la_data_in[30]
port 197 nsew signal input
rlabel metal2 s 226338 0 226394 800 6 la_data_in[31]
port 198 nsew signal input
rlabel metal2 s 229742 0 229798 800 6 la_data_in[32]
port 199 nsew signal input
rlabel metal2 s 233146 0 233202 800 6 la_data_in[33]
port 200 nsew signal input
rlabel metal2 s 236550 0 236606 800 6 la_data_in[34]
port 201 nsew signal input
rlabel metal2 s 239954 0 240010 800 6 la_data_in[35]
port 202 nsew signal input
rlabel metal2 s 243358 0 243414 800 6 la_data_in[36]
port 203 nsew signal input
rlabel metal2 s 246762 0 246818 800 6 la_data_in[37]
port 204 nsew signal input
rlabel metal2 s 250166 0 250222 800 6 la_data_in[38]
port 205 nsew signal input
rlabel metal2 s 253570 0 253626 800 6 la_data_in[39]
port 206 nsew signal input
rlabel metal2 s 131026 0 131082 800 6 la_data_in[3]
port 207 nsew signal input
rlabel metal2 s 256974 0 257030 800 6 la_data_in[40]
port 208 nsew signal input
rlabel metal2 s 260378 0 260434 800 6 la_data_in[41]
port 209 nsew signal input
rlabel metal2 s 263782 0 263838 800 6 la_data_in[42]
port 210 nsew signal input
rlabel metal2 s 267186 0 267242 800 6 la_data_in[43]
port 211 nsew signal input
rlabel metal2 s 270590 0 270646 800 6 la_data_in[44]
port 212 nsew signal input
rlabel metal2 s 273994 0 274050 800 6 la_data_in[45]
port 213 nsew signal input
rlabel metal2 s 277398 0 277454 800 6 la_data_in[46]
port 214 nsew signal input
rlabel metal2 s 280802 0 280858 800 6 la_data_in[47]
port 215 nsew signal input
rlabel metal2 s 284206 0 284262 800 6 la_data_in[48]
port 216 nsew signal input
rlabel metal2 s 287610 0 287666 800 6 la_data_in[49]
port 217 nsew signal input
rlabel metal2 s 134430 0 134486 800 6 la_data_in[4]
port 218 nsew signal input
rlabel metal2 s 291014 0 291070 800 6 la_data_in[50]
port 219 nsew signal input
rlabel metal2 s 294418 0 294474 800 6 la_data_in[51]
port 220 nsew signal input
rlabel metal2 s 297822 0 297878 800 6 la_data_in[52]
port 221 nsew signal input
rlabel metal2 s 301226 0 301282 800 6 la_data_in[53]
port 222 nsew signal input
rlabel metal2 s 304630 0 304686 800 6 la_data_in[54]
port 223 nsew signal input
rlabel metal2 s 308034 0 308090 800 6 la_data_in[55]
port 224 nsew signal input
rlabel metal2 s 311438 0 311494 800 6 la_data_in[56]
port 225 nsew signal input
rlabel metal2 s 314842 0 314898 800 6 la_data_in[57]
port 226 nsew signal input
rlabel metal2 s 318246 0 318302 800 6 la_data_in[58]
port 227 nsew signal input
rlabel metal2 s 321650 0 321706 800 6 la_data_in[59]
port 228 nsew signal input
rlabel metal2 s 137834 0 137890 800 6 la_data_in[5]
port 229 nsew signal input
rlabel metal2 s 325054 0 325110 800 6 la_data_in[60]
port 230 nsew signal input
rlabel metal2 s 328458 0 328514 800 6 la_data_in[61]
port 231 nsew signal input
rlabel metal2 s 331862 0 331918 800 6 la_data_in[62]
port 232 nsew signal input
rlabel metal2 s 335266 0 335322 800 6 la_data_in[63]
port 233 nsew signal input
rlabel metal2 s 338670 0 338726 800 6 la_data_in[64]
port 234 nsew signal input
rlabel metal2 s 342074 0 342130 800 6 la_data_in[65]
port 235 nsew signal input
rlabel metal2 s 345478 0 345534 800 6 la_data_in[66]
port 236 nsew signal input
rlabel metal2 s 348882 0 348938 800 6 la_data_in[67]
port 237 nsew signal input
rlabel metal2 s 352286 0 352342 800 6 la_data_in[68]
port 238 nsew signal input
rlabel metal2 s 355690 0 355746 800 6 la_data_in[69]
port 239 nsew signal input
rlabel metal2 s 141238 0 141294 800 6 la_data_in[6]
port 240 nsew signal input
rlabel metal2 s 359094 0 359150 800 6 la_data_in[70]
port 241 nsew signal input
rlabel metal2 s 362498 0 362554 800 6 la_data_in[71]
port 242 nsew signal input
rlabel metal2 s 365902 0 365958 800 6 la_data_in[72]
port 243 nsew signal input
rlabel metal2 s 369306 0 369362 800 6 la_data_in[73]
port 244 nsew signal input
rlabel metal2 s 372710 0 372766 800 6 la_data_in[74]
port 245 nsew signal input
rlabel metal2 s 376114 0 376170 800 6 la_data_in[75]
port 246 nsew signal input
rlabel metal2 s 379518 0 379574 800 6 la_data_in[76]
port 247 nsew signal input
rlabel metal2 s 382922 0 382978 800 6 la_data_in[77]
port 248 nsew signal input
rlabel metal2 s 386326 0 386382 800 6 la_data_in[78]
port 249 nsew signal input
rlabel metal2 s 389730 0 389786 800 6 la_data_in[79]
port 250 nsew signal input
rlabel metal2 s 144642 0 144698 800 6 la_data_in[7]
port 251 nsew signal input
rlabel metal2 s 393134 0 393190 800 6 la_data_in[80]
port 252 nsew signal input
rlabel metal2 s 396538 0 396594 800 6 la_data_in[81]
port 253 nsew signal input
rlabel metal2 s 399942 0 399998 800 6 la_data_in[82]
port 254 nsew signal input
rlabel metal2 s 403346 0 403402 800 6 la_data_in[83]
port 255 nsew signal input
rlabel metal2 s 406750 0 406806 800 6 la_data_in[84]
port 256 nsew signal input
rlabel metal2 s 410154 0 410210 800 6 la_data_in[85]
port 257 nsew signal input
rlabel metal2 s 413558 0 413614 800 6 la_data_in[86]
port 258 nsew signal input
rlabel metal2 s 416962 0 417018 800 6 la_data_in[87]
port 259 nsew signal input
rlabel metal2 s 420366 0 420422 800 6 la_data_in[88]
port 260 nsew signal input
rlabel metal2 s 423770 0 423826 800 6 la_data_in[89]
port 261 nsew signal input
rlabel metal2 s 148046 0 148102 800 6 la_data_in[8]
port 262 nsew signal input
rlabel metal2 s 427174 0 427230 800 6 la_data_in[90]
port 263 nsew signal input
rlabel metal2 s 430578 0 430634 800 6 la_data_in[91]
port 264 nsew signal input
rlabel metal2 s 433982 0 434038 800 6 la_data_in[92]
port 265 nsew signal input
rlabel metal2 s 437386 0 437442 800 6 la_data_in[93]
port 266 nsew signal input
rlabel metal2 s 440790 0 440846 800 6 la_data_in[94]
port 267 nsew signal input
rlabel metal2 s 444194 0 444250 800 6 la_data_in[95]
port 268 nsew signal input
rlabel metal2 s 447598 0 447654 800 6 la_data_in[96]
port 269 nsew signal input
rlabel metal2 s 451002 0 451058 800 6 la_data_in[97]
port 270 nsew signal input
rlabel metal2 s 454406 0 454462 800 6 la_data_in[98]
port 271 nsew signal input
rlabel metal2 s 457810 0 457866 800 6 la_data_in[99]
port 272 nsew signal input
rlabel metal2 s 151450 0 151506 800 6 la_data_in[9]
port 273 nsew signal input
rlabel metal2 s 121918 0 121974 800 6 la_data_out[0]
port 274 nsew signal output
rlabel metal2 s 462318 0 462374 800 6 la_data_out[100]
port 275 nsew signal output
rlabel metal2 s 465722 0 465778 800 6 la_data_out[101]
port 276 nsew signal output
rlabel metal2 s 469126 0 469182 800 6 la_data_out[102]
port 277 nsew signal output
rlabel metal2 s 472530 0 472586 800 6 la_data_out[103]
port 278 nsew signal output
rlabel metal2 s 475934 0 475990 800 6 la_data_out[104]
port 279 nsew signal output
rlabel metal2 s 479338 0 479394 800 6 la_data_out[105]
port 280 nsew signal output
rlabel metal2 s 482742 0 482798 800 6 la_data_out[106]
port 281 nsew signal output
rlabel metal2 s 486146 0 486202 800 6 la_data_out[107]
port 282 nsew signal output
rlabel metal2 s 489550 0 489606 800 6 la_data_out[108]
port 283 nsew signal output
rlabel metal2 s 492954 0 493010 800 6 la_data_out[109]
port 284 nsew signal output
rlabel metal2 s 155958 0 156014 800 6 la_data_out[10]
port 285 nsew signal output
rlabel metal2 s 496358 0 496414 800 6 la_data_out[110]
port 286 nsew signal output
rlabel metal2 s 499762 0 499818 800 6 la_data_out[111]
port 287 nsew signal output
rlabel metal2 s 503166 0 503222 800 6 la_data_out[112]
port 288 nsew signal output
rlabel metal2 s 506570 0 506626 800 6 la_data_out[113]
port 289 nsew signal output
rlabel metal2 s 509974 0 510030 800 6 la_data_out[114]
port 290 nsew signal output
rlabel metal2 s 513378 0 513434 800 6 la_data_out[115]
port 291 nsew signal output
rlabel metal2 s 516782 0 516838 800 6 la_data_out[116]
port 292 nsew signal output
rlabel metal2 s 520186 0 520242 800 6 la_data_out[117]
port 293 nsew signal output
rlabel metal2 s 523590 0 523646 800 6 la_data_out[118]
port 294 nsew signal output
rlabel metal2 s 526994 0 527050 800 6 la_data_out[119]
port 295 nsew signal output
rlabel metal2 s 159362 0 159418 800 6 la_data_out[11]
port 296 nsew signal output
rlabel metal2 s 530398 0 530454 800 6 la_data_out[120]
port 297 nsew signal output
rlabel metal2 s 533802 0 533858 800 6 la_data_out[121]
port 298 nsew signal output
rlabel metal2 s 537206 0 537262 800 6 la_data_out[122]
port 299 nsew signal output
rlabel metal2 s 540610 0 540666 800 6 la_data_out[123]
port 300 nsew signal output
rlabel metal2 s 544014 0 544070 800 6 la_data_out[124]
port 301 nsew signal output
rlabel metal2 s 547418 0 547474 800 6 la_data_out[125]
port 302 nsew signal output
rlabel metal2 s 550822 0 550878 800 6 la_data_out[126]
port 303 nsew signal output
rlabel metal2 s 554226 0 554282 800 6 la_data_out[127]
port 304 nsew signal output
rlabel metal2 s 162766 0 162822 800 6 la_data_out[12]
port 305 nsew signal output
rlabel metal2 s 166170 0 166226 800 6 la_data_out[13]
port 306 nsew signal output
rlabel metal2 s 169574 0 169630 800 6 la_data_out[14]
port 307 nsew signal output
rlabel metal2 s 172978 0 173034 800 6 la_data_out[15]
port 308 nsew signal output
rlabel metal2 s 176382 0 176438 800 6 la_data_out[16]
port 309 nsew signal output
rlabel metal2 s 179786 0 179842 800 6 la_data_out[17]
port 310 nsew signal output
rlabel metal2 s 183190 0 183246 800 6 la_data_out[18]
port 311 nsew signal output
rlabel metal2 s 186594 0 186650 800 6 la_data_out[19]
port 312 nsew signal output
rlabel metal2 s 125322 0 125378 800 6 la_data_out[1]
port 313 nsew signal output
rlabel metal2 s 189998 0 190054 800 6 la_data_out[20]
port 314 nsew signal output
rlabel metal2 s 193402 0 193458 800 6 la_data_out[21]
port 315 nsew signal output
rlabel metal2 s 196806 0 196862 800 6 la_data_out[22]
port 316 nsew signal output
rlabel metal2 s 200210 0 200266 800 6 la_data_out[23]
port 317 nsew signal output
rlabel metal2 s 203614 0 203670 800 6 la_data_out[24]
port 318 nsew signal output
rlabel metal2 s 207018 0 207074 800 6 la_data_out[25]
port 319 nsew signal output
rlabel metal2 s 210422 0 210478 800 6 la_data_out[26]
port 320 nsew signal output
rlabel metal2 s 213826 0 213882 800 6 la_data_out[27]
port 321 nsew signal output
rlabel metal2 s 217230 0 217286 800 6 la_data_out[28]
port 322 nsew signal output
rlabel metal2 s 220634 0 220690 800 6 la_data_out[29]
port 323 nsew signal output
rlabel metal2 s 128726 0 128782 800 6 la_data_out[2]
port 324 nsew signal output
rlabel metal2 s 224038 0 224094 800 6 la_data_out[30]
port 325 nsew signal output
rlabel metal2 s 227442 0 227498 800 6 la_data_out[31]
port 326 nsew signal output
rlabel metal2 s 230846 0 230902 800 6 la_data_out[32]
port 327 nsew signal output
rlabel metal2 s 234250 0 234306 800 6 la_data_out[33]
port 328 nsew signal output
rlabel metal2 s 237654 0 237710 800 6 la_data_out[34]
port 329 nsew signal output
rlabel metal2 s 241058 0 241114 800 6 la_data_out[35]
port 330 nsew signal output
rlabel metal2 s 244462 0 244518 800 6 la_data_out[36]
port 331 nsew signal output
rlabel metal2 s 247866 0 247922 800 6 la_data_out[37]
port 332 nsew signal output
rlabel metal2 s 251270 0 251326 800 6 la_data_out[38]
port 333 nsew signal output
rlabel metal2 s 254674 0 254730 800 6 la_data_out[39]
port 334 nsew signal output
rlabel metal2 s 132130 0 132186 800 6 la_data_out[3]
port 335 nsew signal output
rlabel metal2 s 258078 0 258134 800 6 la_data_out[40]
port 336 nsew signal output
rlabel metal2 s 261482 0 261538 800 6 la_data_out[41]
port 337 nsew signal output
rlabel metal2 s 264886 0 264942 800 6 la_data_out[42]
port 338 nsew signal output
rlabel metal2 s 268290 0 268346 800 6 la_data_out[43]
port 339 nsew signal output
rlabel metal2 s 271694 0 271750 800 6 la_data_out[44]
port 340 nsew signal output
rlabel metal2 s 275098 0 275154 800 6 la_data_out[45]
port 341 nsew signal output
rlabel metal2 s 278502 0 278558 800 6 la_data_out[46]
port 342 nsew signal output
rlabel metal2 s 281906 0 281962 800 6 la_data_out[47]
port 343 nsew signal output
rlabel metal2 s 285310 0 285366 800 6 la_data_out[48]
port 344 nsew signal output
rlabel metal2 s 288714 0 288770 800 6 la_data_out[49]
port 345 nsew signal output
rlabel metal2 s 135534 0 135590 800 6 la_data_out[4]
port 346 nsew signal output
rlabel metal2 s 292118 0 292174 800 6 la_data_out[50]
port 347 nsew signal output
rlabel metal2 s 295522 0 295578 800 6 la_data_out[51]
port 348 nsew signal output
rlabel metal2 s 298926 0 298982 800 6 la_data_out[52]
port 349 nsew signal output
rlabel metal2 s 302330 0 302386 800 6 la_data_out[53]
port 350 nsew signal output
rlabel metal2 s 305734 0 305790 800 6 la_data_out[54]
port 351 nsew signal output
rlabel metal2 s 309138 0 309194 800 6 la_data_out[55]
port 352 nsew signal output
rlabel metal2 s 312542 0 312598 800 6 la_data_out[56]
port 353 nsew signal output
rlabel metal2 s 315946 0 316002 800 6 la_data_out[57]
port 354 nsew signal output
rlabel metal2 s 319350 0 319406 800 6 la_data_out[58]
port 355 nsew signal output
rlabel metal2 s 322754 0 322810 800 6 la_data_out[59]
port 356 nsew signal output
rlabel metal2 s 138938 0 138994 800 6 la_data_out[5]
port 357 nsew signal output
rlabel metal2 s 326158 0 326214 800 6 la_data_out[60]
port 358 nsew signal output
rlabel metal2 s 329562 0 329618 800 6 la_data_out[61]
port 359 nsew signal output
rlabel metal2 s 332966 0 333022 800 6 la_data_out[62]
port 360 nsew signal output
rlabel metal2 s 336370 0 336426 800 6 la_data_out[63]
port 361 nsew signal output
rlabel metal2 s 339774 0 339830 800 6 la_data_out[64]
port 362 nsew signal output
rlabel metal2 s 343178 0 343234 800 6 la_data_out[65]
port 363 nsew signal output
rlabel metal2 s 346582 0 346638 800 6 la_data_out[66]
port 364 nsew signal output
rlabel metal2 s 349986 0 350042 800 6 la_data_out[67]
port 365 nsew signal output
rlabel metal2 s 353390 0 353446 800 6 la_data_out[68]
port 366 nsew signal output
rlabel metal2 s 356794 0 356850 800 6 la_data_out[69]
port 367 nsew signal output
rlabel metal2 s 142342 0 142398 800 6 la_data_out[6]
port 368 nsew signal output
rlabel metal2 s 360198 0 360254 800 6 la_data_out[70]
port 369 nsew signal output
rlabel metal2 s 363602 0 363658 800 6 la_data_out[71]
port 370 nsew signal output
rlabel metal2 s 367006 0 367062 800 6 la_data_out[72]
port 371 nsew signal output
rlabel metal2 s 370410 0 370466 800 6 la_data_out[73]
port 372 nsew signal output
rlabel metal2 s 373814 0 373870 800 6 la_data_out[74]
port 373 nsew signal output
rlabel metal2 s 377218 0 377274 800 6 la_data_out[75]
port 374 nsew signal output
rlabel metal2 s 380622 0 380678 800 6 la_data_out[76]
port 375 nsew signal output
rlabel metal2 s 384026 0 384082 800 6 la_data_out[77]
port 376 nsew signal output
rlabel metal2 s 387430 0 387486 800 6 la_data_out[78]
port 377 nsew signal output
rlabel metal2 s 390834 0 390890 800 6 la_data_out[79]
port 378 nsew signal output
rlabel metal2 s 145746 0 145802 800 6 la_data_out[7]
port 379 nsew signal output
rlabel metal2 s 394238 0 394294 800 6 la_data_out[80]
port 380 nsew signal output
rlabel metal2 s 397642 0 397698 800 6 la_data_out[81]
port 381 nsew signal output
rlabel metal2 s 401046 0 401102 800 6 la_data_out[82]
port 382 nsew signal output
rlabel metal2 s 404450 0 404506 800 6 la_data_out[83]
port 383 nsew signal output
rlabel metal2 s 407854 0 407910 800 6 la_data_out[84]
port 384 nsew signal output
rlabel metal2 s 411258 0 411314 800 6 la_data_out[85]
port 385 nsew signal output
rlabel metal2 s 414662 0 414718 800 6 la_data_out[86]
port 386 nsew signal output
rlabel metal2 s 418066 0 418122 800 6 la_data_out[87]
port 387 nsew signal output
rlabel metal2 s 421470 0 421526 800 6 la_data_out[88]
port 388 nsew signal output
rlabel metal2 s 424874 0 424930 800 6 la_data_out[89]
port 389 nsew signal output
rlabel metal2 s 149150 0 149206 800 6 la_data_out[8]
port 390 nsew signal output
rlabel metal2 s 428278 0 428334 800 6 la_data_out[90]
port 391 nsew signal output
rlabel metal2 s 431682 0 431738 800 6 la_data_out[91]
port 392 nsew signal output
rlabel metal2 s 435086 0 435142 800 6 la_data_out[92]
port 393 nsew signal output
rlabel metal2 s 438490 0 438546 800 6 la_data_out[93]
port 394 nsew signal output
rlabel metal2 s 441894 0 441950 800 6 la_data_out[94]
port 395 nsew signal output
rlabel metal2 s 445298 0 445354 800 6 la_data_out[95]
port 396 nsew signal output
rlabel metal2 s 448702 0 448758 800 6 la_data_out[96]
port 397 nsew signal output
rlabel metal2 s 452106 0 452162 800 6 la_data_out[97]
port 398 nsew signal output
rlabel metal2 s 455510 0 455566 800 6 la_data_out[98]
port 399 nsew signal output
rlabel metal2 s 458914 0 458970 800 6 la_data_out[99]
port 400 nsew signal output
rlabel metal2 s 152554 0 152610 800 6 la_data_out[9]
port 401 nsew signal output
rlabel metal2 s 123114 0 123170 800 6 la_oen[0]
port 402 nsew signal input
rlabel metal2 s 463514 0 463570 800 6 la_oen[100]
port 403 nsew signal input
rlabel metal2 s 466918 0 466974 800 6 la_oen[101]
port 404 nsew signal input
rlabel metal2 s 470322 0 470378 800 6 la_oen[102]
port 405 nsew signal input
rlabel metal2 s 473726 0 473782 800 6 la_oen[103]
port 406 nsew signal input
rlabel metal2 s 477130 0 477186 800 6 la_oen[104]
port 407 nsew signal input
rlabel metal2 s 480534 0 480590 800 6 la_oen[105]
port 408 nsew signal input
rlabel metal2 s 483938 0 483994 800 6 la_oen[106]
port 409 nsew signal input
rlabel metal2 s 487342 0 487398 800 6 la_oen[107]
port 410 nsew signal input
rlabel metal2 s 490746 0 490802 800 6 la_oen[108]
port 411 nsew signal input
rlabel metal2 s 494150 0 494206 800 6 la_oen[109]
port 412 nsew signal input
rlabel metal2 s 157154 0 157210 800 6 la_oen[10]
port 413 nsew signal input
rlabel metal2 s 497554 0 497610 800 6 la_oen[110]
port 414 nsew signal input
rlabel metal2 s 500958 0 501014 800 6 la_oen[111]
port 415 nsew signal input
rlabel metal2 s 504362 0 504418 800 6 la_oen[112]
port 416 nsew signal input
rlabel metal2 s 507766 0 507822 800 6 la_oen[113]
port 417 nsew signal input
rlabel metal2 s 511170 0 511226 800 6 la_oen[114]
port 418 nsew signal input
rlabel metal2 s 514574 0 514630 800 6 la_oen[115]
port 419 nsew signal input
rlabel metal2 s 517978 0 518034 800 6 la_oen[116]
port 420 nsew signal input
rlabel metal2 s 521382 0 521438 800 6 la_oen[117]
port 421 nsew signal input
rlabel metal2 s 524786 0 524842 800 6 la_oen[118]
port 422 nsew signal input
rlabel metal2 s 528190 0 528246 800 6 la_oen[119]
port 423 nsew signal input
rlabel metal2 s 160558 0 160614 800 6 la_oen[11]
port 424 nsew signal input
rlabel metal2 s 531594 0 531650 800 6 la_oen[120]
port 425 nsew signal input
rlabel metal2 s 534998 0 535054 800 6 la_oen[121]
port 426 nsew signal input
rlabel metal2 s 538402 0 538458 800 6 la_oen[122]
port 427 nsew signal input
rlabel metal2 s 541806 0 541862 800 6 la_oen[123]
port 428 nsew signal input
rlabel metal2 s 545210 0 545266 800 6 la_oen[124]
port 429 nsew signal input
rlabel metal2 s 548614 0 548670 800 6 la_oen[125]
port 430 nsew signal input
rlabel metal2 s 552018 0 552074 800 6 la_oen[126]
port 431 nsew signal input
rlabel metal2 s 555422 0 555478 800 6 la_oen[127]
port 432 nsew signal input
rlabel metal2 s 163962 0 164018 800 6 la_oen[12]
port 433 nsew signal input
rlabel metal2 s 167366 0 167422 800 6 la_oen[13]
port 434 nsew signal input
rlabel metal2 s 170770 0 170826 800 6 la_oen[14]
port 435 nsew signal input
rlabel metal2 s 174174 0 174230 800 6 la_oen[15]
port 436 nsew signal input
rlabel metal2 s 177578 0 177634 800 6 la_oen[16]
port 437 nsew signal input
rlabel metal2 s 180982 0 181038 800 6 la_oen[17]
port 438 nsew signal input
rlabel metal2 s 184386 0 184442 800 6 la_oen[18]
port 439 nsew signal input
rlabel metal2 s 187790 0 187846 800 6 la_oen[19]
port 440 nsew signal input
rlabel metal2 s 126518 0 126574 800 6 la_oen[1]
port 441 nsew signal input
rlabel metal2 s 191194 0 191250 800 6 la_oen[20]
port 442 nsew signal input
rlabel metal2 s 194598 0 194654 800 6 la_oen[21]
port 443 nsew signal input
rlabel metal2 s 198002 0 198058 800 6 la_oen[22]
port 444 nsew signal input
rlabel metal2 s 201406 0 201462 800 6 la_oen[23]
port 445 nsew signal input
rlabel metal2 s 204810 0 204866 800 6 la_oen[24]
port 446 nsew signal input
rlabel metal2 s 208214 0 208270 800 6 la_oen[25]
port 447 nsew signal input
rlabel metal2 s 211618 0 211674 800 6 la_oen[26]
port 448 nsew signal input
rlabel metal2 s 215022 0 215078 800 6 la_oen[27]
port 449 nsew signal input
rlabel metal2 s 218426 0 218482 800 6 la_oen[28]
port 450 nsew signal input
rlabel metal2 s 221830 0 221886 800 6 la_oen[29]
port 451 nsew signal input
rlabel metal2 s 129922 0 129978 800 6 la_oen[2]
port 452 nsew signal input
rlabel metal2 s 225234 0 225290 800 6 la_oen[30]
port 453 nsew signal input
rlabel metal2 s 228638 0 228694 800 6 la_oen[31]
port 454 nsew signal input
rlabel metal2 s 232042 0 232098 800 6 la_oen[32]
port 455 nsew signal input
rlabel metal2 s 235446 0 235502 800 6 la_oen[33]
port 456 nsew signal input
rlabel metal2 s 238850 0 238906 800 6 la_oen[34]
port 457 nsew signal input
rlabel metal2 s 242254 0 242310 800 6 la_oen[35]
port 458 nsew signal input
rlabel metal2 s 245658 0 245714 800 6 la_oen[36]
port 459 nsew signal input
rlabel metal2 s 249062 0 249118 800 6 la_oen[37]
port 460 nsew signal input
rlabel metal2 s 252466 0 252522 800 6 la_oen[38]
port 461 nsew signal input
rlabel metal2 s 255870 0 255926 800 6 la_oen[39]
port 462 nsew signal input
rlabel metal2 s 133326 0 133382 800 6 la_oen[3]
port 463 nsew signal input
rlabel metal2 s 259274 0 259330 800 6 la_oen[40]
port 464 nsew signal input
rlabel metal2 s 262678 0 262734 800 6 la_oen[41]
port 465 nsew signal input
rlabel metal2 s 266082 0 266138 800 6 la_oen[42]
port 466 nsew signal input
rlabel metal2 s 269486 0 269542 800 6 la_oen[43]
port 467 nsew signal input
rlabel metal2 s 272890 0 272946 800 6 la_oen[44]
port 468 nsew signal input
rlabel metal2 s 276294 0 276350 800 6 la_oen[45]
port 469 nsew signal input
rlabel metal2 s 279698 0 279754 800 6 la_oen[46]
port 470 nsew signal input
rlabel metal2 s 283102 0 283158 800 6 la_oen[47]
port 471 nsew signal input
rlabel metal2 s 286506 0 286562 800 6 la_oen[48]
port 472 nsew signal input
rlabel metal2 s 289910 0 289966 800 6 la_oen[49]
port 473 nsew signal input
rlabel metal2 s 136730 0 136786 800 6 la_oen[4]
port 474 nsew signal input
rlabel metal2 s 293314 0 293370 800 6 la_oen[50]
port 475 nsew signal input
rlabel metal2 s 296718 0 296774 800 6 la_oen[51]
port 476 nsew signal input
rlabel metal2 s 300122 0 300178 800 6 la_oen[52]
port 477 nsew signal input
rlabel metal2 s 303526 0 303582 800 6 la_oen[53]
port 478 nsew signal input
rlabel metal2 s 306930 0 306986 800 6 la_oen[54]
port 479 nsew signal input
rlabel metal2 s 310334 0 310390 800 6 la_oen[55]
port 480 nsew signal input
rlabel metal2 s 313738 0 313794 800 6 la_oen[56]
port 481 nsew signal input
rlabel metal2 s 317142 0 317198 800 6 la_oen[57]
port 482 nsew signal input
rlabel metal2 s 320546 0 320602 800 6 la_oen[58]
port 483 nsew signal input
rlabel metal2 s 323950 0 324006 800 6 la_oen[59]
port 484 nsew signal input
rlabel metal2 s 140134 0 140190 800 6 la_oen[5]
port 485 nsew signal input
rlabel metal2 s 327354 0 327410 800 6 la_oen[60]
port 486 nsew signal input
rlabel metal2 s 330758 0 330814 800 6 la_oen[61]
port 487 nsew signal input
rlabel metal2 s 334162 0 334218 800 6 la_oen[62]
port 488 nsew signal input
rlabel metal2 s 337566 0 337622 800 6 la_oen[63]
port 489 nsew signal input
rlabel metal2 s 340970 0 341026 800 6 la_oen[64]
port 490 nsew signal input
rlabel metal2 s 344374 0 344430 800 6 la_oen[65]
port 491 nsew signal input
rlabel metal2 s 347778 0 347834 800 6 la_oen[66]
port 492 nsew signal input
rlabel metal2 s 351182 0 351238 800 6 la_oen[67]
port 493 nsew signal input
rlabel metal2 s 354586 0 354642 800 6 la_oen[68]
port 494 nsew signal input
rlabel metal2 s 357990 0 358046 800 6 la_oen[69]
port 495 nsew signal input
rlabel metal2 s 143538 0 143594 800 6 la_oen[6]
port 496 nsew signal input
rlabel metal2 s 361394 0 361450 800 6 la_oen[70]
port 497 nsew signal input
rlabel metal2 s 364798 0 364854 800 6 la_oen[71]
port 498 nsew signal input
rlabel metal2 s 368202 0 368258 800 6 la_oen[72]
port 499 nsew signal input
rlabel metal2 s 371606 0 371662 800 6 la_oen[73]
port 500 nsew signal input
rlabel metal2 s 375010 0 375066 800 6 la_oen[74]
port 501 nsew signal input
rlabel metal2 s 378414 0 378470 800 6 la_oen[75]
port 502 nsew signal input
rlabel metal2 s 381818 0 381874 800 6 la_oen[76]
port 503 nsew signal input
rlabel metal2 s 385222 0 385278 800 6 la_oen[77]
port 504 nsew signal input
rlabel metal2 s 388626 0 388682 800 6 la_oen[78]
port 505 nsew signal input
rlabel metal2 s 392030 0 392086 800 6 la_oen[79]
port 506 nsew signal input
rlabel metal2 s 146942 0 146998 800 6 la_oen[7]
port 507 nsew signal input
rlabel metal2 s 395434 0 395490 800 6 la_oen[80]
port 508 nsew signal input
rlabel metal2 s 398838 0 398894 800 6 la_oen[81]
port 509 nsew signal input
rlabel metal2 s 402242 0 402298 800 6 la_oen[82]
port 510 nsew signal input
rlabel metal2 s 405646 0 405702 800 6 la_oen[83]
port 511 nsew signal input
rlabel metal2 s 409050 0 409106 800 6 la_oen[84]
port 512 nsew signal input
rlabel metal2 s 412454 0 412510 800 6 la_oen[85]
port 513 nsew signal input
rlabel metal2 s 415858 0 415914 800 6 la_oen[86]
port 514 nsew signal input
rlabel metal2 s 419262 0 419318 800 6 la_oen[87]
port 515 nsew signal input
rlabel metal2 s 422666 0 422722 800 6 la_oen[88]
port 516 nsew signal input
rlabel metal2 s 426070 0 426126 800 6 la_oen[89]
port 517 nsew signal input
rlabel metal2 s 150346 0 150402 800 6 la_oen[8]
port 518 nsew signal input
rlabel metal2 s 429474 0 429530 800 6 la_oen[90]
port 519 nsew signal input
rlabel metal2 s 432878 0 432934 800 6 la_oen[91]
port 520 nsew signal input
rlabel metal2 s 436282 0 436338 800 6 la_oen[92]
port 521 nsew signal input
rlabel metal2 s 439686 0 439742 800 6 la_oen[93]
port 522 nsew signal input
rlabel metal2 s 443090 0 443146 800 6 la_oen[94]
port 523 nsew signal input
rlabel metal2 s 446494 0 446550 800 6 la_oen[95]
port 524 nsew signal input
rlabel metal2 s 449898 0 449954 800 6 la_oen[96]
port 525 nsew signal input
rlabel metal2 s 453302 0 453358 800 6 la_oen[97]
port 526 nsew signal input
rlabel metal2 s 456706 0 456762 800 6 la_oen[98]
port 527 nsew signal input
rlabel metal2 s 460110 0 460166 800 6 la_oen[99]
port 528 nsew signal input
rlabel metal2 s 153750 0 153806 800 6 la_oen[9]
port 529 nsew signal input
rlabel metal2 s 556526 0 556582 800 6 user_clock2
port 530 nsew signal input
rlabel metal2 s 570 0 626 800 6 wb_clk_i
port 531 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wb_rst_i
port 532 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 wbs_ack_o
port 533 nsew signal output
rlabel metal2 s 7378 0 7434 800 6 wbs_adr_i[0]
port 534 nsew signal input
rlabel metal2 s 45926 0 45982 800 6 wbs_adr_i[10]
port 535 nsew signal input
rlabel metal2 s 49330 0 49386 800 6 wbs_adr_i[11]
port 536 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 wbs_adr_i[12]
port 537 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 wbs_adr_i[13]
port 538 nsew signal input
rlabel metal2 s 59542 0 59598 800 6 wbs_adr_i[14]
port 539 nsew signal input
rlabel metal2 s 62946 0 63002 800 6 wbs_adr_i[15]
port 540 nsew signal input
rlabel metal2 s 66350 0 66406 800 6 wbs_adr_i[16]
port 541 nsew signal input
rlabel metal2 s 69754 0 69810 800 6 wbs_adr_i[17]
port 542 nsew signal input
rlabel metal2 s 73158 0 73214 800 6 wbs_adr_i[18]
port 543 nsew signal input
rlabel metal2 s 76562 0 76618 800 6 wbs_adr_i[19]
port 544 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 wbs_adr_i[1]
port 545 nsew signal input
rlabel metal2 s 79966 0 80022 800 6 wbs_adr_i[20]
port 546 nsew signal input
rlabel metal2 s 83370 0 83426 800 6 wbs_adr_i[21]
port 547 nsew signal input
rlabel metal2 s 86774 0 86830 800 6 wbs_adr_i[22]
port 548 nsew signal input
rlabel metal2 s 90178 0 90234 800 6 wbs_adr_i[23]
port 549 nsew signal input
rlabel metal2 s 93582 0 93638 800 6 wbs_adr_i[24]
port 550 nsew signal input
rlabel metal2 s 96986 0 97042 800 6 wbs_adr_i[25]
port 551 nsew signal input
rlabel metal2 s 100390 0 100446 800 6 wbs_adr_i[26]
port 552 nsew signal input
rlabel metal2 s 103794 0 103850 800 6 wbs_adr_i[27]
port 553 nsew signal input
rlabel metal2 s 107198 0 107254 800 6 wbs_adr_i[28]
port 554 nsew signal input
rlabel metal2 s 110602 0 110658 800 6 wbs_adr_i[29]
port 555 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 wbs_adr_i[2]
port 556 nsew signal input
rlabel metal2 s 114006 0 114062 800 6 wbs_adr_i[30]
port 557 nsew signal input
rlabel metal2 s 117410 0 117466 800 6 wbs_adr_i[31]
port 558 nsew signal input
rlabel metal2 s 20994 0 21050 800 6 wbs_adr_i[3]
port 559 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 wbs_adr_i[4]
port 560 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 wbs_adr_i[5]
port 561 nsew signal input
rlabel metal2 s 32310 0 32366 800 6 wbs_adr_i[6]
port 562 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 wbs_adr_i[7]
port 563 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 wbs_adr_i[8]
port 564 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 wbs_adr_i[9]
port 565 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 wbs_cyc_i
port 566 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_dat_i[0]
port 567 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 wbs_dat_i[10]
port 568 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 wbs_dat_i[11]
port 569 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 wbs_dat_i[12]
port 570 nsew signal input
rlabel metal2 s 57242 0 57298 800 6 wbs_dat_i[13]
port 571 nsew signal input
rlabel metal2 s 60646 0 60702 800 6 wbs_dat_i[14]
port 572 nsew signal input
rlabel metal2 s 64050 0 64106 800 6 wbs_dat_i[15]
port 573 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 wbs_dat_i[16]
port 574 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 wbs_dat_i[17]
port 575 nsew signal input
rlabel metal2 s 74262 0 74318 800 6 wbs_dat_i[18]
port 576 nsew signal input
rlabel metal2 s 77666 0 77722 800 6 wbs_dat_i[19]
port 577 nsew signal input
rlabel metal2 s 12990 0 13046 800 6 wbs_dat_i[1]
port 578 nsew signal input
rlabel metal2 s 81070 0 81126 800 6 wbs_dat_i[20]
port 579 nsew signal input
rlabel metal2 s 84474 0 84530 800 6 wbs_dat_i[21]
port 580 nsew signal input
rlabel metal2 s 87878 0 87934 800 6 wbs_dat_i[22]
port 581 nsew signal input
rlabel metal2 s 91282 0 91338 800 6 wbs_dat_i[23]
port 582 nsew signal input
rlabel metal2 s 94686 0 94742 800 6 wbs_dat_i[24]
port 583 nsew signal input
rlabel metal2 s 98090 0 98146 800 6 wbs_dat_i[25]
port 584 nsew signal input
rlabel metal2 s 101494 0 101550 800 6 wbs_dat_i[26]
port 585 nsew signal input
rlabel metal2 s 104898 0 104954 800 6 wbs_dat_i[27]
port 586 nsew signal input
rlabel metal2 s 108302 0 108358 800 6 wbs_dat_i[28]
port 587 nsew signal input
rlabel metal2 s 111706 0 111762 800 6 wbs_dat_i[29]
port 588 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 wbs_dat_i[2]
port 589 nsew signal input
rlabel metal2 s 115110 0 115166 800 6 wbs_dat_i[30]
port 590 nsew signal input
rlabel metal2 s 118514 0 118570 800 6 wbs_dat_i[31]
port 591 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 wbs_dat_i[3]
port 592 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 wbs_dat_i[4]
port 593 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 wbs_dat_i[5]
port 594 nsew signal input
rlabel metal2 s 33414 0 33470 800 6 wbs_dat_i[6]
port 595 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 wbs_dat_i[7]
port 596 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 wbs_dat_i[8]
port 597 nsew signal input
rlabel metal2 s 43626 0 43682 800 6 wbs_dat_i[9]
port 598 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_dat_o[0]
port 599 nsew signal output
rlabel metal2 s 48226 0 48282 800 6 wbs_dat_o[10]
port 600 nsew signal output
rlabel metal2 s 51630 0 51686 800 6 wbs_dat_o[11]
port 601 nsew signal output
rlabel metal2 s 55034 0 55090 800 6 wbs_dat_o[12]
port 602 nsew signal output
rlabel metal2 s 58438 0 58494 800 6 wbs_dat_o[13]
port 603 nsew signal output
rlabel metal2 s 61842 0 61898 800 6 wbs_dat_o[14]
port 604 nsew signal output
rlabel metal2 s 65246 0 65302 800 6 wbs_dat_o[15]
port 605 nsew signal output
rlabel metal2 s 68650 0 68706 800 6 wbs_dat_o[16]
port 606 nsew signal output
rlabel metal2 s 72054 0 72110 800 6 wbs_dat_o[17]
port 607 nsew signal output
rlabel metal2 s 75458 0 75514 800 6 wbs_dat_o[18]
port 608 nsew signal output
rlabel metal2 s 78862 0 78918 800 6 wbs_dat_o[19]
port 609 nsew signal output
rlabel metal2 s 14186 0 14242 800 6 wbs_dat_o[1]
port 610 nsew signal output
rlabel metal2 s 82266 0 82322 800 6 wbs_dat_o[20]
port 611 nsew signal output
rlabel metal2 s 85670 0 85726 800 6 wbs_dat_o[21]
port 612 nsew signal output
rlabel metal2 s 89074 0 89130 800 6 wbs_dat_o[22]
port 613 nsew signal output
rlabel metal2 s 92478 0 92534 800 6 wbs_dat_o[23]
port 614 nsew signal output
rlabel metal2 s 95882 0 95938 800 6 wbs_dat_o[24]
port 615 nsew signal output
rlabel metal2 s 99286 0 99342 800 6 wbs_dat_o[25]
port 616 nsew signal output
rlabel metal2 s 102690 0 102746 800 6 wbs_dat_o[26]
port 617 nsew signal output
rlabel metal2 s 106094 0 106150 800 6 wbs_dat_o[27]
port 618 nsew signal output
rlabel metal2 s 109498 0 109554 800 6 wbs_dat_o[28]
port 619 nsew signal output
rlabel metal2 s 112902 0 112958 800 6 wbs_dat_o[29]
port 620 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 wbs_dat_o[2]
port 621 nsew signal output
rlabel metal2 s 116306 0 116362 800 6 wbs_dat_o[30]
port 622 nsew signal output
rlabel metal2 s 119710 0 119766 800 6 wbs_dat_o[31]
port 623 nsew signal output
rlabel metal2 s 23202 0 23258 800 6 wbs_dat_o[3]
port 624 nsew signal output
rlabel metal2 s 27802 0 27858 800 6 wbs_dat_o[4]
port 625 nsew signal output
rlabel metal2 s 31206 0 31262 800 6 wbs_dat_o[5]
port 626 nsew signal output
rlabel metal2 s 34610 0 34666 800 6 wbs_dat_o[6]
port 627 nsew signal output
rlabel metal2 s 38014 0 38070 800 6 wbs_dat_o[7]
port 628 nsew signal output
rlabel metal2 s 41418 0 41474 800 6 wbs_dat_o[8]
port 629 nsew signal output
rlabel metal2 s 44822 0 44878 800 6 wbs_dat_o[9]
port 630 nsew signal output
rlabel metal2 s 10782 0 10838 800 6 wbs_sel_i[0]
port 631 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 wbs_sel_i[1]
port 632 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 wbs_sel_i[2]
port 633 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 wbs_sel_i[3]
port 634 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 wbs_stb_i
port 635 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wbs_we_i
port 636 nsew signal input
rlabel metal4 s 557168 2128 557488 681680 6 VPWR
port 637 nsew power bidirectional
rlabel metal4 s 526448 2128 526768 681680 6 VPWR
port 638 nsew power bidirectional
rlabel metal4 s 495728 2128 496048 681680 6 VPWR
port 639 nsew power bidirectional
rlabel metal4 s 465008 2128 465328 681680 6 VPWR
port 640 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 681680 6 VPWR
port 641 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 681680 6 VPWR
port 642 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 681680 6 VPWR
port 643 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 681680 6 VPWR
port 644 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 681680 6 VPWR
port 645 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 681680 6 VPWR
port 646 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 681680 6 VPWR
port 647 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 681680 6 VPWR
port 648 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 681680 6 VPWR
port 649 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 681680 6 VPWR
port 650 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 681680 6 VPWR
port 651 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 681680 6 VPWR
port 652 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 681680 6 VPWR
port 653 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 681680 6 VPWR
port 654 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 681680 6 VPWR
port 655 nsew power bidirectional
rlabel metal4 s 541808 2128 542128 681680 6 VGND
port 656 nsew ground bidirectional
rlabel metal4 s 511088 2128 511408 681680 6 VGND
port 657 nsew ground bidirectional
rlabel metal4 s 480368 2128 480688 681680 6 VGND
port 658 nsew ground bidirectional
rlabel metal4 s 449648 2128 449968 681680 6 VGND
port 659 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 681680 6 VGND
port 660 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 681680 6 VGND
port 661 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 681680 6 VGND
port 662 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 681680 6 VGND
port 663 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 681680 6 VGND
port 664 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 681680 6 VGND
port 665 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 681680 6 VGND
port 666 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 681680 6 VGND
port 667 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 681680 6 VGND
port 668 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 681680 6 VGND
port 669 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 681680 6 VGND
port 670 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 681680 6 VGND
port 671 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 681680 6 VGND
port 672 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 681680 6 VGND
port 673 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 564000 684000
string LEFview TRUE
<< end >>

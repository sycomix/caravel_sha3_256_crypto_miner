VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 2840.000 BY 3440.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2836.000 155.760 2840.000 156.360 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2732.950 3436.000 2733.230 3440.000 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2756.870 3436.000 2757.150 3440.000 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1719.760 4.000 1720.360 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2836.000 1406.280 2840.000 1406.880 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2819.890 0.000 2820.170 4.000 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2101.920 4.000 2102.520 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2836.000 1719.080 2840.000 1719.680 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2836.000 2031.880 2840.000 2032.480 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2484.080 4.000 2484.680 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2836.000 2344.680 2840.000 2345.280 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2709.490 3436.000 2709.770 3440.000 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2780.330 3436.000 2780.610 3440.000 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2866.240 4.000 2866.840 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2825.410 0.000 2825.690 4.000 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2804.250 3436.000 2804.530 3440.000 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2827.710 3436.000 2827.990 3440.000 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3248.400 4.000 3249.000 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2831.390 0.000 2831.670 4.000 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2836.000 2657.480 2840.000 2658.080 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2836.910 0.000 2837.190 4.000 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2836.000 2970.280 2840.000 2970.880 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.120 4.000 191.720 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2836.000 3283.080 2840.000 3283.680 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2836.000 467.880 2840.000 468.480 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 573.280 4.000 573.880 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 955.440 4.000 956.040 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2836.000 780.680 2840.000 781.280 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1337.600 4.000 1338.200 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2836.000 1093.480 2840.000 1094.080 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2813.910 0.000 2814.190 4.000 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 3436.000 11.870 3440.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 3436.000 721.650 3440.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.210 3436.000 792.490 3440.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.510 3436.000 863.790 3440.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 934.350 3436.000 934.630 3440.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1005.190 3436.000 1005.470 3440.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.490 3436.000 1076.770 3440.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1147.330 3436.000 1147.610 3440.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1218.170 3436.000 1218.450 3440.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1289.470 3436.000 1289.750 3440.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1360.310 3436.000 1360.590 3440.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 3436.000 82.710 3440.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1431.610 3436.000 1431.890 3440.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1502.450 3436.000 1502.730 3440.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1573.290 3436.000 1573.570 3440.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1644.590 3436.000 1644.870 3440.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1715.430 3436.000 1715.710 3440.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1786.270 3436.000 1786.550 3440.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1857.570 3436.000 1857.850 3440.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1928.410 3436.000 1928.690 3440.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1999.250 3436.000 1999.530 3440.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2070.550 3436.000 2070.830 3440.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 3436.000 153.550 3440.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2141.390 3436.000 2141.670 3440.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2212.230 3436.000 2212.510 3440.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2283.530 3436.000 2283.810 3440.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2354.370 3436.000 2354.650 3440.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2425.210 3436.000 2425.490 3440.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2496.510 3436.000 2496.790 3440.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2567.350 3436.000 2567.630 3440.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2638.190 3436.000 2638.470 3440.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 3436.000 224.850 3440.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 3436.000 295.690 3440.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.250 3436.000 366.530 3440.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.550 3436.000 437.830 3440.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.390 3436.000 508.670 3440.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.230 3436.000 579.510 3440.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.530 3436.000 650.810 3440.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 3436.000 35.330 3440.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.830 3436.000 745.110 3440.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 816.130 3436.000 816.410 3440.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.970 3436.000 887.250 3440.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 958.270 3436.000 958.550 3440.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1029.110 3436.000 1029.390 3440.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1099.950 3436.000 1100.230 3440.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1171.250 3436.000 1171.530 3440.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1242.090 3436.000 1242.370 3440.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1312.930 3436.000 1313.210 3440.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1384.230 3436.000 1384.510 3440.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 3436.000 106.170 3440.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1455.070 3436.000 1455.350 3440.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1525.910 3436.000 1526.190 3440.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1597.210 3436.000 1597.490 3440.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1668.050 3436.000 1668.330 3440.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1738.890 3436.000 1739.170 3440.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1810.190 3436.000 1810.470 3440.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1881.030 3436.000 1881.310 3440.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1951.870 3436.000 1952.150 3440.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2023.170 3436.000 2023.450 3440.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2094.010 3436.000 2094.290 3440.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 3436.000 177.470 3440.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2164.850 3436.000 2165.130 3440.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2236.150 3436.000 2236.430 3440.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2306.990 3436.000 2307.270 3440.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2378.290 3436.000 2378.570 3440.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2449.130 3436.000 2449.410 3440.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2519.970 3436.000 2520.250 3440.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2591.270 3436.000 2591.550 3440.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2662.110 3436.000 2662.390 3440.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 3436.000 248.310 3440.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 3436.000 319.150 3440.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.170 3436.000 390.450 3440.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.010 3436.000 461.290 3440.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.850 3436.000 532.130 3440.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.150 3436.000 603.430 3440.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.990 3436.000 674.270 3440.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 3436.000 58.790 3440.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.750 3436.000 769.030 3440.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.590 3436.000 839.870 3440.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 910.890 3436.000 911.170 3440.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 981.730 3436.000 982.010 3440.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1052.570 3436.000 1052.850 3440.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1123.870 3436.000 1124.150 3440.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1194.710 3436.000 1194.990 3440.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1265.550 3436.000 1265.830 3440.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1336.850 3436.000 1337.130 3440.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1407.690 3436.000 1407.970 3440.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 3436.000 130.090 3440.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1478.530 3436.000 1478.810 3440.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1549.830 3436.000 1550.110 3440.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1620.670 3436.000 1620.950 3440.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1691.510 3436.000 1691.790 3440.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1762.810 3436.000 1763.090 3440.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1833.650 3436.000 1833.930 3440.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1904.950 3436.000 1905.230 3440.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1975.790 3436.000 1976.070 3440.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2046.630 3436.000 2046.910 3440.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2117.930 3436.000 2118.210 3440.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 3436.000 200.930 3440.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2188.770 3436.000 2189.050 3440.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2259.610 3436.000 2259.890 3440.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2330.910 3436.000 2331.190 3440.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2401.750 3436.000 2402.030 3440.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2472.590 3436.000 2472.870 3440.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2543.890 3436.000 2544.170 3440.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2614.730 3436.000 2615.010 3440.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2685.570 3436.000 2685.850 3440.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 3436.000 271.770 3440.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 3436.000 343.070 3440.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.630 3436.000 413.910 3440.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.930 3436.000 485.210 3440.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.770 3436.000 556.050 3440.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.610 3436.000 626.890 3440.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.910 3436.000 698.190 3440.000 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.590 0.000 609.870 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2327.230 0.000 2327.510 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2344.710 0.000 2344.990 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2361.730 0.000 2362.010 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2378.750 0.000 2379.030 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2396.230 0.000 2396.510 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2413.250 0.000 2413.530 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2430.270 0.000 2430.550 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2447.750 0.000 2448.030 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2464.770 0.000 2465.050 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2481.790 0.000 2482.070 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.170 0.000 781.450 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2499.270 0.000 2499.550 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2516.290 0.000 2516.570 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2533.310 0.000 2533.590 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2550.790 0.000 2551.070 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2567.810 0.000 2568.090 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2584.830 0.000 2585.110 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2602.310 0.000 2602.590 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2619.330 0.000 2619.610 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2636.350 0.000 2636.630 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2653.830 0.000 2654.110 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.650 0.000 798.930 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2670.850 0.000 2671.130 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2687.870 0.000 2688.150 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2705.350 0.000 2705.630 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2722.370 0.000 2722.650 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2739.390 0.000 2739.670 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2756.870 0.000 2757.150 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2773.890 0.000 2774.170 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2790.910 0.000 2791.190 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.670 0.000 815.950 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 832.690 0.000 832.970 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.170 0.000 850.450 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 867.190 0.000 867.470 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 884.210 0.000 884.490 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.690 0.000 901.970 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.710 0.000 918.990 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 935.730 0.000 936.010 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.610 0.000 626.890 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.210 0.000 953.490 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 970.230 0.000 970.510 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 987.250 0.000 987.530 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1004.730 0.000 1005.010 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1021.750 0.000 1022.030 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1039.230 0.000 1039.510 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.250 0.000 1056.530 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1073.270 0.000 1073.550 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.750 0.000 1091.030 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.770 0.000 1108.050 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 0.000 644.370 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1124.790 0.000 1125.070 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1142.270 0.000 1142.550 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1159.290 0.000 1159.570 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1176.310 0.000 1176.590 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1193.790 0.000 1194.070 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1210.810 0.000 1211.090 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1227.830 0.000 1228.110 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1245.310 0.000 1245.590 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1262.330 0.000 1262.610 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1279.350 0.000 1279.630 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.110 0.000 661.390 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1296.830 0.000 1297.110 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1313.850 0.000 1314.130 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1330.870 0.000 1331.150 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1348.350 0.000 1348.630 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1365.370 0.000 1365.650 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1382.390 0.000 1382.670 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1399.870 0.000 1400.150 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1416.890 0.000 1417.170 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1433.910 0.000 1434.190 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1451.390 0.000 1451.670 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.130 0.000 678.410 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.410 0.000 1468.690 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1485.430 0.000 1485.710 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1502.910 0.000 1503.190 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1519.930 0.000 1520.210 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1536.950 0.000 1537.230 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1554.430 0.000 1554.710 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1571.450 0.000 1571.730 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1588.470 0.000 1588.750 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1605.950 0.000 1606.230 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1622.970 0.000 1623.250 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 0.000 695.890 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1640.450 0.000 1640.730 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1657.470 0.000 1657.750 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1674.490 0.000 1674.770 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1691.970 0.000 1692.250 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1708.990 0.000 1709.270 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1726.010 0.000 1726.290 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1743.490 0.000 1743.770 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1760.510 0.000 1760.790 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1777.530 0.000 1777.810 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1795.010 0.000 1795.290 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.630 0.000 712.910 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1812.030 0.000 1812.310 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1829.050 0.000 1829.330 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1846.530 0.000 1846.810 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1863.550 0.000 1863.830 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1880.570 0.000 1880.850 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1898.050 0.000 1898.330 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1915.070 0.000 1915.350 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1932.090 0.000 1932.370 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1949.570 0.000 1949.850 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1966.590 0.000 1966.870 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.650 0.000 729.930 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1983.610 0.000 1983.890 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2001.090 0.000 2001.370 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2018.110 0.000 2018.390 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2035.130 0.000 2035.410 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2052.610 0.000 2052.890 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2069.630 0.000 2069.910 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2086.650 0.000 2086.930 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2104.130 0.000 2104.410 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2121.150 0.000 2121.430 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2138.170 0.000 2138.450 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 0.000 747.410 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2155.650 0.000 2155.930 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2172.670 0.000 2172.950 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2189.690 0.000 2189.970 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2207.170 0.000 2207.450 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2224.190 0.000 2224.470 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2241.670 0.000 2241.950 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2258.690 0.000 2258.970 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2275.710 0.000 2275.990 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2293.190 0.000 2293.470 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2310.210 0.000 2310.490 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.150 0.000 764.430 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.110 0.000 615.390 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2333.210 0.000 2333.490 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2350.230 0.000 2350.510 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2367.250 0.000 2367.530 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2384.730 0.000 2385.010 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2401.750 0.000 2402.030 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2418.770 0.000 2419.050 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2436.250 0.000 2436.530 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2453.270 0.000 2453.550 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2470.290 0.000 2470.570 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2487.770 0.000 2488.050 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.150 0.000 787.430 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2504.790 0.000 2505.070 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2521.810 0.000 2522.090 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2539.290 0.000 2539.570 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2556.310 0.000 2556.590 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2573.330 0.000 2573.610 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2590.810 0.000 2591.090 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2607.830 0.000 2608.110 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2624.850 0.000 2625.130 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2642.330 0.000 2642.610 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2659.350 0.000 2659.630 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.170 0.000 804.450 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2676.830 0.000 2677.110 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2693.850 0.000 2694.130 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2710.870 0.000 2711.150 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2728.350 0.000 2728.630 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2745.370 0.000 2745.650 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2762.390 0.000 2762.670 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2779.870 0.000 2780.150 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2796.890 0.000 2797.170 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.650 0.000 821.930 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 838.670 0.000 838.950 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.690 0.000 855.970 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 873.170 0.000 873.450 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 890.190 0.000 890.470 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.210 0.000 907.490 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.690 0.000 924.970 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 941.710 0.000 941.990 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.590 0.000 632.870 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 958.730 0.000 959.010 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.210 0.000 976.490 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 993.230 0.000 993.510 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1010.250 0.000 1010.530 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1027.730 0.000 1028.010 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1044.750 0.000 1045.030 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1061.770 0.000 1062.050 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1079.250 0.000 1079.530 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1096.270 0.000 1096.550 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1113.290 0.000 1113.570 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.610 0.000 649.890 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1130.770 0.000 1131.050 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1147.790 0.000 1148.070 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1164.810 0.000 1165.090 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1182.290 0.000 1182.570 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1199.310 0.000 1199.590 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1216.330 0.000 1216.610 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1233.810 0.000 1234.090 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1250.830 0.000 1251.110 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1267.850 0.000 1268.130 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1285.330 0.000 1285.610 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.630 0.000 666.910 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1302.350 0.000 1302.630 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1319.370 0.000 1319.650 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1336.850 0.000 1337.130 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1353.870 0.000 1354.150 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1370.890 0.000 1371.170 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1388.370 0.000 1388.650 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1405.390 0.000 1405.670 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1422.870 0.000 1423.150 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1439.890 0.000 1440.170 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1456.910 0.000 1457.190 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.110 0.000 684.390 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1474.390 0.000 1474.670 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1491.410 0.000 1491.690 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1508.430 0.000 1508.710 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1525.910 0.000 1526.190 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1542.930 0.000 1543.210 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1559.950 0.000 1560.230 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1577.430 0.000 1577.710 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1594.450 0.000 1594.730 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1611.470 0.000 1611.750 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1628.950 0.000 1629.230 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.130 0.000 701.410 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1645.970 0.000 1646.250 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1662.990 0.000 1663.270 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1680.470 0.000 1680.750 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1697.490 0.000 1697.770 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1714.510 0.000 1714.790 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1731.990 0.000 1732.270 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1749.010 0.000 1749.290 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1766.030 0.000 1766.310 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1783.510 0.000 1783.790 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1800.530 0.000 1800.810 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.150 0.000 718.430 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1817.550 0.000 1817.830 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1835.030 0.000 1835.310 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1852.050 0.000 1852.330 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1869.070 0.000 1869.350 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1886.550 0.000 1886.830 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1903.570 0.000 1903.850 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1920.590 0.000 1920.870 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1938.070 0.000 1938.350 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1955.090 0.000 1955.370 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1972.110 0.000 1972.390 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.630 0.000 735.910 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1989.590 0.000 1989.870 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2006.610 0.000 2006.890 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2023.630 0.000 2023.910 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2041.110 0.000 2041.390 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2058.130 0.000 2058.410 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2075.610 0.000 2075.890 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2092.630 0.000 2092.910 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2109.650 0.000 2109.930 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2127.130 0.000 2127.410 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2144.150 0.000 2144.430 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.650 0.000 752.930 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2161.170 0.000 2161.450 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2178.650 0.000 2178.930 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2195.670 0.000 2195.950 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2212.690 0.000 2212.970 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.170 0.000 2230.450 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2247.190 0.000 2247.470 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2264.210 0.000 2264.490 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2281.690 0.000 2281.970 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2298.710 0.000 2298.990 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2315.730 0.000 2316.010 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.670 0.000 769.950 4.000 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.090 0.000 621.370 4.000 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2338.730 0.000 2339.010 4.000 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2355.750 0.000 2356.030 4.000 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2373.230 0.000 2373.510 4.000 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2390.250 0.000 2390.530 4.000 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2407.270 0.000 2407.550 4.000 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2424.750 0.000 2425.030 4.000 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2441.770 0.000 2442.050 4.000 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2459.250 0.000 2459.530 4.000 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2476.270 0.000 2476.550 4.000 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2493.290 0.000 2493.570 4.000 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.670 0.000 792.950 4.000 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2510.770 0.000 2511.050 4.000 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2527.790 0.000 2528.070 4.000 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2544.810 0.000 2545.090 4.000 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2562.290 0.000 2562.570 4.000 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2579.310 0.000 2579.590 4.000 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2596.330 0.000 2596.610 4.000 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2613.810 0.000 2614.090 4.000 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2630.830 0.000 2631.110 4.000 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2647.850 0.000 2648.130 4.000 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2665.330 0.000 2665.610 4.000 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.150 0.000 810.430 4.000 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2682.350 0.000 2682.630 4.000 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2699.370 0.000 2699.650 4.000 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2716.850 0.000 2717.130 4.000 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2733.870 0.000 2734.150 4.000 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2750.890 0.000 2751.170 4.000 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2768.370 0.000 2768.650 4.000 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2785.390 0.000 2785.670 4.000 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2802.410 0.000 2802.690 4.000 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.170 0.000 827.450 4.000 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 844.190 0.000 844.470 4.000 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.670 0.000 861.950 4.000 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 878.690 0.000 878.970 4.000 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.710 0.000 895.990 4.000 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 913.190 0.000 913.470 4.000 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.210 0.000 930.490 4.000 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 947.230 0.000 947.510 4.000 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.110 0.000 638.390 4.000 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 964.710 0.000 964.990 4.000 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 981.730 0.000 982.010 4.000 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.750 0.000 999.030 4.000 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1016.230 0.000 1016.510 4.000 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.250 0.000 1033.530 4.000 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1050.270 0.000 1050.550 4.000 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1067.750 0.000 1068.030 4.000 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1084.770 0.000 1085.050 4.000 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1101.790 0.000 1102.070 4.000 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1119.270 0.000 1119.550 4.000 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.590 0.000 655.870 4.000 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1136.290 0.000 1136.570 4.000 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1153.310 0.000 1153.590 4.000 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1170.790 0.000 1171.070 4.000 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1187.810 0.000 1188.090 4.000 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1204.830 0.000 1205.110 4.000 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1222.310 0.000 1222.590 4.000 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1239.330 0.000 1239.610 4.000 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1256.810 0.000 1257.090 4.000 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1273.830 0.000 1274.110 4.000 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1290.850 0.000 1291.130 4.000 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.610 0.000 672.890 4.000 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1308.330 0.000 1308.610 4.000 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1325.350 0.000 1325.630 4.000 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1342.370 0.000 1342.650 4.000 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1359.850 0.000 1360.130 4.000 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1376.870 0.000 1377.150 4.000 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1393.890 0.000 1394.170 4.000 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1411.370 0.000 1411.650 4.000 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1428.390 0.000 1428.670 4.000 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1445.410 0.000 1445.690 4.000 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1462.890 0.000 1463.170 4.000 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.630 0.000 689.910 4.000 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1479.910 0.000 1480.190 4.000 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1496.930 0.000 1497.210 4.000 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1514.410 0.000 1514.690 4.000 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1531.430 0.000 1531.710 4.000 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1548.450 0.000 1548.730 4.000 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1565.930 0.000 1566.210 4.000 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1582.950 0.000 1583.230 4.000 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1599.970 0.000 1600.250 4.000 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1617.450 0.000 1617.730 4.000 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1634.470 0.000 1634.750 4.000 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.110 0.000 707.390 4.000 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.490 0.000 1651.770 4.000 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1668.970 0.000 1669.250 4.000 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1685.990 0.000 1686.270 4.000 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1703.010 0.000 1703.290 4.000 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1720.490 0.000 1720.770 4.000 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1737.510 0.000 1737.790 4.000 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1754.530 0.000 1754.810 4.000 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1772.010 0.000 1772.290 4.000 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1789.030 0.000 1789.310 4.000 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1806.050 0.000 1806.330 4.000 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.130 0.000 724.410 4.000 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1823.530 0.000 1823.810 4.000 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1840.550 0.000 1840.830 4.000 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1858.030 0.000 1858.310 4.000 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1875.050 0.000 1875.330 4.000 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1892.070 0.000 1892.350 4.000 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1909.550 0.000 1909.830 4.000 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1926.570 0.000 1926.850 4.000 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1943.590 0.000 1943.870 4.000 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1961.070 0.000 1961.350 4.000 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1978.090 0.000 1978.370 4.000 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.150 0.000 741.430 4.000 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1995.110 0.000 1995.390 4.000 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2012.590 0.000 2012.870 4.000 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2029.610 0.000 2029.890 4.000 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2046.630 0.000 2046.910 4.000 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2064.110 0.000 2064.390 4.000 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2081.130 0.000 2081.410 4.000 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2098.150 0.000 2098.430 4.000 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2115.630 0.000 2115.910 4.000 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2132.650 0.000 2132.930 4.000 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2149.670 0.000 2149.950 4.000 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.630 0.000 758.910 4.000 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2167.150 0.000 2167.430 4.000 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2184.170 0.000 2184.450 4.000 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2201.190 0.000 2201.470 4.000 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2218.670 0.000 2218.950 4.000 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2235.690 0.000 2235.970 4.000 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2252.710 0.000 2252.990 4.000 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2270.190 0.000 2270.470 4.000 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2287.210 0.000 2287.490 4.000 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2304.230 0.000 2304.510 4.000 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2321.710 0.000 2321.990 4.000 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.650 0.000 775.930 4.000 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2808.390 0.000 2808.670 4.000 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.470 0.000 231.750 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.950 0.000 249.230 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.970 0.000 266.250 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.990 0.000 283.270 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.470 0.000 300.750 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 0.000 317.770 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.510 0.000 334.790 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 0.000 352.270 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.010 0.000 369.290 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.030 0.000 386.310 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.510 0.000 403.790 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.530 0.000 420.810 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 0.000 438.290 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.030 0.000 455.310 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.050 0.000 472.330 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 0.000 489.810 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.550 0.000 506.830 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.570 0.000 523.850 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 0.000 541.330 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.070 0.000 558.350 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.090 0.000 575.370 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 0.000 592.850 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 0.000 128.710 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 0.000 146.190 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.930 0.000 163.210 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 0.000 180.230 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 0.000 197.710 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 0.000 214.730 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 0.000 20.150 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 0.000 237.730 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 0.000 272.230 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.970 0.000 289.250 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.470 0.000 323.750 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.490 0.000 340.770 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.990 0.000 375.270 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 0.000 392.290 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 0.000 409.310 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.510 0.000 426.790 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.530 0.000 443.810 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 0.000 460.830 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.030 0.000 478.310 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.050 0.000 495.330 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 0.000 512.350 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.550 0.000 529.830 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.570 0.000 546.850 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 0.000 563.870 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.070 0.000 581.350 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.090 0.000 598.370 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 0.000 134.690 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.430 0.000 220.710 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 0.000 243.250 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.450 0.000 260.730 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 0.000 277.750 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 0.000 294.770 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 0.000 312.250 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.990 0.000 329.270 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.010 0.000 346.290 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 0.000 363.770 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.510 0.000 380.790 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.530 0.000 397.810 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.010 0.000 415.290 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.030 0.000 432.310 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.050 0.000 449.330 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.530 0.000 466.810 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.550 0.000 483.830 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.570 0.000 500.850 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.050 0.000 518.330 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.070 0.000 535.350 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.090 0.000 552.370 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.570 0.000 569.850 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.590 0.000 586.870 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.610 0.000 603.890 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.930 0.000 140.210 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 0.000 157.690 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 0.000 174.710 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 0.000 191.730 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 0.000 209.210 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.950 0.000 226.230 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.650 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 0.000 123.190 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 4.000 ;
    END
  END wbs_we_i
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2785.840 10.640 2787.440 3427.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2632.240 10.640 2633.840 3427.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2478.640 10.640 2480.240 3427.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2325.040 10.640 2326.640 3427.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2171.440 10.640 2173.040 3427.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2017.840 10.640 2019.440 3427.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1864.240 10.640 1865.840 3427.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 3427.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 3427.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 3427.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 3427.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 3427.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 3427.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 3427.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 3427.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 3427.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 3427.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 3427.440 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 3427.440 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2709.040 10.640 2710.640 3427.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2555.440 10.640 2557.040 3427.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2401.840 10.640 2403.440 3427.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2248.240 10.640 2249.840 3427.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2094.640 10.640 2096.240 3427.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1941.040 10.640 1942.640 3427.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 3427.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 3427.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 3427.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 3427.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 3427.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 3427.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 3427.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 3427.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 3427.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 3427.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 3427.440 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 3427.440 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2834.060 3427.285 ;
      LAYER met1 ;
        RECT 0.070 6.160 2834.060 3427.440 ;
      LAYER met2 ;
        RECT 0.100 3435.720 11.310 3436.000 ;
        RECT 12.150 3435.720 34.770 3436.000 ;
        RECT 35.610 3435.720 58.230 3436.000 ;
        RECT 59.070 3435.720 82.150 3436.000 ;
        RECT 82.990 3435.720 105.610 3436.000 ;
        RECT 106.450 3435.720 129.530 3436.000 ;
        RECT 130.370 3435.720 152.990 3436.000 ;
        RECT 153.830 3435.720 176.910 3436.000 ;
        RECT 177.750 3435.720 200.370 3436.000 ;
        RECT 201.210 3435.720 224.290 3436.000 ;
        RECT 225.130 3435.720 247.750 3436.000 ;
        RECT 248.590 3435.720 271.210 3436.000 ;
        RECT 272.050 3435.720 295.130 3436.000 ;
        RECT 295.970 3435.720 318.590 3436.000 ;
        RECT 319.430 3435.720 342.510 3436.000 ;
        RECT 343.350 3435.720 365.970 3436.000 ;
        RECT 366.810 3435.720 389.890 3436.000 ;
        RECT 390.730 3435.720 413.350 3436.000 ;
        RECT 414.190 3435.720 437.270 3436.000 ;
        RECT 438.110 3435.720 460.730 3436.000 ;
        RECT 461.570 3435.720 484.650 3436.000 ;
        RECT 485.490 3435.720 508.110 3436.000 ;
        RECT 508.950 3435.720 531.570 3436.000 ;
        RECT 532.410 3435.720 555.490 3436.000 ;
        RECT 556.330 3435.720 578.950 3436.000 ;
        RECT 579.790 3435.720 602.870 3436.000 ;
        RECT 603.710 3435.720 626.330 3436.000 ;
        RECT 627.170 3435.720 650.250 3436.000 ;
        RECT 651.090 3435.720 673.710 3436.000 ;
        RECT 674.550 3435.720 697.630 3436.000 ;
        RECT 698.470 3435.720 721.090 3436.000 ;
        RECT 721.930 3435.720 744.550 3436.000 ;
        RECT 745.390 3435.720 768.470 3436.000 ;
        RECT 769.310 3435.720 791.930 3436.000 ;
        RECT 792.770 3435.720 815.850 3436.000 ;
        RECT 816.690 3435.720 839.310 3436.000 ;
        RECT 840.150 3435.720 863.230 3436.000 ;
        RECT 864.070 3435.720 886.690 3436.000 ;
        RECT 887.530 3435.720 910.610 3436.000 ;
        RECT 911.450 3435.720 934.070 3436.000 ;
        RECT 934.910 3435.720 957.990 3436.000 ;
        RECT 958.830 3435.720 981.450 3436.000 ;
        RECT 982.290 3435.720 1004.910 3436.000 ;
        RECT 1005.750 3435.720 1028.830 3436.000 ;
        RECT 1029.670 3435.720 1052.290 3436.000 ;
        RECT 1053.130 3435.720 1076.210 3436.000 ;
        RECT 1077.050 3435.720 1099.670 3436.000 ;
        RECT 1100.510 3435.720 1123.590 3436.000 ;
        RECT 1124.430 3435.720 1147.050 3436.000 ;
        RECT 1147.890 3435.720 1170.970 3436.000 ;
        RECT 1171.810 3435.720 1194.430 3436.000 ;
        RECT 1195.270 3435.720 1217.890 3436.000 ;
        RECT 1218.730 3435.720 1241.810 3436.000 ;
        RECT 1242.650 3435.720 1265.270 3436.000 ;
        RECT 1266.110 3435.720 1289.190 3436.000 ;
        RECT 1290.030 3435.720 1312.650 3436.000 ;
        RECT 1313.490 3435.720 1336.570 3436.000 ;
        RECT 1337.410 3435.720 1360.030 3436.000 ;
        RECT 1360.870 3435.720 1383.950 3436.000 ;
        RECT 1384.790 3435.720 1407.410 3436.000 ;
        RECT 1408.250 3435.720 1431.330 3436.000 ;
        RECT 1432.170 3435.720 1454.790 3436.000 ;
        RECT 1455.630 3435.720 1478.250 3436.000 ;
        RECT 1479.090 3435.720 1502.170 3436.000 ;
        RECT 1503.010 3435.720 1525.630 3436.000 ;
        RECT 1526.470 3435.720 1549.550 3436.000 ;
        RECT 1550.390 3435.720 1573.010 3436.000 ;
        RECT 1573.850 3435.720 1596.930 3436.000 ;
        RECT 1597.770 3435.720 1620.390 3436.000 ;
        RECT 1621.230 3435.720 1644.310 3436.000 ;
        RECT 1645.150 3435.720 1667.770 3436.000 ;
        RECT 1668.610 3435.720 1691.230 3436.000 ;
        RECT 1692.070 3435.720 1715.150 3436.000 ;
        RECT 1715.990 3435.720 1738.610 3436.000 ;
        RECT 1739.450 3435.720 1762.530 3436.000 ;
        RECT 1763.370 3435.720 1785.990 3436.000 ;
        RECT 1786.830 3435.720 1809.910 3436.000 ;
        RECT 1810.750 3435.720 1833.370 3436.000 ;
        RECT 1834.210 3435.720 1857.290 3436.000 ;
        RECT 1858.130 3435.720 1880.750 3436.000 ;
        RECT 1881.590 3435.720 1904.670 3436.000 ;
        RECT 1905.510 3435.720 1928.130 3436.000 ;
        RECT 1928.970 3435.720 1951.590 3436.000 ;
        RECT 1952.430 3435.720 1975.510 3436.000 ;
        RECT 1976.350 3435.720 1998.970 3436.000 ;
        RECT 1999.810 3435.720 2022.890 3436.000 ;
        RECT 2023.730 3435.720 2046.350 3436.000 ;
        RECT 2047.190 3435.720 2070.270 3436.000 ;
        RECT 2071.110 3435.720 2093.730 3436.000 ;
        RECT 2094.570 3435.720 2117.650 3436.000 ;
        RECT 2118.490 3435.720 2141.110 3436.000 ;
        RECT 2141.950 3435.720 2164.570 3436.000 ;
        RECT 2165.410 3435.720 2188.490 3436.000 ;
        RECT 2189.330 3435.720 2211.950 3436.000 ;
        RECT 2212.790 3435.720 2235.870 3436.000 ;
        RECT 2236.710 3435.720 2259.330 3436.000 ;
        RECT 2260.170 3435.720 2283.250 3436.000 ;
        RECT 2284.090 3435.720 2306.710 3436.000 ;
        RECT 2307.550 3435.720 2330.630 3436.000 ;
        RECT 2331.470 3435.720 2354.090 3436.000 ;
        RECT 2354.930 3435.720 2378.010 3436.000 ;
        RECT 2378.850 3435.720 2401.470 3436.000 ;
        RECT 2402.310 3435.720 2424.930 3436.000 ;
        RECT 2425.770 3435.720 2448.850 3436.000 ;
        RECT 2449.690 3435.720 2472.310 3436.000 ;
        RECT 2473.150 3435.720 2496.230 3436.000 ;
        RECT 2497.070 3435.720 2519.690 3436.000 ;
        RECT 2520.530 3435.720 2543.610 3436.000 ;
        RECT 2544.450 3435.720 2567.070 3436.000 ;
        RECT 2567.910 3435.720 2590.990 3436.000 ;
        RECT 2591.830 3435.720 2614.450 3436.000 ;
        RECT 2615.290 3435.720 2637.910 3436.000 ;
        RECT 2638.750 3435.720 2661.830 3436.000 ;
        RECT 2662.670 3435.720 2685.290 3436.000 ;
        RECT 2686.130 3435.720 2709.210 3436.000 ;
        RECT 2710.050 3435.720 2732.670 3436.000 ;
        RECT 2733.510 3435.720 2756.590 3436.000 ;
        RECT 2757.430 3435.720 2780.050 3436.000 ;
        RECT 2780.890 3435.720 2803.970 3436.000 ;
        RECT 2804.810 3435.720 2808.670 3436.000 ;
        RECT 0.100 4.280 2808.670 3435.720 ;
        RECT 0.100 4.000 2.570 4.280 ;
        RECT 3.410 4.000 8.090 4.280 ;
        RECT 8.930 4.000 13.610 4.280 ;
        RECT 14.450 4.000 19.590 4.280 ;
        RECT 20.430 4.000 25.110 4.280 ;
        RECT 25.950 4.000 31.090 4.280 ;
        RECT 31.930 4.000 36.610 4.280 ;
        RECT 37.450 4.000 42.590 4.280 ;
        RECT 43.430 4.000 48.110 4.280 ;
        RECT 48.950 4.000 54.090 4.280 ;
        RECT 54.930 4.000 59.610 4.280 ;
        RECT 60.450 4.000 65.130 4.280 ;
        RECT 65.970 4.000 71.110 4.280 ;
        RECT 71.950 4.000 76.630 4.280 ;
        RECT 77.470 4.000 82.610 4.280 ;
        RECT 83.450 4.000 88.130 4.280 ;
        RECT 88.970 4.000 94.110 4.280 ;
        RECT 94.950 4.000 99.630 4.280 ;
        RECT 100.470 4.000 105.610 4.280 ;
        RECT 106.450 4.000 111.130 4.280 ;
        RECT 111.970 4.000 116.650 4.280 ;
        RECT 117.490 4.000 122.630 4.280 ;
        RECT 123.470 4.000 128.150 4.280 ;
        RECT 128.990 4.000 134.130 4.280 ;
        RECT 134.970 4.000 139.650 4.280 ;
        RECT 140.490 4.000 145.630 4.280 ;
        RECT 146.470 4.000 151.150 4.280 ;
        RECT 151.990 4.000 157.130 4.280 ;
        RECT 157.970 4.000 162.650 4.280 ;
        RECT 163.490 4.000 168.170 4.280 ;
        RECT 169.010 4.000 174.150 4.280 ;
        RECT 174.990 4.000 179.670 4.280 ;
        RECT 180.510 4.000 185.650 4.280 ;
        RECT 186.490 4.000 191.170 4.280 ;
        RECT 192.010 4.000 197.150 4.280 ;
        RECT 197.990 4.000 202.670 4.280 ;
        RECT 203.510 4.000 208.650 4.280 ;
        RECT 209.490 4.000 214.170 4.280 ;
        RECT 215.010 4.000 220.150 4.280 ;
        RECT 220.990 4.000 225.670 4.280 ;
        RECT 226.510 4.000 231.190 4.280 ;
        RECT 232.030 4.000 237.170 4.280 ;
        RECT 238.010 4.000 242.690 4.280 ;
        RECT 243.530 4.000 248.670 4.280 ;
        RECT 249.510 4.000 254.190 4.280 ;
        RECT 255.030 4.000 260.170 4.280 ;
        RECT 261.010 4.000 265.690 4.280 ;
        RECT 266.530 4.000 271.670 4.280 ;
        RECT 272.510 4.000 277.190 4.280 ;
        RECT 278.030 4.000 282.710 4.280 ;
        RECT 283.550 4.000 288.690 4.280 ;
        RECT 289.530 4.000 294.210 4.280 ;
        RECT 295.050 4.000 300.190 4.280 ;
        RECT 301.030 4.000 305.710 4.280 ;
        RECT 306.550 4.000 311.690 4.280 ;
        RECT 312.530 4.000 317.210 4.280 ;
        RECT 318.050 4.000 323.190 4.280 ;
        RECT 324.030 4.000 328.710 4.280 ;
        RECT 329.550 4.000 334.230 4.280 ;
        RECT 335.070 4.000 340.210 4.280 ;
        RECT 341.050 4.000 345.730 4.280 ;
        RECT 346.570 4.000 351.710 4.280 ;
        RECT 352.550 4.000 357.230 4.280 ;
        RECT 358.070 4.000 363.210 4.280 ;
        RECT 364.050 4.000 368.730 4.280 ;
        RECT 369.570 4.000 374.710 4.280 ;
        RECT 375.550 4.000 380.230 4.280 ;
        RECT 381.070 4.000 385.750 4.280 ;
        RECT 386.590 4.000 391.730 4.280 ;
        RECT 392.570 4.000 397.250 4.280 ;
        RECT 398.090 4.000 403.230 4.280 ;
        RECT 404.070 4.000 408.750 4.280 ;
        RECT 409.590 4.000 414.730 4.280 ;
        RECT 415.570 4.000 420.250 4.280 ;
        RECT 421.090 4.000 426.230 4.280 ;
        RECT 427.070 4.000 431.750 4.280 ;
        RECT 432.590 4.000 437.730 4.280 ;
        RECT 438.570 4.000 443.250 4.280 ;
        RECT 444.090 4.000 448.770 4.280 ;
        RECT 449.610 4.000 454.750 4.280 ;
        RECT 455.590 4.000 460.270 4.280 ;
        RECT 461.110 4.000 466.250 4.280 ;
        RECT 467.090 4.000 471.770 4.280 ;
        RECT 472.610 4.000 477.750 4.280 ;
        RECT 478.590 4.000 483.270 4.280 ;
        RECT 484.110 4.000 489.250 4.280 ;
        RECT 490.090 4.000 494.770 4.280 ;
        RECT 495.610 4.000 500.290 4.280 ;
        RECT 501.130 4.000 506.270 4.280 ;
        RECT 507.110 4.000 511.790 4.280 ;
        RECT 512.630 4.000 517.770 4.280 ;
        RECT 518.610 4.000 523.290 4.280 ;
        RECT 524.130 4.000 529.270 4.280 ;
        RECT 530.110 4.000 534.790 4.280 ;
        RECT 535.630 4.000 540.770 4.280 ;
        RECT 541.610 4.000 546.290 4.280 ;
        RECT 547.130 4.000 551.810 4.280 ;
        RECT 552.650 4.000 557.790 4.280 ;
        RECT 558.630 4.000 563.310 4.280 ;
        RECT 564.150 4.000 569.290 4.280 ;
        RECT 570.130 4.000 574.810 4.280 ;
        RECT 575.650 4.000 580.790 4.280 ;
        RECT 581.630 4.000 586.310 4.280 ;
        RECT 587.150 4.000 592.290 4.280 ;
        RECT 593.130 4.000 597.810 4.280 ;
        RECT 598.650 4.000 603.330 4.280 ;
        RECT 604.170 4.000 609.310 4.280 ;
        RECT 610.150 4.000 614.830 4.280 ;
        RECT 615.670 4.000 620.810 4.280 ;
        RECT 621.650 4.000 626.330 4.280 ;
        RECT 627.170 4.000 632.310 4.280 ;
        RECT 633.150 4.000 637.830 4.280 ;
        RECT 638.670 4.000 643.810 4.280 ;
        RECT 644.650 4.000 649.330 4.280 ;
        RECT 650.170 4.000 655.310 4.280 ;
        RECT 656.150 4.000 660.830 4.280 ;
        RECT 661.670 4.000 666.350 4.280 ;
        RECT 667.190 4.000 672.330 4.280 ;
        RECT 673.170 4.000 677.850 4.280 ;
        RECT 678.690 4.000 683.830 4.280 ;
        RECT 684.670 4.000 689.350 4.280 ;
        RECT 690.190 4.000 695.330 4.280 ;
        RECT 696.170 4.000 700.850 4.280 ;
        RECT 701.690 4.000 706.830 4.280 ;
        RECT 707.670 4.000 712.350 4.280 ;
        RECT 713.190 4.000 717.870 4.280 ;
        RECT 718.710 4.000 723.850 4.280 ;
        RECT 724.690 4.000 729.370 4.280 ;
        RECT 730.210 4.000 735.350 4.280 ;
        RECT 736.190 4.000 740.870 4.280 ;
        RECT 741.710 4.000 746.850 4.280 ;
        RECT 747.690 4.000 752.370 4.280 ;
        RECT 753.210 4.000 758.350 4.280 ;
        RECT 759.190 4.000 763.870 4.280 ;
        RECT 764.710 4.000 769.390 4.280 ;
        RECT 770.230 4.000 775.370 4.280 ;
        RECT 776.210 4.000 780.890 4.280 ;
        RECT 781.730 4.000 786.870 4.280 ;
        RECT 787.710 4.000 792.390 4.280 ;
        RECT 793.230 4.000 798.370 4.280 ;
        RECT 799.210 4.000 803.890 4.280 ;
        RECT 804.730 4.000 809.870 4.280 ;
        RECT 810.710 4.000 815.390 4.280 ;
        RECT 816.230 4.000 821.370 4.280 ;
        RECT 822.210 4.000 826.890 4.280 ;
        RECT 827.730 4.000 832.410 4.280 ;
        RECT 833.250 4.000 838.390 4.280 ;
        RECT 839.230 4.000 843.910 4.280 ;
        RECT 844.750 4.000 849.890 4.280 ;
        RECT 850.730 4.000 855.410 4.280 ;
        RECT 856.250 4.000 861.390 4.280 ;
        RECT 862.230 4.000 866.910 4.280 ;
        RECT 867.750 4.000 872.890 4.280 ;
        RECT 873.730 4.000 878.410 4.280 ;
        RECT 879.250 4.000 883.930 4.280 ;
        RECT 884.770 4.000 889.910 4.280 ;
        RECT 890.750 4.000 895.430 4.280 ;
        RECT 896.270 4.000 901.410 4.280 ;
        RECT 902.250 4.000 906.930 4.280 ;
        RECT 907.770 4.000 912.910 4.280 ;
        RECT 913.750 4.000 918.430 4.280 ;
        RECT 919.270 4.000 924.410 4.280 ;
        RECT 925.250 4.000 929.930 4.280 ;
        RECT 930.770 4.000 935.450 4.280 ;
        RECT 936.290 4.000 941.430 4.280 ;
        RECT 942.270 4.000 946.950 4.280 ;
        RECT 947.790 4.000 952.930 4.280 ;
        RECT 953.770 4.000 958.450 4.280 ;
        RECT 959.290 4.000 964.430 4.280 ;
        RECT 965.270 4.000 969.950 4.280 ;
        RECT 970.790 4.000 975.930 4.280 ;
        RECT 976.770 4.000 981.450 4.280 ;
        RECT 982.290 4.000 986.970 4.280 ;
        RECT 987.810 4.000 992.950 4.280 ;
        RECT 993.790 4.000 998.470 4.280 ;
        RECT 999.310 4.000 1004.450 4.280 ;
        RECT 1005.290 4.000 1009.970 4.280 ;
        RECT 1010.810 4.000 1015.950 4.280 ;
        RECT 1016.790 4.000 1021.470 4.280 ;
        RECT 1022.310 4.000 1027.450 4.280 ;
        RECT 1028.290 4.000 1032.970 4.280 ;
        RECT 1033.810 4.000 1038.950 4.280 ;
        RECT 1039.790 4.000 1044.470 4.280 ;
        RECT 1045.310 4.000 1049.990 4.280 ;
        RECT 1050.830 4.000 1055.970 4.280 ;
        RECT 1056.810 4.000 1061.490 4.280 ;
        RECT 1062.330 4.000 1067.470 4.280 ;
        RECT 1068.310 4.000 1072.990 4.280 ;
        RECT 1073.830 4.000 1078.970 4.280 ;
        RECT 1079.810 4.000 1084.490 4.280 ;
        RECT 1085.330 4.000 1090.470 4.280 ;
        RECT 1091.310 4.000 1095.990 4.280 ;
        RECT 1096.830 4.000 1101.510 4.280 ;
        RECT 1102.350 4.000 1107.490 4.280 ;
        RECT 1108.330 4.000 1113.010 4.280 ;
        RECT 1113.850 4.000 1118.990 4.280 ;
        RECT 1119.830 4.000 1124.510 4.280 ;
        RECT 1125.350 4.000 1130.490 4.280 ;
        RECT 1131.330 4.000 1136.010 4.280 ;
        RECT 1136.850 4.000 1141.990 4.280 ;
        RECT 1142.830 4.000 1147.510 4.280 ;
        RECT 1148.350 4.000 1153.030 4.280 ;
        RECT 1153.870 4.000 1159.010 4.280 ;
        RECT 1159.850 4.000 1164.530 4.280 ;
        RECT 1165.370 4.000 1170.510 4.280 ;
        RECT 1171.350 4.000 1176.030 4.280 ;
        RECT 1176.870 4.000 1182.010 4.280 ;
        RECT 1182.850 4.000 1187.530 4.280 ;
        RECT 1188.370 4.000 1193.510 4.280 ;
        RECT 1194.350 4.000 1199.030 4.280 ;
        RECT 1199.870 4.000 1204.550 4.280 ;
        RECT 1205.390 4.000 1210.530 4.280 ;
        RECT 1211.370 4.000 1216.050 4.280 ;
        RECT 1216.890 4.000 1222.030 4.280 ;
        RECT 1222.870 4.000 1227.550 4.280 ;
        RECT 1228.390 4.000 1233.530 4.280 ;
        RECT 1234.370 4.000 1239.050 4.280 ;
        RECT 1239.890 4.000 1245.030 4.280 ;
        RECT 1245.870 4.000 1250.550 4.280 ;
        RECT 1251.390 4.000 1256.530 4.280 ;
        RECT 1257.370 4.000 1262.050 4.280 ;
        RECT 1262.890 4.000 1267.570 4.280 ;
        RECT 1268.410 4.000 1273.550 4.280 ;
        RECT 1274.390 4.000 1279.070 4.280 ;
        RECT 1279.910 4.000 1285.050 4.280 ;
        RECT 1285.890 4.000 1290.570 4.280 ;
        RECT 1291.410 4.000 1296.550 4.280 ;
        RECT 1297.390 4.000 1302.070 4.280 ;
        RECT 1302.910 4.000 1308.050 4.280 ;
        RECT 1308.890 4.000 1313.570 4.280 ;
        RECT 1314.410 4.000 1319.090 4.280 ;
        RECT 1319.930 4.000 1325.070 4.280 ;
        RECT 1325.910 4.000 1330.590 4.280 ;
        RECT 1331.430 4.000 1336.570 4.280 ;
        RECT 1337.410 4.000 1342.090 4.280 ;
        RECT 1342.930 4.000 1348.070 4.280 ;
        RECT 1348.910 4.000 1353.590 4.280 ;
        RECT 1354.430 4.000 1359.570 4.280 ;
        RECT 1360.410 4.000 1365.090 4.280 ;
        RECT 1365.930 4.000 1370.610 4.280 ;
        RECT 1371.450 4.000 1376.590 4.280 ;
        RECT 1377.430 4.000 1382.110 4.280 ;
        RECT 1382.950 4.000 1388.090 4.280 ;
        RECT 1388.930 4.000 1393.610 4.280 ;
        RECT 1394.450 4.000 1399.590 4.280 ;
        RECT 1400.430 4.000 1405.110 4.280 ;
        RECT 1405.950 4.000 1411.090 4.280 ;
        RECT 1411.930 4.000 1416.610 4.280 ;
        RECT 1417.450 4.000 1422.590 4.280 ;
        RECT 1423.430 4.000 1428.110 4.280 ;
        RECT 1428.950 4.000 1433.630 4.280 ;
        RECT 1434.470 4.000 1439.610 4.280 ;
        RECT 1440.450 4.000 1445.130 4.280 ;
        RECT 1445.970 4.000 1451.110 4.280 ;
        RECT 1451.950 4.000 1456.630 4.280 ;
        RECT 1457.470 4.000 1462.610 4.280 ;
        RECT 1463.450 4.000 1468.130 4.280 ;
        RECT 1468.970 4.000 1474.110 4.280 ;
        RECT 1474.950 4.000 1479.630 4.280 ;
        RECT 1480.470 4.000 1485.150 4.280 ;
        RECT 1485.990 4.000 1491.130 4.280 ;
        RECT 1491.970 4.000 1496.650 4.280 ;
        RECT 1497.490 4.000 1502.630 4.280 ;
        RECT 1503.470 4.000 1508.150 4.280 ;
        RECT 1508.990 4.000 1514.130 4.280 ;
        RECT 1514.970 4.000 1519.650 4.280 ;
        RECT 1520.490 4.000 1525.630 4.280 ;
        RECT 1526.470 4.000 1531.150 4.280 ;
        RECT 1531.990 4.000 1536.670 4.280 ;
        RECT 1537.510 4.000 1542.650 4.280 ;
        RECT 1543.490 4.000 1548.170 4.280 ;
        RECT 1549.010 4.000 1554.150 4.280 ;
        RECT 1554.990 4.000 1559.670 4.280 ;
        RECT 1560.510 4.000 1565.650 4.280 ;
        RECT 1566.490 4.000 1571.170 4.280 ;
        RECT 1572.010 4.000 1577.150 4.280 ;
        RECT 1577.990 4.000 1582.670 4.280 ;
        RECT 1583.510 4.000 1588.190 4.280 ;
        RECT 1589.030 4.000 1594.170 4.280 ;
        RECT 1595.010 4.000 1599.690 4.280 ;
        RECT 1600.530 4.000 1605.670 4.280 ;
        RECT 1606.510 4.000 1611.190 4.280 ;
        RECT 1612.030 4.000 1617.170 4.280 ;
        RECT 1618.010 4.000 1622.690 4.280 ;
        RECT 1623.530 4.000 1628.670 4.280 ;
        RECT 1629.510 4.000 1634.190 4.280 ;
        RECT 1635.030 4.000 1640.170 4.280 ;
        RECT 1641.010 4.000 1645.690 4.280 ;
        RECT 1646.530 4.000 1651.210 4.280 ;
        RECT 1652.050 4.000 1657.190 4.280 ;
        RECT 1658.030 4.000 1662.710 4.280 ;
        RECT 1663.550 4.000 1668.690 4.280 ;
        RECT 1669.530 4.000 1674.210 4.280 ;
        RECT 1675.050 4.000 1680.190 4.280 ;
        RECT 1681.030 4.000 1685.710 4.280 ;
        RECT 1686.550 4.000 1691.690 4.280 ;
        RECT 1692.530 4.000 1697.210 4.280 ;
        RECT 1698.050 4.000 1702.730 4.280 ;
        RECT 1703.570 4.000 1708.710 4.280 ;
        RECT 1709.550 4.000 1714.230 4.280 ;
        RECT 1715.070 4.000 1720.210 4.280 ;
        RECT 1721.050 4.000 1725.730 4.280 ;
        RECT 1726.570 4.000 1731.710 4.280 ;
        RECT 1732.550 4.000 1737.230 4.280 ;
        RECT 1738.070 4.000 1743.210 4.280 ;
        RECT 1744.050 4.000 1748.730 4.280 ;
        RECT 1749.570 4.000 1754.250 4.280 ;
        RECT 1755.090 4.000 1760.230 4.280 ;
        RECT 1761.070 4.000 1765.750 4.280 ;
        RECT 1766.590 4.000 1771.730 4.280 ;
        RECT 1772.570 4.000 1777.250 4.280 ;
        RECT 1778.090 4.000 1783.230 4.280 ;
        RECT 1784.070 4.000 1788.750 4.280 ;
        RECT 1789.590 4.000 1794.730 4.280 ;
        RECT 1795.570 4.000 1800.250 4.280 ;
        RECT 1801.090 4.000 1805.770 4.280 ;
        RECT 1806.610 4.000 1811.750 4.280 ;
        RECT 1812.590 4.000 1817.270 4.280 ;
        RECT 1818.110 4.000 1823.250 4.280 ;
        RECT 1824.090 4.000 1828.770 4.280 ;
        RECT 1829.610 4.000 1834.750 4.280 ;
        RECT 1835.590 4.000 1840.270 4.280 ;
        RECT 1841.110 4.000 1846.250 4.280 ;
        RECT 1847.090 4.000 1851.770 4.280 ;
        RECT 1852.610 4.000 1857.750 4.280 ;
        RECT 1858.590 4.000 1863.270 4.280 ;
        RECT 1864.110 4.000 1868.790 4.280 ;
        RECT 1869.630 4.000 1874.770 4.280 ;
        RECT 1875.610 4.000 1880.290 4.280 ;
        RECT 1881.130 4.000 1886.270 4.280 ;
        RECT 1887.110 4.000 1891.790 4.280 ;
        RECT 1892.630 4.000 1897.770 4.280 ;
        RECT 1898.610 4.000 1903.290 4.280 ;
        RECT 1904.130 4.000 1909.270 4.280 ;
        RECT 1910.110 4.000 1914.790 4.280 ;
        RECT 1915.630 4.000 1920.310 4.280 ;
        RECT 1921.150 4.000 1926.290 4.280 ;
        RECT 1927.130 4.000 1931.810 4.280 ;
        RECT 1932.650 4.000 1937.790 4.280 ;
        RECT 1938.630 4.000 1943.310 4.280 ;
        RECT 1944.150 4.000 1949.290 4.280 ;
        RECT 1950.130 4.000 1954.810 4.280 ;
        RECT 1955.650 4.000 1960.790 4.280 ;
        RECT 1961.630 4.000 1966.310 4.280 ;
        RECT 1967.150 4.000 1971.830 4.280 ;
        RECT 1972.670 4.000 1977.810 4.280 ;
        RECT 1978.650 4.000 1983.330 4.280 ;
        RECT 1984.170 4.000 1989.310 4.280 ;
        RECT 1990.150 4.000 1994.830 4.280 ;
        RECT 1995.670 4.000 2000.810 4.280 ;
        RECT 2001.650 4.000 2006.330 4.280 ;
        RECT 2007.170 4.000 2012.310 4.280 ;
        RECT 2013.150 4.000 2017.830 4.280 ;
        RECT 2018.670 4.000 2023.350 4.280 ;
        RECT 2024.190 4.000 2029.330 4.280 ;
        RECT 2030.170 4.000 2034.850 4.280 ;
        RECT 2035.690 4.000 2040.830 4.280 ;
        RECT 2041.670 4.000 2046.350 4.280 ;
        RECT 2047.190 4.000 2052.330 4.280 ;
        RECT 2053.170 4.000 2057.850 4.280 ;
        RECT 2058.690 4.000 2063.830 4.280 ;
        RECT 2064.670 4.000 2069.350 4.280 ;
        RECT 2070.190 4.000 2075.330 4.280 ;
        RECT 2076.170 4.000 2080.850 4.280 ;
        RECT 2081.690 4.000 2086.370 4.280 ;
        RECT 2087.210 4.000 2092.350 4.280 ;
        RECT 2093.190 4.000 2097.870 4.280 ;
        RECT 2098.710 4.000 2103.850 4.280 ;
        RECT 2104.690 4.000 2109.370 4.280 ;
        RECT 2110.210 4.000 2115.350 4.280 ;
        RECT 2116.190 4.000 2120.870 4.280 ;
        RECT 2121.710 4.000 2126.850 4.280 ;
        RECT 2127.690 4.000 2132.370 4.280 ;
        RECT 2133.210 4.000 2137.890 4.280 ;
        RECT 2138.730 4.000 2143.870 4.280 ;
        RECT 2144.710 4.000 2149.390 4.280 ;
        RECT 2150.230 4.000 2155.370 4.280 ;
        RECT 2156.210 4.000 2160.890 4.280 ;
        RECT 2161.730 4.000 2166.870 4.280 ;
        RECT 2167.710 4.000 2172.390 4.280 ;
        RECT 2173.230 4.000 2178.370 4.280 ;
        RECT 2179.210 4.000 2183.890 4.280 ;
        RECT 2184.730 4.000 2189.410 4.280 ;
        RECT 2190.250 4.000 2195.390 4.280 ;
        RECT 2196.230 4.000 2200.910 4.280 ;
        RECT 2201.750 4.000 2206.890 4.280 ;
        RECT 2207.730 4.000 2212.410 4.280 ;
        RECT 2213.250 4.000 2218.390 4.280 ;
        RECT 2219.230 4.000 2223.910 4.280 ;
        RECT 2224.750 4.000 2229.890 4.280 ;
        RECT 2230.730 4.000 2235.410 4.280 ;
        RECT 2236.250 4.000 2241.390 4.280 ;
        RECT 2242.230 4.000 2246.910 4.280 ;
        RECT 2247.750 4.000 2252.430 4.280 ;
        RECT 2253.270 4.000 2258.410 4.280 ;
        RECT 2259.250 4.000 2263.930 4.280 ;
        RECT 2264.770 4.000 2269.910 4.280 ;
        RECT 2270.750 4.000 2275.430 4.280 ;
        RECT 2276.270 4.000 2281.410 4.280 ;
        RECT 2282.250 4.000 2286.930 4.280 ;
        RECT 2287.770 4.000 2292.910 4.280 ;
        RECT 2293.750 4.000 2298.430 4.280 ;
        RECT 2299.270 4.000 2303.950 4.280 ;
        RECT 2304.790 4.000 2309.930 4.280 ;
        RECT 2310.770 4.000 2315.450 4.280 ;
        RECT 2316.290 4.000 2321.430 4.280 ;
        RECT 2322.270 4.000 2326.950 4.280 ;
        RECT 2327.790 4.000 2332.930 4.280 ;
        RECT 2333.770 4.000 2338.450 4.280 ;
        RECT 2339.290 4.000 2344.430 4.280 ;
        RECT 2345.270 4.000 2349.950 4.280 ;
        RECT 2350.790 4.000 2355.470 4.280 ;
        RECT 2356.310 4.000 2361.450 4.280 ;
        RECT 2362.290 4.000 2366.970 4.280 ;
        RECT 2367.810 4.000 2372.950 4.280 ;
        RECT 2373.790 4.000 2378.470 4.280 ;
        RECT 2379.310 4.000 2384.450 4.280 ;
        RECT 2385.290 4.000 2389.970 4.280 ;
        RECT 2390.810 4.000 2395.950 4.280 ;
        RECT 2396.790 4.000 2401.470 4.280 ;
        RECT 2402.310 4.000 2406.990 4.280 ;
        RECT 2407.830 4.000 2412.970 4.280 ;
        RECT 2413.810 4.000 2418.490 4.280 ;
        RECT 2419.330 4.000 2424.470 4.280 ;
        RECT 2425.310 4.000 2429.990 4.280 ;
        RECT 2430.830 4.000 2435.970 4.280 ;
        RECT 2436.810 4.000 2441.490 4.280 ;
        RECT 2442.330 4.000 2447.470 4.280 ;
        RECT 2448.310 4.000 2452.990 4.280 ;
        RECT 2453.830 4.000 2458.970 4.280 ;
        RECT 2459.810 4.000 2464.490 4.280 ;
        RECT 2465.330 4.000 2470.010 4.280 ;
        RECT 2470.850 4.000 2475.990 4.280 ;
        RECT 2476.830 4.000 2481.510 4.280 ;
        RECT 2482.350 4.000 2487.490 4.280 ;
        RECT 2488.330 4.000 2493.010 4.280 ;
        RECT 2493.850 4.000 2498.990 4.280 ;
        RECT 2499.830 4.000 2504.510 4.280 ;
        RECT 2505.350 4.000 2510.490 4.280 ;
        RECT 2511.330 4.000 2516.010 4.280 ;
        RECT 2516.850 4.000 2521.530 4.280 ;
        RECT 2522.370 4.000 2527.510 4.280 ;
        RECT 2528.350 4.000 2533.030 4.280 ;
        RECT 2533.870 4.000 2539.010 4.280 ;
        RECT 2539.850 4.000 2544.530 4.280 ;
        RECT 2545.370 4.000 2550.510 4.280 ;
        RECT 2551.350 4.000 2556.030 4.280 ;
        RECT 2556.870 4.000 2562.010 4.280 ;
        RECT 2562.850 4.000 2567.530 4.280 ;
        RECT 2568.370 4.000 2573.050 4.280 ;
        RECT 2573.890 4.000 2579.030 4.280 ;
        RECT 2579.870 4.000 2584.550 4.280 ;
        RECT 2585.390 4.000 2590.530 4.280 ;
        RECT 2591.370 4.000 2596.050 4.280 ;
        RECT 2596.890 4.000 2602.030 4.280 ;
        RECT 2602.870 4.000 2607.550 4.280 ;
        RECT 2608.390 4.000 2613.530 4.280 ;
        RECT 2614.370 4.000 2619.050 4.280 ;
        RECT 2619.890 4.000 2624.570 4.280 ;
        RECT 2625.410 4.000 2630.550 4.280 ;
        RECT 2631.390 4.000 2636.070 4.280 ;
        RECT 2636.910 4.000 2642.050 4.280 ;
        RECT 2642.890 4.000 2647.570 4.280 ;
        RECT 2648.410 4.000 2653.550 4.280 ;
        RECT 2654.390 4.000 2659.070 4.280 ;
        RECT 2659.910 4.000 2665.050 4.280 ;
        RECT 2665.890 4.000 2670.570 4.280 ;
        RECT 2671.410 4.000 2676.550 4.280 ;
        RECT 2677.390 4.000 2682.070 4.280 ;
        RECT 2682.910 4.000 2687.590 4.280 ;
        RECT 2688.430 4.000 2693.570 4.280 ;
        RECT 2694.410 4.000 2699.090 4.280 ;
        RECT 2699.930 4.000 2705.070 4.280 ;
        RECT 2705.910 4.000 2710.590 4.280 ;
        RECT 2711.430 4.000 2716.570 4.280 ;
        RECT 2717.410 4.000 2722.090 4.280 ;
        RECT 2722.930 4.000 2728.070 4.280 ;
        RECT 2728.910 4.000 2733.590 4.280 ;
        RECT 2734.430 4.000 2739.110 4.280 ;
        RECT 2739.950 4.000 2745.090 4.280 ;
        RECT 2745.930 4.000 2750.610 4.280 ;
        RECT 2751.450 4.000 2756.590 4.280 ;
        RECT 2757.430 4.000 2762.110 4.280 ;
        RECT 2762.950 4.000 2768.090 4.280 ;
        RECT 2768.930 4.000 2773.610 4.280 ;
        RECT 2774.450 4.000 2779.590 4.280 ;
        RECT 2780.430 4.000 2785.110 4.280 ;
        RECT 2785.950 4.000 2790.630 4.280 ;
        RECT 2791.470 4.000 2796.610 4.280 ;
        RECT 2797.450 4.000 2802.130 4.280 ;
        RECT 2802.970 4.000 2808.110 4.280 ;
      LAYER met3 ;
        RECT 12.025 10.715 2808.695 3427.365 ;
      LAYER met4 ;
        RECT 15.015 12.415 20.640 3418.185 ;
        RECT 23.040 12.415 97.440 3418.185 ;
        RECT 99.840 12.415 174.240 3418.185 ;
        RECT 176.640 12.415 251.040 3418.185 ;
        RECT 253.440 12.415 327.840 3418.185 ;
        RECT 330.240 12.415 404.640 3418.185 ;
        RECT 407.040 12.415 481.440 3418.185 ;
        RECT 483.840 12.415 558.240 3418.185 ;
        RECT 560.640 12.415 635.040 3418.185 ;
        RECT 637.440 12.415 711.840 3418.185 ;
        RECT 714.240 12.415 788.640 3418.185 ;
        RECT 791.040 12.415 865.440 3418.185 ;
        RECT 867.840 12.415 942.240 3418.185 ;
        RECT 944.640 12.415 1019.040 3418.185 ;
        RECT 1021.440 12.415 1095.840 3418.185 ;
        RECT 1098.240 12.415 1172.640 3418.185 ;
        RECT 1175.040 12.415 1249.440 3418.185 ;
        RECT 1251.840 12.415 1326.240 3418.185 ;
        RECT 1328.640 12.415 1403.040 3418.185 ;
        RECT 1405.440 12.415 1479.840 3418.185 ;
        RECT 1482.240 12.415 1556.640 3418.185 ;
        RECT 1559.040 12.415 1633.440 3418.185 ;
        RECT 1635.840 12.415 1710.240 3418.185 ;
        RECT 1712.640 12.415 1787.040 3418.185 ;
        RECT 1789.440 12.415 1863.840 3418.185 ;
        RECT 1866.240 12.415 1940.640 3418.185 ;
        RECT 1943.040 12.415 2017.440 3418.185 ;
        RECT 2019.840 12.415 2094.240 3418.185 ;
        RECT 2096.640 12.415 2171.040 3418.185 ;
        RECT 2173.440 12.415 2247.840 3418.185 ;
        RECT 2250.240 12.415 2324.640 3418.185 ;
        RECT 2327.040 12.415 2401.440 3418.185 ;
        RECT 2403.840 12.415 2478.240 3418.185 ;
        RECT 2480.640 12.415 2555.040 3418.185 ;
        RECT 2557.440 12.415 2631.840 3418.185 ;
        RECT 2634.240 12.415 2708.640 3418.185 ;
        RECT 2711.040 12.415 2748.665 3418.185 ;
  END
END user_proj_example
END LIBRARY


magic
tech sky130A
magscale 1 2
timestamp 1610237017
<< obsli1 >>
rect 1104 2159 566812 685457
<< obsm1 >>
rect 566 1232 566812 685488
<< metal2 >>
rect 2318 687200 2374 688000
rect 7010 687200 7066 688000
rect 11702 687200 11758 688000
rect 16486 687200 16542 688000
rect 21178 687200 21234 688000
rect 25962 687200 26018 688000
rect 30654 687200 30710 688000
rect 35438 687200 35494 688000
rect 40130 687200 40186 688000
rect 44914 687200 44970 688000
rect 49606 687200 49662 688000
rect 54298 687200 54354 688000
rect 59082 687200 59138 688000
rect 63774 687200 63830 688000
rect 68558 687200 68614 688000
rect 73250 687200 73306 688000
rect 78034 687200 78090 688000
rect 82726 687200 82782 688000
rect 87510 687200 87566 688000
rect 92202 687200 92258 688000
rect 96986 687200 97042 688000
rect 101678 687200 101734 688000
rect 106370 687200 106426 688000
rect 111154 687200 111210 688000
rect 115846 687200 115902 688000
rect 120630 687200 120686 688000
rect 125322 687200 125378 688000
rect 130106 687200 130162 688000
rect 134798 687200 134854 688000
rect 139582 687200 139638 688000
rect 144274 687200 144330 688000
rect 148966 687200 149022 688000
rect 153750 687200 153806 688000
rect 158442 687200 158498 688000
rect 163226 687200 163282 688000
rect 167918 687200 167974 688000
rect 172702 687200 172758 688000
rect 177394 687200 177450 688000
rect 182178 687200 182234 688000
rect 186870 687200 186926 688000
rect 191654 687200 191710 688000
rect 196346 687200 196402 688000
rect 201038 687200 201094 688000
rect 205822 687200 205878 688000
rect 210514 687200 210570 688000
rect 215298 687200 215354 688000
rect 219990 687200 220046 688000
rect 224774 687200 224830 688000
rect 229466 687200 229522 688000
rect 234250 687200 234306 688000
rect 238942 687200 238998 688000
rect 243634 687200 243690 688000
rect 248418 687200 248474 688000
rect 253110 687200 253166 688000
rect 257894 687200 257950 688000
rect 262586 687200 262642 688000
rect 267370 687200 267426 688000
rect 272062 687200 272118 688000
rect 276846 687200 276902 688000
rect 281538 687200 281594 688000
rect 286322 687200 286378 688000
rect 291014 687200 291070 688000
rect 295706 687200 295762 688000
rect 300490 687200 300546 688000
rect 305182 687200 305238 688000
rect 309966 687200 310022 688000
rect 314658 687200 314714 688000
rect 319442 687200 319498 688000
rect 324134 687200 324190 688000
rect 328918 687200 328974 688000
rect 333610 687200 333666 688000
rect 338302 687200 338358 688000
rect 343086 687200 343142 688000
rect 347778 687200 347834 688000
rect 352562 687200 352618 688000
rect 357254 687200 357310 688000
rect 362038 687200 362094 688000
rect 366730 687200 366786 688000
rect 371514 687200 371570 688000
rect 376206 687200 376262 688000
rect 380990 687200 381046 688000
rect 385682 687200 385738 688000
rect 390374 687200 390430 688000
rect 395158 687200 395214 688000
rect 399850 687200 399906 688000
rect 404634 687200 404690 688000
rect 409326 687200 409382 688000
rect 414110 687200 414166 688000
rect 418802 687200 418858 688000
rect 423586 687200 423642 688000
rect 428278 687200 428334 688000
rect 432970 687200 433026 688000
rect 437754 687200 437810 688000
rect 442446 687200 442502 688000
rect 447230 687200 447286 688000
rect 451922 687200 451978 688000
rect 456706 687200 456762 688000
rect 461398 687200 461454 688000
rect 466182 687200 466238 688000
rect 470874 687200 470930 688000
rect 475658 687200 475714 688000
rect 480350 687200 480406 688000
rect 485042 687200 485098 688000
rect 489826 687200 489882 688000
rect 494518 687200 494574 688000
rect 499302 687200 499358 688000
rect 503994 687200 504050 688000
rect 508778 687200 508834 688000
rect 513470 687200 513526 688000
rect 518254 687200 518310 688000
rect 522946 687200 523002 688000
rect 527638 687200 527694 688000
rect 532422 687200 532478 688000
rect 537114 687200 537170 688000
rect 541898 687200 541954 688000
rect 546590 687200 546646 688000
rect 551374 687200 551430 688000
rect 556066 687200 556122 688000
rect 560850 687200 560906 688000
rect 565542 687200 565598 688000
rect 570 0 626 800
rect 1674 0 1730 800
rect 2778 0 2834 800
rect 3882 0 3938 800
rect 5078 0 5134 800
rect 6182 0 6238 800
rect 7286 0 7342 800
rect 8482 0 8538 800
rect 9586 0 9642 800
rect 10690 0 10746 800
rect 11886 0 11942 800
rect 12990 0 13046 800
rect 14094 0 14150 800
rect 15290 0 15346 800
rect 16394 0 16450 800
rect 17498 0 17554 800
rect 18694 0 18750 800
rect 19798 0 19854 800
rect 20902 0 20958 800
rect 22098 0 22154 800
rect 23202 0 23258 800
rect 24306 0 24362 800
rect 25502 0 25558 800
rect 26606 0 26662 800
rect 27710 0 27766 800
rect 28906 0 28962 800
rect 30010 0 30066 800
rect 31114 0 31170 800
rect 32310 0 32366 800
rect 33414 0 33470 800
rect 34518 0 34574 800
rect 35714 0 35770 800
rect 36818 0 36874 800
rect 37922 0 37978 800
rect 39026 0 39082 800
rect 40222 0 40278 800
rect 41326 0 41382 800
rect 42430 0 42486 800
rect 43626 0 43682 800
rect 44730 0 44786 800
rect 45834 0 45890 800
rect 47030 0 47086 800
rect 48134 0 48190 800
rect 49238 0 49294 800
rect 50434 0 50490 800
rect 51538 0 51594 800
rect 52642 0 52698 800
rect 53838 0 53894 800
rect 54942 0 54998 800
rect 56046 0 56102 800
rect 57242 0 57298 800
rect 58346 0 58402 800
rect 59450 0 59506 800
rect 60646 0 60702 800
rect 61750 0 61806 800
rect 62854 0 62910 800
rect 64050 0 64106 800
rect 65154 0 65210 800
rect 66258 0 66314 800
rect 67454 0 67510 800
rect 68558 0 68614 800
rect 69662 0 69718 800
rect 70858 0 70914 800
rect 71962 0 72018 800
rect 73066 0 73122 800
rect 74262 0 74318 800
rect 75366 0 75422 800
rect 76470 0 76526 800
rect 77574 0 77630 800
rect 78770 0 78826 800
rect 79874 0 79930 800
rect 80978 0 81034 800
rect 82174 0 82230 800
rect 83278 0 83334 800
rect 84382 0 84438 800
rect 85578 0 85634 800
rect 86682 0 86738 800
rect 87786 0 87842 800
rect 88982 0 89038 800
rect 90086 0 90142 800
rect 91190 0 91246 800
rect 92386 0 92442 800
rect 93490 0 93546 800
rect 94594 0 94650 800
rect 95790 0 95846 800
rect 96894 0 96950 800
rect 97998 0 98054 800
rect 99194 0 99250 800
rect 100298 0 100354 800
rect 101402 0 101458 800
rect 102598 0 102654 800
rect 103702 0 103758 800
rect 104806 0 104862 800
rect 106002 0 106058 800
rect 107106 0 107162 800
rect 108210 0 108266 800
rect 109406 0 109462 800
rect 110510 0 110566 800
rect 111614 0 111670 800
rect 112810 0 112866 800
rect 113914 0 113970 800
rect 115018 0 115074 800
rect 116122 0 116178 800
rect 117318 0 117374 800
rect 118422 0 118478 800
rect 119526 0 119582 800
rect 120722 0 120778 800
rect 121826 0 121882 800
rect 122930 0 122986 800
rect 124126 0 124182 800
rect 125230 0 125286 800
rect 126334 0 126390 800
rect 127530 0 127586 800
rect 128634 0 128690 800
rect 129738 0 129794 800
rect 130934 0 130990 800
rect 132038 0 132094 800
rect 133142 0 133198 800
rect 134338 0 134394 800
rect 135442 0 135498 800
rect 136546 0 136602 800
rect 137742 0 137798 800
rect 138846 0 138902 800
rect 139950 0 140006 800
rect 141146 0 141202 800
rect 142250 0 142306 800
rect 143354 0 143410 800
rect 144550 0 144606 800
rect 145654 0 145710 800
rect 146758 0 146814 800
rect 147954 0 148010 800
rect 149058 0 149114 800
rect 150162 0 150218 800
rect 151358 0 151414 800
rect 152462 0 152518 800
rect 153566 0 153622 800
rect 154670 0 154726 800
rect 155866 0 155922 800
rect 156970 0 157026 800
rect 158074 0 158130 800
rect 159270 0 159326 800
rect 160374 0 160430 800
rect 161478 0 161534 800
rect 162674 0 162730 800
rect 163778 0 163834 800
rect 164882 0 164938 800
rect 166078 0 166134 800
rect 167182 0 167238 800
rect 168286 0 168342 800
rect 169482 0 169538 800
rect 170586 0 170642 800
rect 171690 0 171746 800
rect 172886 0 172942 800
rect 173990 0 174046 800
rect 175094 0 175150 800
rect 176290 0 176346 800
rect 177394 0 177450 800
rect 178498 0 178554 800
rect 179694 0 179750 800
rect 180798 0 180854 800
rect 181902 0 181958 800
rect 183098 0 183154 800
rect 184202 0 184258 800
rect 185306 0 185362 800
rect 186502 0 186558 800
rect 187606 0 187662 800
rect 188710 0 188766 800
rect 189906 0 189962 800
rect 191010 0 191066 800
rect 192114 0 192170 800
rect 193218 0 193274 800
rect 194414 0 194470 800
rect 195518 0 195574 800
rect 196622 0 196678 800
rect 197818 0 197874 800
rect 198922 0 198978 800
rect 200026 0 200082 800
rect 201222 0 201278 800
rect 202326 0 202382 800
rect 203430 0 203486 800
rect 204626 0 204682 800
rect 205730 0 205786 800
rect 206834 0 206890 800
rect 208030 0 208086 800
rect 209134 0 209190 800
rect 210238 0 210294 800
rect 211434 0 211490 800
rect 212538 0 212594 800
rect 213642 0 213698 800
rect 214838 0 214894 800
rect 215942 0 215998 800
rect 217046 0 217102 800
rect 218242 0 218298 800
rect 219346 0 219402 800
rect 220450 0 220506 800
rect 221646 0 221702 800
rect 222750 0 222806 800
rect 223854 0 223910 800
rect 225050 0 225106 800
rect 226154 0 226210 800
rect 227258 0 227314 800
rect 228362 0 228418 800
rect 229558 0 229614 800
rect 230662 0 230718 800
rect 231766 0 231822 800
rect 232962 0 233018 800
rect 234066 0 234122 800
rect 235170 0 235226 800
rect 236366 0 236422 800
rect 237470 0 237526 800
rect 238574 0 238630 800
rect 239770 0 239826 800
rect 240874 0 240930 800
rect 241978 0 242034 800
rect 243174 0 243230 800
rect 244278 0 244334 800
rect 245382 0 245438 800
rect 246578 0 246634 800
rect 247682 0 247738 800
rect 248786 0 248842 800
rect 249982 0 250038 800
rect 251086 0 251142 800
rect 252190 0 252246 800
rect 253386 0 253442 800
rect 254490 0 254546 800
rect 255594 0 255650 800
rect 256790 0 256846 800
rect 257894 0 257950 800
rect 258998 0 259054 800
rect 260194 0 260250 800
rect 261298 0 261354 800
rect 262402 0 262458 800
rect 263598 0 263654 800
rect 264702 0 264758 800
rect 265806 0 265862 800
rect 266910 0 266966 800
rect 268106 0 268162 800
rect 269210 0 269266 800
rect 270314 0 270370 800
rect 271510 0 271566 800
rect 272614 0 272670 800
rect 273718 0 273774 800
rect 274914 0 274970 800
rect 276018 0 276074 800
rect 277122 0 277178 800
rect 278318 0 278374 800
rect 279422 0 279478 800
rect 280526 0 280582 800
rect 281722 0 281778 800
rect 282826 0 282882 800
rect 283930 0 283986 800
rect 285126 0 285182 800
rect 286230 0 286286 800
rect 287334 0 287390 800
rect 288530 0 288586 800
rect 289634 0 289690 800
rect 290738 0 290794 800
rect 291934 0 291990 800
rect 293038 0 293094 800
rect 294142 0 294198 800
rect 295338 0 295394 800
rect 296442 0 296498 800
rect 297546 0 297602 800
rect 298742 0 298798 800
rect 299846 0 299902 800
rect 300950 0 301006 800
rect 302146 0 302202 800
rect 303250 0 303306 800
rect 304354 0 304410 800
rect 305458 0 305514 800
rect 306654 0 306710 800
rect 307758 0 307814 800
rect 308862 0 308918 800
rect 310058 0 310114 800
rect 311162 0 311218 800
rect 312266 0 312322 800
rect 313462 0 313518 800
rect 314566 0 314622 800
rect 315670 0 315726 800
rect 316866 0 316922 800
rect 317970 0 318026 800
rect 319074 0 319130 800
rect 320270 0 320326 800
rect 321374 0 321430 800
rect 322478 0 322534 800
rect 323674 0 323730 800
rect 324778 0 324834 800
rect 325882 0 325938 800
rect 327078 0 327134 800
rect 328182 0 328238 800
rect 329286 0 329342 800
rect 330482 0 330538 800
rect 331586 0 331642 800
rect 332690 0 332746 800
rect 333886 0 333942 800
rect 334990 0 335046 800
rect 336094 0 336150 800
rect 337290 0 337346 800
rect 338394 0 338450 800
rect 339498 0 339554 800
rect 340694 0 340750 800
rect 341798 0 341854 800
rect 342902 0 342958 800
rect 344006 0 344062 800
rect 345202 0 345258 800
rect 346306 0 346362 800
rect 347410 0 347466 800
rect 348606 0 348662 800
rect 349710 0 349766 800
rect 350814 0 350870 800
rect 352010 0 352066 800
rect 353114 0 353170 800
rect 354218 0 354274 800
rect 355414 0 355470 800
rect 356518 0 356574 800
rect 357622 0 357678 800
rect 358818 0 358874 800
rect 359922 0 359978 800
rect 361026 0 361082 800
rect 362222 0 362278 800
rect 363326 0 363382 800
rect 364430 0 364486 800
rect 365626 0 365682 800
rect 366730 0 366786 800
rect 367834 0 367890 800
rect 369030 0 369086 800
rect 370134 0 370190 800
rect 371238 0 371294 800
rect 372434 0 372490 800
rect 373538 0 373594 800
rect 374642 0 374698 800
rect 375838 0 375894 800
rect 376942 0 376998 800
rect 378046 0 378102 800
rect 379242 0 379298 800
rect 380346 0 380402 800
rect 381450 0 381506 800
rect 382554 0 382610 800
rect 383750 0 383806 800
rect 384854 0 384910 800
rect 385958 0 386014 800
rect 387154 0 387210 800
rect 388258 0 388314 800
rect 389362 0 389418 800
rect 390558 0 390614 800
rect 391662 0 391718 800
rect 392766 0 392822 800
rect 393962 0 394018 800
rect 395066 0 395122 800
rect 396170 0 396226 800
rect 397366 0 397422 800
rect 398470 0 398526 800
rect 399574 0 399630 800
rect 400770 0 400826 800
rect 401874 0 401930 800
rect 402978 0 403034 800
rect 404174 0 404230 800
rect 405278 0 405334 800
rect 406382 0 406438 800
rect 407578 0 407634 800
rect 408682 0 408738 800
rect 409786 0 409842 800
rect 410982 0 411038 800
rect 412086 0 412142 800
rect 413190 0 413246 800
rect 414386 0 414442 800
rect 415490 0 415546 800
rect 416594 0 416650 800
rect 417698 0 417754 800
rect 418894 0 418950 800
rect 419998 0 420054 800
rect 421102 0 421158 800
rect 422298 0 422354 800
rect 423402 0 423458 800
rect 424506 0 424562 800
rect 425702 0 425758 800
rect 426806 0 426862 800
rect 427910 0 427966 800
rect 429106 0 429162 800
rect 430210 0 430266 800
rect 431314 0 431370 800
rect 432510 0 432566 800
rect 433614 0 433670 800
rect 434718 0 434774 800
rect 435914 0 435970 800
rect 437018 0 437074 800
rect 438122 0 438178 800
rect 439318 0 439374 800
rect 440422 0 440478 800
rect 441526 0 441582 800
rect 442722 0 442778 800
rect 443826 0 443882 800
rect 444930 0 444986 800
rect 446126 0 446182 800
rect 447230 0 447286 800
rect 448334 0 448390 800
rect 449530 0 449586 800
rect 450634 0 450690 800
rect 451738 0 451794 800
rect 452934 0 452990 800
rect 454038 0 454094 800
rect 455142 0 455198 800
rect 456246 0 456302 800
rect 457442 0 457498 800
rect 458546 0 458602 800
rect 459650 0 459706 800
rect 460846 0 460902 800
rect 461950 0 462006 800
rect 463054 0 463110 800
rect 464250 0 464306 800
rect 465354 0 465410 800
rect 466458 0 466514 800
rect 467654 0 467710 800
rect 468758 0 468814 800
rect 469862 0 469918 800
rect 471058 0 471114 800
rect 472162 0 472218 800
rect 473266 0 473322 800
rect 474462 0 474518 800
rect 475566 0 475622 800
rect 476670 0 476726 800
rect 477866 0 477922 800
rect 478970 0 479026 800
rect 480074 0 480130 800
rect 481270 0 481326 800
rect 482374 0 482430 800
rect 483478 0 483534 800
rect 484674 0 484730 800
rect 485778 0 485834 800
rect 486882 0 486938 800
rect 488078 0 488134 800
rect 489182 0 489238 800
rect 490286 0 490342 800
rect 491482 0 491538 800
rect 492586 0 492642 800
rect 493690 0 493746 800
rect 494794 0 494850 800
rect 495990 0 496046 800
rect 497094 0 497150 800
rect 498198 0 498254 800
rect 499394 0 499450 800
rect 500498 0 500554 800
rect 501602 0 501658 800
rect 502798 0 502854 800
rect 503902 0 503958 800
rect 505006 0 505062 800
rect 506202 0 506258 800
rect 507306 0 507362 800
rect 508410 0 508466 800
rect 509606 0 509662 800
rect 510710 0 510766 800
rect 511814 0 511870 800
rect 513010 0 513066 800
rect 514114 0 514170 800
rect 515218 0 515274 800
rect 516414 0 516470 800
rect 517518 0 517574 800
rect 518622 0 518678 800
rect 519818 0 519874 800
rect 520922 0 520978 800
rect 522026 0 522082 800
rect 523222 0 523278 800
rect 524326 0 524382 800
rect 525430 0 525486 800
rect 526626 0 526682 800
rect 527730 0 527786 800
rect 528834 0 528890 800
rect 530030 0 530086 800
rect 531134 0 531190 800
rect 532238 0 532294 800
rect 533342 0 533398 800
rect 534538 0 534594 800
rect 535642 0 535698 800
rect 536746 0 536802 800
rect 537942 0 537998 800
rect 539046 0 539102 800
rect 540150 0 540206 800
rect 541346 0 541402 800
rect 542450 0 542506 800
rect 543554 0 543610 800
rect 544750 0 544806 800
rect 545854 0 545910 800
rect 546958 0 547014 800
rect 548154 0 548210 800
rect 549258 0 549314 800
rect 550362 0 550418 800
rect 551558 0 551614 800
rect 552662 0 552718 800
rect 553766 0 553822 800
rect 554962 0 555018 800
rect 556066 0 556122 800
rect 557170 0 557226 800
rect 558366 0 558422 800
rect 559470 0 559526 800
rect 560574 0 560630 800
rect 561770 0 561826 800
rect 562874 0 562930 800
rect 563978 0 564034 800
rect 565174 0 565230 800
rect 566278 0 566334 800
rect 567382 0 567438 800
<< obsm2 >>
rect 572 687144 2262 687200
rect 2430 687144 6954 687200
rect 7122 687144 11646 687200
rect 11814 687144 16430 687200
rect 16598 687144 21122 687200
rect 21290 687144 25906 687200
rect 26074 687144 30598 687200
rect 30766 687144 35382 687200
rect 35550 687144 40074 687200
rect 40242 687144 44858 687200
rect 45026 687144 49550 687200
rect 49718 687144 54242 687200
rect 54410 687144 59026 687200
rect 59194 687144 63718 687200
rect 63886 687144 68502 687200
rect 68670 687144 73194 687200
rect 73362 687144 77978 687200
rect 78146 687144 82670 687200
rect 82838 687144 87454 687200
rect 87622 687144 92146 687200
rect 92314 687144 96930 687200
rect 97098 687144 101622 687200
rect 101790 687144 106314 687200
rect 106482 687144 111098 687200
rect 111266 687144 115790 687200
rect 115958 687144 120574 687200
rect 120742 687144 125266 687200
rect 125434 687144 130050 687200
rect 130218 687144 134742 687200
rect 134910 687144 139526 687200
rect 139694 687144 144218 687200
rect 144386 687144 148910 687200
rect 149078 687144 153694 687200
rect 153862 687144 158386 687200
rect 158554 687144 163170 687200
rect 163338 687144 167862 687200
rect 168030 687144 172646 687200
rect 172814 687144 177338 687200
rect 177506 687144 182122 687200
rect 182290 687144 186814 687200
rect 186982 687144 191598 687200
rect 191766 687144 196290 687200
rect 196458 687144 200982 687200
rect 201150 687144 205766 687200
rect 205934 687144 210458 687200
rect 210626 687144 215242 687200
rect 215410 687144 219934 687200
rect 220102 687144 224718 687200
rect 224886 687144 229410 687200
rect 229578 687144 234194 687200
rect 234362 687144 238886 687200
rect 239054 687144 243578 687200
rect 243746 687144 248362 687200
rect 248530 687144 253054 687200
rect 253222 687144 257838 687200
rect 258006 687144 262530 687200
rect 262698 687144 267314 687200
rect 267482 687144 272006 687200
rect 272174 687144 276790 687200
rect 276958 687144 281482 687200
rect 281650 687144 286266 687200
rect 286434 687144 290958 687200
rect 291126 687144 295650 687200
rect 295818 687144 300434 687200
rect 300602 687144 305126 687200
rect 305294 687144 309910 687200
rect 310078 687144 314602 687200
rect 314770 687144 319386 687200
rect 319554 687144 324078 687200
rect 324246 687144 328862 687200
rect 329030 687144 333554 687200
rect 333722 687144 338246 687200
rect 338414 687144 343030 687200
rect 343198 687144 347722 687200
rect 347890 687144 352506 687200
rect 352674 687144 357198 687200
rect 357366 687144 361982 687200
rect 362150 687144 366674 687200
rect 366842 687144 371458 687200
rect 371626 687144 376150 687200
rect 376318 687144 380934 687200
rect 381102 687144 385626 687200
rect 385794 687144 390318 687200
rect 390486 687144 395102 687200
rect 395270 687144 399794 687200
rect 399962 687144 404578 687200
rect 404746 687144 409270 687200
rect 409438 687144 414054 687200
rect 414222 687144 418746 687200
rect 418914 687144 423530 687200
rect 423698 687144 428222 687200
rect 428390 687144 432914 687200
rect 433082 687144 437698 687200
rect 437866 687144 442390 687200
rect 442558 687144 447174 687200
rect 447342 687144 451866 687200
rect 452034 687144 456650 687200
rect 456818 687144 461342 687200
rect 461510 687144 466126 687200
rect 466294 687144 470818 687200
rect 470986 687144 475602 687200
rect 475770 687144 480294 687200
rect 480462 687144 484986 687200
rect 485154 687144 489770 687200
rect 489938 687144 494462 687200
rect 494630 687144 499246 687200
rect 499414 687144 503938 687200
rect 504106 687144 508722 687200
rect 508890 687144 513414 687200
rect 513582 687144 518198 687200
rect 518366 687144 522890 687200
rect 523058 687144 527582 687200
rect 527750 687144 532366 687200
rect 532534 687144 537058 687200
rect 537226 687144 541842 687200
rect 542010 687144 546534 687200
rect 546702 687144 551318 687200
rect 551486 687144 556010 687200
rect 556178 687144 557476 687200
rect 572 856 557476 687144
rect 682 800 1618 856
rect 1786 800 2722 856
rect 2890 800 3826 856
rect 3994 800 5022 856
rect 5190 800 6126 856
rect 6294 800 7230 856
rect 7398 800 8426 856
rect 8594 800 9530 856
rect 9698 800 10634 856
rect 10802 800 11830 856
rect 11998 800 12934 856
rect 13102 800 14038 856
rect 14206 800 15234 856
rect 15402 800 16338 856
rect 16506 800 17442 856
rect 17610 800 18638 856
rect 18806 800 19742 856
rect 19910 800 20846 856
rect 21014 800 22042 856
rect 22210 800 23146 856
rect 23314 800 24250 856
rect 24418 800 25446 856
rect 25614 800 26550 856
rect 26718 800 27654 856
rect 27822 800 28850 856
rect 29018 800 29954 856
rect 30122 800 31058 856
rect 31226 800 32254 856
rect 32422 800 33358 856
rect 33526 800 34462 856
rect 34630 800 35658 856
rect 35826 800 36762 856
rect 36930 800 37866 856
rect 38034 800 38970 856
rect 39138 800 40166 856
rect 40334 800 41270 856
rect 41438 800 42374 856
rect 42542 800 43570 856
rect 43738 800 44674 856
rect 44842 800 45778 856
rect 45946 800 46974 856
rect 47142 800 48078 856
rect 48246 800 49182 856
rect 49350 800 50378 856
rect 50546 800 51482 856
rect 51650 800 52586 856
rect 52754 800 53782 856
rect 53950 800 54886 856
rect 55054 800 55990 856
rect 56158 800 57186 856
rect 57354 800 58290 856
rect 58458 800 59394 856
rect 59562 800 60590 856
rect 60758 800 61694 856
rect 61862 800 62798 856
rect 62966 800 63994 856
rect 64162 800 65098 856
rect 65266 800 66202 856
rect 66370 800 67398 856
rect 67566 800 68502 856
rect 68670 800 69606 856
rect 69774 800 70802 856
rect 70970 800 71906 856
rect 72074 800 73010 856
rect 73178 800 74206 856
rect 74374 800 75310 856
rect 75478 800 76414 856
rect 76582 800 77518 856
rect 77686 800 78714 856
rect 78882 800 79818 856
rect 79986 800 80922 856
rect 81090 800 82118 856
rect 82286 800 83222 856
rect 83390 800 84326 856
rect 84494 800 85522 856
rect 85690 800 86626 856
rect 86794 800 87730 856
rect 87898 800 88926 856
rect 89094 800 90030 856
rect 90198 800 91134 856
rect 91302 800 92330 856
rect 92498 800 93434 856
rect 93602 800 94538 856
rect 94706 800 95734 856
rect 95902 800 96838 856
rect 97006 800 97942 856
rect 98110 800 99138 856
rect 99306 800 100242 856
rect 100410 800 101346 856
rect 101514 800 102542 856
rect 102710 800 103646 856
rect 103814 800 104750 856
rect 104918 800 105946 856
rect 106114 800 107050 856
rect 107218 800 108154 856
rect 108322 800 109350 856
rect 109518 800 110454 856
rect 110622 800 111558 856
rect 111726 800 112754 856
rect 112922 800 113858 856
rect 114026 800 114962 856
rect 115130 800 116066 856
rect 116234 800 117262 856
rect 117430 800 118366 856
rect 118534 800 119470 856
rect 119638 800 120666 856
rect 120834 800 121770 856
rect 121938 800 122874 856
rect 123042 800 124070 856
rect 124238 800 125174 856
rect 125342 800 126278 856
rect 126446 800 127474 856
rect 127642 800 128578 856
rect 128746 800 129682 856
rect 129850 800 130878 856
rect 131046 800 131982 856
rect 132150 800 133086 856
rect 133254 800 134282 856
rect 134450 800 135386 856
rect 135554 800 136490 856
rect 136658 800 137686 856
rect 137854 800 138790 856
rect 138958 800 139894 856
rect 140062 800 141090 856
rect 141258 800 142194 856
rect 142362 800 143298 856
rect 143466 800 144494 856
rect 144662 800 145598 856
rect 145766 800 146702 856
rect 146870 800 147898 856
rect 148066 800 149002 856
rect 149170 800 150106 856
rect 150274 800 151302 856
rect 151470 800 152406 856
rect 152574 800 153510 856
rect 153678 800 154614 856
rect 154782 800 155810 856
rect 155978 800 156914 856
rect 157082 800 158018 856
rect 158186 800 159214 856
rect 159382 800 160318 856
rect 160486 800 161422 856
rect 161590 800 162618 856
rect 162786 800 163722 856
rect 163890 800 164826 856
rect 164994 800 166022 856
rect 166190 800 167126 856
rect 167294 800 168230 856
rect 168398 800 169426 856
rect 169594 800 170530 856
rect 170698 800 171634 856
rect 171802 800 172830 856
rect 172998 800 173934 856
rect 174102 800 175038 856
rect 175206 800 176234 856
rect 176402 800 177338 856
rect 177506 800 178442 856
rect 178610 800 179638 856
rect 179806 800 180742 856
rect 180910 800 181846 856
rect 182014 800 183042 856
rect 183210 800 184146 856
rect 184314 800 185250 856
rect 185418 800 186446 856
rect 186614 800 187550 856
rect 187718 800 188654 856
rect 188822 800 189850 856
rect 190018 800 190954 856
rect 191122 800 192058 856
rect 192226 800 193162 856
rect 193330 800 194358 856
rect 194526 800 195462 856
rect 195630 800 196566 856
rect 196734 800 197762 856
rect 197930 800 198866 856
rect 199034 800 199970 856
rect 200138 800 201166 856
rect 201334 800 202270 856
rect 202438 800 203374 856
rect 203542 800 204570 856
rect 204738 800 205674 856
rect 205842 800 206778 856
rect 206946 800 207974 856
rect 208142 800 209078 856
rect 209246 800 210182 856
rect 210350 800 211378 856
rect 211546 800 212482 856
rect 212650 800 213586 856
rect 213754 800 214782 856
rect 214950 800 215886 856
rect 216054 800 216990 856
rect 217158 800 218186 856
rect 218354 800 219290 856
rect 219458 800 220394 856
rect 220562 800 221590 856
rect 221758 800 222694 856
rect 222862 800 223798 856
rect 223966 800 224994 856
rect 225162 800 226098 856
rect 226266 800 227202 856
rect 227370 800 228306 856
rect 228474 800 229502 856
rect 229670 800 230606 856
rect 230774 800 231710 856
rect 231878 800 232906 856
rect 233074 800 234010 856
rect 234178 800 235114 856
rect 235282 800 236310 856
rect 236478 800 237414 856
rect 237582 800 238518 856
rect 238686 800 239714 856
rect 239882 800 240818 856
rect 240986 800 241922 856
rect 242090 800 243118 856
rect 243286 800 244222 856
rect 244390 800 245326 856
rect 245494 800 246522 856
rect 246690 800 247626 856
rect 247794 800 248730 856
rect 248898 800 249926 856
rect 250094 800 251030 856
rect 251198 800 252134 856
rect 252302 800 253330 856
rect 253498 800 254434 856
rect 254602 800 255538 856
rect 255706 800 256734 856
rect 256902 800 257838 856
rect 258006 800 258942 856
rect 259110 800 260138 856
rect 260306 800 261242 856
rect 261410 800 262346 856
rect 262514 800 263542 856
rect 263710 800 264646 856
rect 264814 800 265750 856
rect 265918 800 266854 856
rect 267022 800 268050 856
rect 268218 800 269154 856
rect 269322 800 270258 856
rect 270426 800 271454 856
rect 271622 800 272558 856
rect 272726 800 273662 856
rect 273830 800 274858 856
rect 275026 800 275962 856
rect 276130 800 277066 856
rect 277234 800 278262 856
rect 278430 800 279366 856
rect 279534 800 280470 856
rect 280638 800 281666 856
rect 281834 800 282770 856
rect 282938 800 283874 856
rect 284042 800 285070 856
rect 285238 800 286174 856
rect 286342 800 287278 856
rect 287446 800 288474 856
rect 288642 800 289578 856
rect 289746 800 290682 856
rect 290850 800 291878 856
rect 292046 800 292982 856
rect 293150 800 294086 856
rect 294254 800 295282 856
rect 295450 800 296386 856
rect 296554 800 297490 856
rect 297658 800 298686 856
rect 298854 800 299790 856
rect 299958 800 300894 856
rect 301062 800 302090 856
rect 302258 800 303194 856
rect 303362 800 304298 856
rect 304466 800 305402 856
rect 305570 800 306598 856
rect 306766 800 307702 856
rect 307870 800 308806 856
rect 308974 800 310002 856
rect 310170 800 311106 856
rect 311274 800 312210 856
rect 312378 800 313406 856
rect 313574 800 314510 856
rect 314678 800 315614 856
rect 315782 800 316810 856
rect 316978 800 317914 856
rect 318082 800 319018 856
rect 319186 800 320214 856
rect 320382 800 321318 856
rect 321486 800 322422 856
rect 322590 800 323618 856
rect 323786 800 324722 856
rect 324890 800 325826 856
rect 325994 800 327022 856
rect 327190 800 328126 856
rect 328294 800 329230 856
rect 329398 800 330426 856
rect 330594 800 331530 856
rect 331698 800 332634 856
rect 332802 800 333830 856
rect 333998 800 334934 856
rect 335102 800 336038 856
rect 336206 800 337234 856
rect 337402 800 338338 856
rect 338506 800 339442 856
rect 339610 800 340638 856
rect 340806 800 341742 856
rect 341910 800 342846 856
rect 343014 800 343950 856
rect 344118 800 345146 856
rect 345314 800 346250 856
rect 346418 800 347354 856
rect 347522 800 348550 856
rect 348718 800 349654 856
rect 349822 800 350758 856
rect 350926 800 351954 856
rect 352122 800 353058 856
rect 353226 800 354162 856
rect 354330 800 355358 856
rect 355526 800 356462 856
rect 356630 800 357566 856
rect 357734 800 358762 856
rect 358930 800 359866 856
rect 360034 800 360970 856
rect 361138 800 362166 856
rect 362334 800 363270 856
rect 363438 800 364374 856
rect 364542 800 365570 856
rect 365738 800 366674 856
rect 366842 800 367778 856
rect 367946 800 368974 856
rect 369142 800 370078 856
rect 370246 800 371182 856
rect 371350 800 372378 856
rect 372546 800 373482 856
rect 373650 800 374586 856
rect 374754 800 375782 856
rect 375950 800 376886 856
rect 377054 800 377990 856
rect 378158 800 379186 856
rect 379354 800 380290 856
rect 380458 800 381394 856
rect 381562 800 382498 856
rect 382666 800 383694 856
rect 383862 800 384798 856
rect 384966 800 385902 856
rect 386070 800 387098 856
rect 387266 800 388202 856
rect 388370 800 389306 856
rect 389474 800 390502 856
rect 390670 800 391606 856
rect 391774 800 392710 856
rect 392878 800 393906 856
rect 394074 800 395010 856
rect 395178 800 396114 856
rect 396282 800 397310 856
rect 397478 800 398414 856
rect 398582 800 399518 856
rect 399686 800 400714 856
rect 400882 800 401818 856
rect 401986 800 402922 856
rect 403090 800 404118 856
rect 404286 800 405222 856
rect 405390 800 406326 856
rect 406494 800 407522 856
rect 407690 800 408626 856
rect 408794 800 409730 856
rect 409898 800 410926 856
rect 411094 800 412030 856
rect 412198 800 413134 856
rect 413302 800 414330 856
rect 414498 800 415434 856
rect 415602 800 416538 856
rect 416706 800 417642 856
rect 417810 800 418838 856
rect 419006 800 419942 856
rect 420110 800 421046 856
rect 421214 800 422242 856
rect 422410 800 423346 856
rect 423514 800 424450 856
rect 424618 800 425646 856
rect 425814 800 426750 856
rect 426918 800 427854 856
rect 428022 800 429050 856
rect 429218 800 430154 856
rect 430322 800 431258 856
rect 431426 800 432454 856
rect 432622 800 433558 856
rect 433726 800 434662 856
rect 434830 800 435858 856
rect 436026 800 436962 856
rect 437130 800 438066 856
rect 438234 800 439262 856
rect 439430 800 440366 856
rect 440534 800 441470 856
rect 441638 800 442666 856
rect 442834 800 443770 856
rect 443938 800 444874 856
rect 445042 800 446070 856
rect 446238 800 447174 856
rect 447342 800 448278 856
rect 448446 800 449474 856
rect 449642 800 450578 856
rect 450746 800 451682 856
rect 451850 800 452878 856
rect 453046 800 453982 856
rect 454150 800 455086 856
rect 455254 800 456190 856
rect 456358 800 457386 856
rect 457554 800 458490 856
rect 458658 800 459594 856
rect 459762 800 460790 856
rect 460958 800 461894 856
rect 462062 800 462998 856
rect 463166 800 464194 856
rect 464362 800 465298 856
rect 465466 800 466402 856
rect 466570 800 467598 856
rect 467766 800 468702 856
rect 468870 800 469806 856
rect 469974 800 471002 856
rect 471170 800 472106 856
rect 472274 800 473210 856
rect 473378 800 474406 856
rect 474574 800 475510 856
rect 475678 800 476614 856
rect 476782 800 477810 856
rect 477978 800 478914 856
rect 479082 800 480018 856
rect 480186 800 481214 856
rect 481382 800 482318 856
rect 482486 800 483422 856
rect 483590 800 484618 856
rect 484786 800 485722 856
rect 485890 800 486826 856
rect 486994 800 488022 856
rect 488190 800 489126 856
rect 489294 800 490230 856
rect 490398 800 491426 856
rect 491594 800 492530 856
rect 492698 800 493634 856
rect 493802 800 494738 856
rect 494906 800 495934 856
rect 496102 800 497038 856
rect 497206 800 498142 856
rect 498310 800 499338 856
rect 499506 800 500442 856
rect 500610 800 501546 856
rect 501714 800 502742 856
rect 502910 800 503846 856
rect 504014 800 504950 856
rect 505118 800 506146 856
rect 506314 800 507250 856
rect 507418 800 508354 856
rect 508522 800 509550 856
rect 509718 800 510654 856
rect 510822 800 511758 856
rect 511926 800 512954 856
rect 513122 800 514058 856
rect 514226 800 515162 856
rect 515330 800 516358 856
rect 516526 800 517462 856
rect 517630 800 518566 856
rect 518734 800 519762 856
rect 519930 800 520866 856
rect 521034 800 521970 856
rect 522138 800 523166 856
rect 523334 800 524270 856
rect 524438 800 525374 856
rect 525542 800 526570 856
rect 526738 800 527674 856
rect 527842 800 528778 856
rect 528946 800 529974 856
rect 530142 800 531078 856
rect 531246 800 532182 856
rect 532350 800 533286 856
rect 533454 800 534482 856
rect 534650 800 535586 856
rect 535754 800 536690 856
rect 536858 800 537886 856
rect 538054 800 538990 856
rect 539158 800 540094 856
rect 540262 800 541290 856
rect 541458 800 542394 856
rect 542562 800 543498 856
rect 543666 800 544694 856
rect 544862 800 545798 856
rect 545966 800 546902 856
rect 547070 800 548098 856
rect 548266 800 549202 856
rect 549370 800 550306 856
rect 550474 800 551502 856
rect 551670 800 552606 856
rect 552774 800 553710 856
rect 553878 800 554906 856
rect 555074 800 556010 856
rect 556178 800 557114 856
rect 557282 800 557476 856
<< metal3 >>
rect 0 653488 800 653608
rect 0 584672 800 584792
rect 0 515856 800 515976
rect 0 447040 800 447160
rect 0 378224 800 378344
rect 0 309408 800 309528
rect 0 240592 800 240712
rect 0 171776 800 171896
rect 0 102960 800 103080
rect 0 34280 800 34400
rect 567200 619080 568000 619200
rect 567200 481448 568000 481568
rect 567200 343816 568000 343936
rect 567200 206184 568000 206304
rect 567200 68688 568000 68808
<< obsm3 >>
rect 2497 2143 557488 685473
<< metal4 >>
rect 4208 2128 4528 685488
rect 19568 2128 19888 685488
rect 34928 2128 35248 685488
rect 50288 2128 50608 685488
rect 65648 2128 65968 685488
rect 81008 2128 81328 685488
rect 96368 2128 96688 685488
rect 111728 2128 112048 685488
rect 127088 2128 127408 685488
rect 142448 2128 142768 685488
rect 157808 2128 158128 685488
rect 173168 2128 173488 685488
rect 188528 2128 188848 685488
rect 203888 2128 204208 685488
rect 219248 2128 219568 685488
rect 234608 2128 234928 685488
rect 249968 2128 250288 685488
rect 265328 2128 265648 685488
rect 280688 2128 281008 685488
rect 296048 2128 296368 685488
rect 311408 2128 311728 685488
rect 326768 2128 327088 685488
rect 342128 2128 342448 685488
rect 357488 2128 357808 685488
rect 372848 2128 373168 685488
rect 388208 2128 388528 685488
rect 403568 2128 403888 685488
rect 418928 2128 419248 685488
rect 434288 2128 434608 685488
rect 449648 2128 449968 685488
rect 465008 2128 465328 685488
rect 480368 2128 480688 685488
rect 495728 2128 496048 685488
rect 511088 2128 511408 685488
rect 526448 2128 526768 685488
rect 541808 2128 542128 685488
rect 557168 2128 557488 685488
<< obsm4 >>
rect 3003 2211 4128 683229
rect 4608 2211 19488 683229
rect 19968 2211 34848 683229
rect 35328 2211 50208 683229
rect 50688 2211 65568 683229
rect 66048 2211 80928 683229
rect 81408 2211 96288 683229
rect 96768 2211 111648 683229
rect 112128 2211 127008 683229
rect 127488 2211 142368 683229
rect 142848 2211 157728 683229
rect 158208 2211 173088 683229
rect 173568 2211 188448 683229
rect 188928 2211 203808 683229
rect 204288 2211 219168 683229
rect 219648 2211 234528 683229
rect 235008 2211 249888 683229
rect 250368 2211 265248 683229
rect 265728 2211 280608 683229
rect 281088 2211 295968 683229
rect 296448 2211 311328 683229
rect 311808 2211 326688 683229
rect 327168 2211 342048 683229
rect 342528 2211 357408 683229
rect 357888 2211 372768 683229
rect 373248 2211 388128 683229
rect 388608 2211 403488 683229
rect 403968 2211 418848 683229
rect 419328 2211 434208 683229
rect 434688 2211 449568 683229
rect 450048 2211 464928 683229
rect 465408 2211 480288 683229
rect 480768 2211 495648 683229
rect 496128 2211 511008 683229
rect 511488 2211 526368 683229
rect 526848 2211 541728 683229
rect 542208 2211 549181 683229
<< labels >>
rlabel metal3 s 0 34280 800 34400 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal3 s 0 309408 800 309528 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 560574 0 560630 800 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 546590 687200 546646 688000 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal3 s 0 378224 800 378344 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal3 s 0 447040 800 447160 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 551374 687200 551430 688000 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal3 s 567200 343816 568000 343936 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal2 s 556066 687200 556122 688000 6 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal2 s 561770 0 561826 800 6 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal2 s 560850 687200 560906 688000 6 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal2 s 557170 0 557226 800 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s 567200 481448 568000 481568 6 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal2 s 565542 687200 565598 688000 6 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s 0 515856 800 515976 6 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal2 s 562874 0 562930 800 6 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s 567200 619080 568000 619200 6 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s 0 584672 800 584792 6 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal2 s 563978 0 564034 800 6 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal2 s 565174 0 565230 800 6 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal2 s 566278 0 566334 800 6 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 0 653488 800 653608 6 analog_io[29]
port 22 nsew signal bidirectional
rlabel metal3 s 567200 68688 568000 68808 6 analog_io[2]
port 23 nsew signal bidirectional
rlabel metal2 s 567382 0 567438 800 6 analog_io[30]
port 24 nsew signal bidirectional
rlabel metal2 s 558366 0 558422 800 6 analog_io[3]
port 25 nsew signal bidirectional
rlabel metal3 s 0 102960 800 103080 6 analog_io[4]
port 26 nsew signal bidirectional
rlabel metal3 s 0 171776 800 171896 6 analog_io[5]
port 27 nsew signal bidirectional
rlabel metal3 s 0 240592 800 240712 6 analog_io[6]
port 28 nsew signal bidirectional
rlabel metal3 s 567200 206184 568000 206304 6 analog_io[7]
port 29 nsew signal bidirectional
rlabel metal2 s 559470 0 559526 800 6 analog_io[8]
port 30 nsew signal bidirectional
rlabel metal2 s 541898 687200 541954 688000 6 analog_io[9]
port 31 nsew signal bidirectional
rlabel metal2 s 2318 687200 2374 688000 6 io_in[0]
port 32 nsew signal input
rlabel metal2 s 144274 687200 144330 688000 6 io_in[10]
port 33 nsew signal input
rlabel metal2 s 158442 687200 158498 688000 6 io_in[11]
port 34 nsew signal input
rlabel metal2 s 172702 687200 172758 688000 6 io_in[12]
port 35 nsew signal input
rlabel metal2 s 186870 687200 186926 688000 6 io_in[13]
port 36 nsew signal input
rlabel metal2 s 201038 687200 201094 688000 6 io_in[14]
port 37 nsew signal input
rlabel metal2 s 215298 687200 215354 688000 6 io_in[15]
port 38 nsew signal input
rlabel metal2 s 229466 687200 229522 688000 6 io_in[16]
port 39 nsew signal input
rlabel metal2 s 243634 687200 243690 688000 6 io_in[17]
port 40 nsew signal input
rlabel metal2 s 257894 687200 257950 688000 6 io_in[18]
port 41 nsew signal input
rlabel metal2 s 272062 687200 272118 688000 6 io_in[19]
port 42 nsew signal input
rlabel metal2 s 16486 687200 16542 688000 6 io_in[1]
port 43 nsew signal input
rlabel metal2 s 286322 687200 286378 688000 6 io_in[20]
port 44 nsew signal input
rlabel metal2 s 300490 687200 300546 688000 6 io_in[21]
port 45 nsew signal input
rlabel metal2 s 314658 687200 314714 688000 6 io_in[22]
port 46 nsew signal input
rlabel metal2 s 328918 687200 328974 688000 6 io_in[23]
port 47 nsew signal input
rlabel metal2 s 343086 687200 343142 688000 6 io_in[24]
port 48 nsew signal input
rlabel metal2 s 357254 687200 357310 688000 6 io_in[25]
port 49 nsew signal input
rlabel metal2 s 371514 687200 371570 688000 6 io_in[26]
port 50 nsew signal input
rlabel metal2 s 385682 687200 385738 688000 6 io_in[27]
port 51 nsew signal input
rlabel metal2 s 399850 687200 399906 688000 6 io_in[28]
port 52 nsew signal input
rlabel metal2 s 414110 687200 414166 688000 6 io_in[29]
port 53 nsew signal input
rlabel metal2 s 30654 687200 30710 688000 6 io_in[2]
port 54 nsew signal input
rlabel metal2 s 428278 687200 428334 688000 6 io_in[30]
port 55 nsew signal input
rlabel metal2 s 442446 687200 442502 688000 6 io_in[31]
port 56 nsew signal input
rlabel metal2 s 456706 687200 456762 688000 6 io_in[32]
port 57 nsew signal input
rlabel metal2 s 470874 687200 470930 688000 6 io_in[33]
port 58 nsew signal input
rlabel metal2 s 485042 687200 485098 688000 6 io_in[34]
port 59 nsew signal input
rlabel metal2 s 499302 687200 499358 688000 6 io_in[35]
port 60 nsew signal input
rlabel metal2 s 513470 687200 513526 688000 6 io_in[36]
port 61 nsew signal input
rlabel metal2 s 527638 687200 527694 688000 6 io_in[37]
port 62 nsew signal input
rlabel metal2 s 44914 687200 44970 688000 6 io_in[3]
port 63 nsew signal input
rlabel metal2 s 59082 687200 59138 688000 6 io_in[4]
port 64 nsew signal input
rlabel metal2 s 73250 687200 73306 688000 6 io_in[5]
port 65 nsew signal input
rlabel metal2 s 87510 687200 87566 688000 6 io_in[6]
port 66 nsew signal input
rlabel metal2 s 101678 687200 101734 688000 6 io_in[7]
port 67 nsew signal input
rlabel metal2 s 115846 687200 115902 688000 6 io_in[8]
port 68 nsew signal input
rlabel metal2 s 130106 687200 130162 688000 6 io_in[9]
port 69 nsew signal input
rlabel metal2 s 7010 687200 7066 688000 6 io_oeb[0]
port 70 nsew signal output
rlabel metal2 s 148966 687200 149022 688000 6 io_oeb[10]
port 71 nsew signal output
rlabel metal2 s 163226 687200 163282 688000 6 io_oeb[11]
port 72 nsew signal output
rlabel metal2 s 177394 687200 177450 688000 6 io_oeb[12]
port 73 nsew signal output
rlabel metal2 s 191654 687200 191710 688000 6 io_oeb[13]
port 74 nsew signal output
rlabel metal2 s 205822 687200 205878 688000 6 io_oeb[14]
port 75 nsew signal output
rlabel metal2 s 219990 687200 220046 688000 6 io_oeb[15]
port 76 nsew signal output
rlabel metal2 s 234250 687200 234306 688000 6 io_oeb[16]
port 77 nsew signal output
rlabel metal2 s 248418 687200 248474 688000 6 io_oeb[17]
port 78 nsew signal output
rlabel metal2 s 262586 687200 262642 688000 6 io_oeb[18]
port 79 nsew signal output
rlabel metal2 s 276846 687200 276902 688000 6 io_oeb[19]
port 80 nsew signal output
rlabel metal2 s 21178 687200 21234 688000 6 io_oeb[1]
port 81 nsew signal output
rlabel metal2 s 291014 687200 291070 688000 6 io_oeb[20]
port 82 nsew signal output
rlabel metal2 s 305182 687200 305238 688000 6 io_oeb[21]
port 83 nsew signal output
rlabel metal2 s 319442 687200 319498 688000 6 io_oeb[22]
port 84 nsew signal output
rlabel metal2 s 333610 687200 333666 688000 6 io_oeb[23]
port 85 nsew signal output
rlabel metal2 s 347778 687200 347834 688000 6 io_oeb[24]
port 86 nsew signal output
rlabel metal2 s 362038 687200 362094 688000 6 io_oeb[25]
port 87 nsew signal output
rlabel metal2 s 376206 687200 376262 688000 6 io_oeb[26]
port 88 nsew signal output
rlabel metal2 s 390374 687200 390430 688000 6 io_oeb[27]
port 89 nsew signal output
rlabel metal2 s 404634 687200 404690 688000 6 io_oeb[28]
port 90 nsew signal output
rlabel metal2 s 418802 687200 418858 688000 6 io_oeb[29]
port 91 nsew signal output
rlabel metal2 s 35438 687200 35494 688000 6 io_oeb[2]
port 92 nsew signal output
rlabel metal2 s 432970 687200 433026 688000 6 io_oeb[30]
port 93 nsew signal output
rlabel metal2 s 447230 687200 447286 688000 6 io_oeb[31]
port 94 nsew signal output
rlabel metal2 s 461398 687200 461454 688000 6 io_oeb[32]
port 95 nsew signal output
rlabel metal2 s 475658 687200 475714 688000 6 io_oeb[33]
port 96 nsew signal output
rlabel metal2 s 489826 687200 489882 688000 6 io_oeb[34]
port 97 nsew signal output
rlabel metal2 s 503994 687200 504050 688000 6 io_oeb[35]
port 98 nsew signal output
rlabel metal2 s 518254 687200 518310 688000 6 io_oeb[36]
port 99 nsew signal output
rlabel metal2 s 532422 687200 532478 688000 6 io_oeb[37]
port 100 nsew signal output
rlabel metal2 s 49606 687200 49662 688000 6 io_oeb[3]
port 101 nsew signal output
rlabel metal2 s 63774 687200 63830 688000 6 io_oeb[4]
port 102 nsew signal output
rlabel metal2 s 78034 687200 78090 688000 6 io_oeb[5]
port 103 nsew signal output
rlabel metal2 s 92202 687200 92258 688000 6 io_oeb[6]
port 104 nsew signal output
rlabel metal2 s 106370 687200 106426 688000 6 io_oeb[7]
port 105 nsew signal output
rlabel metal2 s 120630 687200 120686 688000 6 io_oeb[8]
port 106 nsew signal output
rlabel metal2 s 134798 687200 134854 688000 6 io_oeb[9]
port 107 nsew signal output
rlabel metal2 s 11702 687200 11758 688000 6 io_out[0]
port 108 nsew signal output
rlabel metal2 s 153750 687200 153806 688000 6 io_out[10]
port 109 nsew signal output
rlabel metal2 s 167918 687200 167974 688000 6 io_out[11]
port 110 nsew signal output
rlabel metal2 s 182178 687200 182234 688000 6 io_out[12]
port 111 nsew signal output
rlabel metal2 s 196346 687200 196402 688000 6 io_out[13]
port 112 nsew signal output
rlabel metal2 s 210514 687200 210570 688000 6 io_out[14]
port 113 nsew signal output
rlabel metal2 s 224774 687200 224830 688000 6 io_out[15]
port 114 nsew signal output
rlabel metal2 s 238942 687200 238998 688000 6 io_out[16]
port 115 nsew signal output
rlabel metal2 s 253110 687200 253166 688000 6 io_out[17]
port 116 nsew signal output
rlabel metal2 s 267370 687200 267426 688000 6 io_out[18]
port 117 nsew signal output
rlabel metal2 s 281538 687200 281594 688000 6 io_out[19]
port 118 nsew signal output
rlabel metal2 s 25962 687200 26018 688000 6 io_out[1]
port 119 nsew signal output
rlabel metal2 s 295706 687200 295762 688000 6 io_out[20]
port 120 nsew signal output
rlabel metal2 s 309966 687200 310022 688000 6 io_out[21]
port 121 nsew signal output
rlabel metal2 s 324134 687200 324190 688000 6 io_out[22]
port 122 nsew signal output
rlabel metal2 s 338302 687200 338358 688000 6 io_out[23]
port 123 nsew signal output
rlabel metal2 s 352562 687200 352618 688000 6 io_out[24]
port 124 nsew signal output
rlabel metal2 s 366730 687200 366786 688000 6 io_out[25]
port 125 nsew signal output
rlabel metal2 s 380990 687200 381046 688000 6 io_out[26]
port 126 nsew signal output
rlabel metal2 s 395158 687200 395214 688000 6 io_out[27]
port 127 nsew signal output
rlabel metal2 s 409326 687200 409382 688000 6 io_out[28]
port 128 nsew signal output
rlabel metal2 s 423586 687200 423642 688000 6 io_out[29]
port 129 nsew signal output
rlabel metal2 s 40130 687200 40186 688000 6 io_out[2]
port 130 nsew signal output
rlabel metal2 s 437754 687200 437810 688000 6 io_out[30]
port 131 nsew signal output
rlabel metal2 s 451922 687200 451978 688000 6 io_out[31]
port 132 nsew signal output
rlabel metal2 s 466182 687200 466238 688000 6 io_out[32]
port 133 nsew signal output
rlabel metal2 s 480350 687200 480406 688000 6 io_out[33]
port 134 nsew signal output
rlabel metal2 s 494518 687200 494574 688000 6 io_out[34]
port 135 nsew signal output
rlabel metal2 s 508778 687200 508834 688000 6 io_out[35]
port 136 nsew signal output
rlabel metal2 s 522946 687200 523002 688000 6 io_out[36]
port 137 nsew signal output
rlabel metal2 s 537114 687200 537170 688000 6 io_out[37]
port 138 nsew signal output
rlabel metal2 s 54298 687200 54354 688000 6 io_out[3]
port 139 nsew signal output
rlabel metal2 s 68558 687200 68614 688000 6 io_out[4]
port 140 nsew signal output
rlabel metal2 s 82726 687200 82782 688000 6 io_out[5]
port 141 nsew signal output
rlabel metal2 s 96986 687200 97042 688000 6 io_out[6]
port 142 nsew signal output
rlabel metal2 s 111154 687200 111210 688000 6 io_out[7]
port 143 nsew signal output
rlabel metal2 s 125322 687200 125378 688000 6 io_out[8]
port 144 nsew signal output
rlabel metal2 s 139582 687200 139638 688000 6 io_out[9]
port 145 nsew signal output
rlabel metal2 s 120722 0 120778 800 6 la_data_in[0]
port 146 nsew signal input
rlabel metal2 s 460846 0 460902 800 6 la_data_in[100]
port 147 nsew signal input
rlabel metal2 s 464250 0 464306 800 6 la_data_in[101]
port 148 nsew signal input
rlabel metal2 s 467654 0 467710 800 6 la_data_in[102]
port 149 nsew signal input
rlabel metal2 s 471058 0 471114 800 6 la_data_in[103]
port 150 nsew signal input
rlabel metal2 s 474462 0 474518 800 6 la_data_in[104]
port 151 nsew signal input
rlabel metal2 s 477866 0 477922 800 6 la_data_in[105]
port 152 nsew signal input
rlabel metal2 s 481270 0 481326 800 6 la_data_in[106]
port 153 nsew signal input
rlabel metal2 s 484674 0 484730 800 6 la_data_in[107]
port 154 nsew signal input
rlabel metal2 s 488078 0 488134 800 6 la_data_in[108]
port 155 nsew signal input
rlabel metal2 s 491482 0 491538 800 6 la_data_in[109]
port 156 nsew signal input
rlabel metal2 s 154670 0 154726 800 6 la_data_in[10]
port 157 nsew signal input
rlabel metal2 s 494794 0 494850 800 6 la_data_in[110]
port 158 nsew signal input
rlabel metal2 s 498198 0 498254 800 6 la_data_in[111]
port 159 nsew signal input
rlabel metal2 s 501602 0 501658 800 6 la_data_in[112]
port 160 nsew signal input
rlabel metal2 s 505006 0 505062 800 6 la_data_in[113]
port 161 nsew signal input
rlabel metal2 s 508410 0 508466 800 6 la_data_in[114]
port 162 nsew signal input
rlabel metal2 s 511814 0 511870 800 6 la_data_in[115]
port 163 nsew signal input
rlabel metal2 s 515218 0 515274 800 6 la_data_in[116]
port 164 nsew signal input
rlabel metal2 s 518622 0 518678 800 6 la_data_in[117]
port 165 nsew signal input
rlabel metal2 s 522026 0 522082 800 6 la_data_in[118]
port 166 nsew signal input
rlabel metal2 s 525430 0 525486 800 6 la_data_in[119]
port 167 nsew signal input
rlabel metal2 s 158074 0 158130 800 6 la_data_in[11]
port 168 nsew signal input
rlabel metal2 s 528834 0 528890 800 6 la_data_in[120]
port 169 nsew signal input
rlabel metal2 s 532238 0 532294 800 6 la_data_in[121]
port 170 nsew signal input
rlabel metal2 s 535642 0 535698 800 6 la_data_in[122]
port 171 nsew signal input
rlabel metal2 s 539046 0 539102 800 6 la_data_in[123]
port 172 nsew signal input
rlabel metal2 s 542450 0 542506 800 6 la_data_in[124]
port 173 nsew signal input
rlabel metal2 s 545854 0 545910 800 6 la_data_in[125]
port 174 nsew signal input
rlabel metal2 s 549258 0 549314 800 6 la_data_in[126]
port 175 nsew signal input
rlabel metal2 s 552662 0 552718 800 6 la_data_in[127]
port 176 nsew signal input
rlabel metal2 s 161478 0 161534 800 6 la_data_in[12]
port 177 nsew signal input
rlabel metal2 s 164882 0 164938 800 6 la_data_in[13]
port 178 nsew signal input
rlabel metal2 s 168286 0 168342 800 6 la_data_in[14]
port 179 nsew signal input
rlabel metal2 s 171690 0 171746 800 6 la_data_in[15]
port 180 nsew signal input
rlabel metal2 s 175094 0 175150 800 6 la_data_in[16]
port 181 nsew signal input
rlabel metal2 s 178498 0 178554 800 6 la_data_in[17]
port 182 nsew signal input
rlabel metal2 s 181902 0 181958 800 6 la_data_in[18]
port 183 nsew signal input
rlabel metal2 s 185306 0 185362 800 6 la_data_in[19]
port 184 nsew signal input
rlabel metal2 s 124126 0 124182 800 6 la_data_in[1]
port 185 nsew signal input
rlabel metal2 s 188710 0 188766 800 6 la_data_in[20]
port 186 nsew signal input
rlabel metal2 s 192114 0 192170 800 6 la_data_in[21]
port 187 nsew signal input
rlabel metal2 s 195518 0 195574 800 6 la_data_in[22]
port 188 nsew signal input
rlabel metal2 s 198922 0 198978 800 6 la_data_in[23]
port 189 nsew signal input
rlabel metal2 s 202326 0 202382 800 6 la_data_in[24]
port 190 nsew signal input
rlabel metal2 s 205730 0 205786 800 6 la_data_in[25]
port 191 nsew signal input
rlabel metal2 s 209134 0 209190 800 6 la_data_in[26]
port 192 nsew signal input
rlabel metal2 s 212538 0 212594 800 6 la_data_in[27]
port 193 nsew signal input
rlabel metal2 s 215942 0 215998 800 6 la_data_in[28]
port 194 nsew signal input
rlabel metal2 s 219346 0 219402 800 6 la_data_in[29]
port 195 nsew signal input
rlabel metal2 s 127530 0 127586 800 6 la_data_in[2]
port 196 nsew signal input
rlabel metal2 s 222750 0 222806 800 6 la_data_in[30]
port 197 nsew signal input
rlabel metal2 s 226154 0 226210 800 6 la_data_in[31]
port 198 nsew signal input
rlabel metal2 s 229558 0 229614 800 6 la_data_in[32]
port 199 nsew signal input
rlabel metal2 s 232962 0 233018 800 6 la_data_in[33]
port 200 nsew signal input
rlabel metal2 s 236366 0 236422 800 6 la_data_in[34]
port 201 nsew signal input
rlabel metal2 s 239770 0 239826 800 6 la_data_in[35]
port 202 nsew signal input
rlabel metal2 s 243174 0 243230 800 6 la_data_in[36]
port 203 nsew signal input
rlabel metal2 s 246578 0 246634 800 6 la_data_in[37]
port 204 nsew signal input
rlabel metal2 s 249982 0 250038 800 6 la_data_in[38]
port 205 nsew signal input
rlabel metal2 s 253386 0 253442 800 6 la_data_in[39]
port 206 nsew signal input
rlabel metal2 s 130934 0 130990 800 6 la_data_in[3]
port 207 nsew signal input
rlabel metal2 s 256790 0 256846 800 6 la_data_in[40]
port 208 nsew signal input
rlabel metal2 s 260194 0 260250 800 6 la_data_in[41]
port 209 nsew signal input
rlabel metal2 s 263598 0 263654 800 6 la_data_in[42]
port 210 nsew signal input
rlabel metal2 s 266910 0 266966 800 6 la_data_in[43]
port 211 nsew signal input
rlabel metal2 s 270314 0 270370 800 6 la_data_in[44]
port 212 nsew signal input
rlabel metal2 s 273718 0 273774 800 6 la_data_in[45]
port 213 nsew signal input
rlabel metal2 s 277122 0 277178 800 6 la_data_in[46]
port 214 nsew signal input
rlabel metal2 s 280526 0 280582 800 6 la_data_in[47]
port 215 nsew signal input
rlabel metal2 s 283930 0 283986 800 6 la_data_in[48]
port 216 nsew signal input
rlabel metal2 s 287334 0 287390 800 6 la_data_in[49]
port 217 nsew signal input
rlabel metal2 s 134338 0 134394 800 6 la_data_in[4]
port 218 nsew signal input
rlabel metal2 s 290738 0 290794 800 6 la_data_in[50]
port 219 nsew signal input
rlabel metal2 s 294142 0 294198 800 6 la_data_in[51]
port 220 nsew signal input
rlabel metal2 s 297546 0 297602 800 6 la_data_in[52]
port 221 nsew signal input
rlabel metal2 s 300950 0 301006 800 6 la_data_in[53]
port 222 nsew signal input
rlabel metal2 s 304354 0 304410 800 6 la_data_in[54]
port 223 nsew signal input
rlabel metal2 s 307758 0 307814 800 6 la_data_in[55]
port 224 nsew signal input
rlabel metal2 s 311162 0 311218 800 6 la_data_in[56]
port 225 nsew signal input
rlabel metal2 s 314566 0 314622 800 6 la_data_in[57]
port 226 nsew signal input
rlabel metal2 s 317970 0 318026 800 6 la_data_in[58]
port 227 nsew signal input
rlabel metal2 s 321374 0 321430 800 6 la_data_in[59]
port 228 nsew signal input
rlabel metal2 s 137742 0 137798 800 6 la_data_in[5]
port 229 nsew signal input
rlabel metal2 s 324778 0 324834 800 6 la_data_in[60]
port 230 nsew signal input
rlabel metal2 s 328182 0 328238 800 6 la_data_in[61]
port 231 nsew signal input
rlabel metal2 s 331586 0 331642 800 6 la_data_in[62]
port 232 nsew signal input
rlabel metal2 s 334990 0 335046 800 6 la_data_in[63]
port 233 nsew signal input
rlabel metal2 s 338394 0 338450 800 6 la_data_in[64]
port 234 nsew signal input
rlabel metal2 s 341798 0 341854 800 6 la_data_in[65]
port 235 nsew signal input
rlabel metal2 s 345202 0 345258 800 6 la_data_in[66]
port 236 nsew signal input
rlabel metal2 s 348606 0 348662 800 6 la_data_in[67]
port 237 nsew signal input
rlabel metal2 s 352010 0 352066 800 6 la_data_in[68]
port 238 nsew signal input
rlabel metal2 s 355414 0 355470 800 6 la_data_in[69]
port 239 nsew signal input
rlabel metal2 s 141146 0 141202 800 6 la_data_in[6]
port 240 nsew signal input
rlabel metal2 s 358818 0 358874 800 6 la_data_in[70]
port 241 nsew signal input
rlabel metal2 s 362222 0 362278 800 6 la_data_in[71]
port 242 nsew signal input
rlabel metal2 s 365626 0 365682 800 6 la_data_in[72]
port 243 nsew signal input
rlabel metal2 s 369030 0 369086 800 6 la_data_in[73]
port 244 nsew signal input
rlabel metal2 s 372434 0 372490 800 6 la_data_in[74]
port 245 nsew signal input
rlabel metal2 s 375838 0 375894 800 6 la_data_in[75]
port 246 nsew signal input
rlabel metal2 s 379242 0 379298 800 6 la_data_in[76]
port 247 nsew signal input
rlabel metal2 s 382554 0 382610 800 6 la_data_in[77]
port 248 nsew signal input
rlabel metal2 s 385958 0 386014 800 6 la_data_in[78]
port 249 nsew signal input
rlabel metal2 s 389362 0 389418 800 6 la_data_in[79]
port 250 nsew signal input
rlabel metal2 s 144550 0 144606 800 6 la_data_in[7]
port 251 nsew signal input
rlabel metal2 s 392766 0 392822 800 6 la_data_in[80]
port 252 nsew signal input
rlabel metal2 s 396170 0 396226 800 6 la_data_in[81]
port 253 nsew signal input
rlabel metal2 s 399574 0 399630 800 6 la_data_in[82]
port 254 nsew signal input
rlabel metal2 s 402978 0 403034 800 6 la_data_in[83]
port 255 nsew signal input
rlabel metal2 s 406382 0 406438 800 6 la_data_in[84]
port 256 nsew signal input
rlabel metal2 s 409786 0 409842 800 6 la_data_in[85]
port 257 nsew signal input
rlabel metal2 s 413190 0 413246 800 6 la_data_in[86]
port 258 nsew signal input
rlabel metal2 s 416594 0 416650 800 6 la_data_in[87]
port 259 nsew signal input
rlabel metal2 s 419998 0 420054 800 6 la_data_in[88]
port 260 nsew signal input
rlabel metal2 s 423402 0 423458 800 6 la_data_in[89]
port 261 nsew signal input
rlabel metal2 s 147954 0 148010 800 6 la_data_in[8]
port 262 nsew signal input
rlabel metal2 s 426806 0 426862 800 6 la_data_in[90]
port 263 nsew signal input
rlabel metal2 s 430210 0 430266 800 6 la_data_in[91]
port 264 nsew signal input
rlabel metal2 s 433614 0 433670 800 6 la_data_in[92]
port 265 nsew signal input
rlabel metal2 s 437018 0 437074 800 6 la_data_in[93]
port 266 nsew signal input
rlabel metal2 s 440422 0 440478 800 6 la_data_in[94]
port 267 nsew signal input
rlabel metal2 s 443826 0 443882 800 6 la_data_in[95]
port 268 nsew signal input
rlabel metal2 s 447230 0 447286 800 6 la_data_in[96]
port 269 nsew signal input
rlabel metal2 s 450634 0 450690 800 6 la_data_in[97]
port 270 nsew signal input
rlabel metal2 s 454038 0 454094 800 6 la_data_in[98]
port 271 nsew signal input
rlabel metal2 s 457442 0 457498 800 6 la_data_in[99]
port 272 nsew signal input
rlabel metal2 s 151358 0 151414 800 6 la_data_in[9]
port 273 nsew signal input
rlabel metal2 s 121826 0 121882 800 6 la_data_out[0]
port 274 nsew signal output
rlabel metal2 s 461950 0 462006 800 6 la_data_out[100]
port 275 nsew signal output
rlabel metal2 s 465354 0 465410 800 6 la_data_out[101]
port 276 nsew signal output
rlabel metal2 s 468758 0 468814 800 6 la_data_out[102]
port 277 nsew signal output
rlabel metal2 s 472162 0 472218 800 6 la_data_out[103]
port 278 nsew signal output
rlabel metal2 s 475566 0 475622 800 6 la_data_out[104]
port 279 nsew signal output
rlabel metal2 s 478970 0 479026 800 6 la_data_out[105]
port 280 nsew signal output
rlabel metal2 s 482374 0 482430 800 6 la_data_out[106]
port 281 nsew signal output
rlabel metal2 s 485778 0 485834 800 6 la_data_out[107]
port 282 nsew signal output
rlabel metal2 s 489182 0 489238 800 6 la_data_out[108]
port 283 nsew signal output
rlabel metal2 s 492586 0 492642 800 6 la_data_out[109]
port 284 nsew signal output
rlabel metal2 s 155866 0 155922 800 6 la_data_out[10]
port 285 nsew signal output
rlabel metal2 s 495990 0 496046 800 6 la_data_out[110]
port 286 nsew signal output
rlabel metal2 s 499394 0 499450 800 6 la_data_out[111]
port 287 nsew signal output
rlabel metal2 s 502798 0 502854 800 6 la_data_out[112]
port 288 nsew signal output
rlabel metal2 s 506202 0 506258 800 6 la_data_out[113]
port 289 nsew signal output
rlabel metal2 s 509606 0 509662 800 6 la_data_out[114]
port 290 nsew signal output
rlabel metal2 s 513010 0 513066 800 6 la_data_out[115]
port 291 nsew signal output
rlabel metal2 s 516414 0 516470 800 6 la_data_out[116]
port 292 nsew signal output
rlabel metal2 s 519818 0 519874 800 6 la_data_out[117]
port 293 nsew signal output
rlabel metal2 s 523222 0 523278 800 6 la_data_out[118]
port 294 nsew signal output
rlabel metal2 s 526626 0 526682 800 6 la_data_out[119]
port 295 nsew signal output
rlabel metal2 s 159270 0 159326 800 6 la_data_out[11]
port 296 nsew signal output
rlabel metal2 s 530030 0 530086 800 6 la_data_out[120]
port 297 nsew signal output
rlabel metal2 s 533342 0 533398 800 6 la_data_out[121]
port 298 nsew signal output
rlabel metal2 s 536746 0 536802 800 6 la_data_out[122]
port 299 nsew signal output
rlabel metal2 s 540150 0 540206 800 6 la_data_out[123]
port 300 nsew signal output
rlabel metal2 s 543554 0 543610 800 6 la_data_out[124]
port 301 nsew signal output
rlabel metal2 s 546958 0 547014 800 6 la_data_out[125]
port 302 nsew signal output
rlabel metal2 s 550362 0 550418 800 6 la_data_out[126]
port 303 nsew signal output
rlabel metal2 s 553766 0 553822 800 6 la_data_out[127]
port 304 nsew signal output
rlabel metal2 s 162674 0 162730 800 6 la_data_out[12]
port 305 nsew signal output
rlabel metal2 s 166078 0 166134 800 6 la_data_out[13]
port 306 nsew signal output
rlabel metal2 s 169482 0 169538 800 6 la_data_out[14]
port 307 nsew signal output
rlabel metal2 s 172886 0 172942 800 6 la_data_out[15]
port 308 nsew signal output
rlabel metal2 s 176290 0 176346 800 6 la_data_out[16]
port 309 nsew signal output
rlabel metal2 s 179694 0 179750 800 6 la_data_out[17]
port 310 nsew signal output
rlabel metal2 s 183098 0 183154 800 6 la_data_out[18]
port 311 nsew signal output
rlabel metal2 s 186502 0 186558 800 6 la_data_out[19]
port 312 nsew signal output
rlabel metal2 s 125230 0 125286 800 6 la_data_out[1]
port 313 nsew signal output
rlabel metal2 s 189906 0 189962 800 6 la_data_out[20]
port 314 nsew signal output
rlabel metal2 s 193218 0 193274 800 6 la_data_out[21]
port 315 nsew signal output
rlabel metal2 s 196622 0 196678 800 6 la_data_out[22]
port 316 nsew signal output
rlabel metal2 s 200026 0 200082 800 6 la_data_out[23]
port 317 nsew signal output
rlabel metal2 s 203430 0 203486 800 6 la_data_out[24]
port 318 nsew signal output
rlabel metal2 s 206834 0 206890 800 6 la_data_out[25]
port 319 nsew signal output
rlabel metal2 s 210238 0 210294 800 6 la_data_out[26]
port 320 nsew signal output
rlabel metal2 s 213642 0 213698 800 6 la_data_out[27]
port 321 nsew signal output
rlabel metal2 s 217046 0 217102 800 6 la_data_out[28]
port 322 nsew signal output
rlabel metal2 s 220450 0 220506 800 6 la_data_out[29]
port 323 nsew signal output
rlabel metal2 s 128634 0 128690 800 6 la_data_out[2]
port 324 nsew signal output
rlabel metal2 s 223854 0 223910 800 6 la_data_out[30]
port 325 nsew signal output
rlabel metal2 s 227258 0 227314 800 6 la_data_out[31]
port 326 nsew signal output
rlabel metal2 s 230662 0 230718 800 6 la_data_out[32]
port 327 nsew signal output
rlabel metal2 s 234066 0 234122 800 6 la_data_out[33]
port 328 nsew signal output
rlabel metal2 s 237470 0 237526 800 6 la_data_out[34]
port 329 nsew signal output
rlabel metal2 s 240874 0 240930 800 6 la_data_out[35]
port 330 nsew signal output
rlabel metal2 s 244278 0 244334 800 6 la_data_out[36]
port 331 nsew signal output
rlabel metal2 s 247682 0 247738 800 6 la_data_out[37]
port 332 nsew signal output
rlabel metal2 s 251086 0 251142 800 6 la_data_out[38]
port 333 nsew signal output
rlabel metal2 s 254490 0 254546 800 6 la_data_out[39]
port 334 nsew signal output
rlabel metal2 s 132038 0 132094 800 6 la_data_out[3]
port 335 nsew signal output
rlabel metal2 s 257894 0 257950 800 6 la_data_out[40]
port 336 nsew signal output
rlabel metal2 s 261298 0 261354 800 6 la_data_out[41]
port 337 nsew signal output
rlabel metal2 s 264702 0 264758 800 6 la_data_out[42]
port 338 nsew signal output
rlabel metal2 s 268106 0 268162 800 6 la_data_out[43]
port 339 nsew signal output
rlabel metal2 s 271510 0 271566 800 6 la_data_out[44]
port 340 nsew signal output
rlabel metal2 s 274914 0 274970 800 6 la_data_out[45]
port 341 nsew signal output
rlabel metal2 s 278318 0 278374 800 6 la_data_out[46]
port 342 nsew signal output
rlabel metal2 s 281722 0 281778 800 6 la_data_out[47]
port 343 nsew signal output
rlabel metal2 s 285126 0 285182 800 6 la_data_out[48]
port 344 nsew signal output
rlabel metal2 s 288530 0 288586 800 6 la_data_out[49]
port 345 nsew signal output
rlabel metal2 s 135442 0 135498 800 6 la_data_out[4]
port 346 nsew signal output
rlabel metal2 s 291934 0 291990 800 6 la_data_out[50]
port 347 nsew signal output
rlabel metal2 s 295338 0 295394 800 6 la_data_out[51]
port 348 nsew signal output
rlabel metal2 s 298742 0 298798 800 6 la_data_out[52]
port 349 nsew signal output
rlabel metal2 s 302146 0 302202 800 6 la_data_out[53]
port 350 nsew signal output
rlabel metal2 s 305458 0 305514 800 6 la_data_out[54]
port 351 nsew signal output
rlabel metal2 s 308862 0 308918 800 6 la_data_out[55]
port 352 nsew signal output
rlabel metal2 s 312266 0 312322 800 6 la_data_out[56]
port 353 nsew signal output
rlabel metal2 s 315670 0 315726 800 6 la_data_out[57]
port 354 nsew signal output
rlabel metal2 s 319074 0 319130 800 6 la_data_out[58]
port 355 nsew signal output
rlabel metal2 s 322478 0 322534 800 6 la_data_out[59]
port 356 nsew signal output
rlabel metal2 s 138846 0 138902 800 6 la_data_out[5]
port 357 nsew signal output
rlabel metal2 s 325882 0 325938 800 6 la_data_out[60]
port 358 nsew signal output
rlabel metal2 s 329286 0 329342 800 6 la_data_out[61]
port 359 nsew signal output
rlabel metal2 s 332690 0 332746 800 6 la_data_out[62]
port 360 nsew signal output
rlabel metal2 s 336094 0 336150 800 6 la_data_out[63]
port 361 nsew signal output
rlabel metal2 s 339498 0 339554 800 6 la_data_out[64]
port 362 nsew signal output
rlabel metal2 s 342902 0 342958 800 6 la_data_out[65]
port 363 nsew signal output
rlabel metal2 s 346306 0 346362 800 6 la_data_out[66]
port 364 nsew signal output
rlabel metal2 s 349710 0 349766 800 6 la_data_out[67]
port 365 nsew signal output
rlabel metal2 s 353114 0 353170 800 6 la_data_out[68]
port 366 nsew signal output
rlabel metal2 s 356518 0 356574 800 6 la_data_out[69]
port 367 nsew signal output
rlabel metal2 s 142250 0 142306 800 6 la_data_out[6]
port 368 nsew signal output
rlabel metal2 s 359922 0 359978 800 6 la_data_out[70]
port 369 nsew signal output
rlabel metal2 s 363326 0 363382 800 6 la_data_out[71]
port 370 nsew signal output
rlabel metal2 s 366730 0 366786 800 6 la_data_out[72]
port 371 nsew signal output
rlabel metal2 s 370134 0 370190 800 6 la_data_out[73]
port 372 nsew signal output
rlabel metal2 s 373538 0 373594 800 6 la_data_out[74]
port 373 nsew signal output
rlabel metal2 s 376942 0 376998 800 6 la_data_out[75]
port 374 nsew signal output
rlabel metal2 s 380346 0 380402 800 6 la_data_out[76]
port 375 nsew signal output
rlabel metal2 s 383750 0 383806 800 6 la_data_out[77]
port 376 nsew signal output
rlabel metal2 s 387154 0 387210 800 6 la_data_out[78]
port 377 nsew signal output
rlabel metal2 s 390558 0 390614 800 6 la_data_out[79]
port 378 nsew signal output
rlabel metal2 s 145654 0 145710 800 6 la_data_out[7]
port 379 nsew signal output
rlabel metal2 s 393962 0 394018 800 6 la_data_out[80]
port 380 nsew signal output
rlabel metal2 s 397366 0 397422 800 6 la_data_out[81]
port 381 nsew signal output
rlabel metal2 s 400770 0 400826 800 6 la_data_out[82]
port 382 nsew signal output
rlabel metal2 s 404174 0 404230 800 6 la_data_out[83]
port 383 nsew signal output
rlabel metal2 s 407578 0 407634 800 6 la_data_out[84]
port 384 nsew signal output
rlabel metal2 s 410982 0 411038 800 6 la_data_out[85]
port 385 nsew signal output
rlabel metal2 s 414386 0 414442 800 6 la_data_out[86]
port 386 nsew signal output
rlabel metal2 s 417698 0 417754 800 6 la_data_out[87]
port 387 nsew signal output
rlabel metal2 s 421102 0 421158 800 6 la_data_out[88]
port 388 nsew signal output
rlabel metal2 s 424506 0 424562 800 6 la_data_out[89]
port 389 nsew signal output
rlabel metal2 s 149058 0 149114 800 6 la_data_out[8]
port 390 nsew signal output
rlabel metal2 s 427910 0 427966 800 6 la_data_out[90]
port 391 nsew signal output
rlabel metal2 s 431314 0 431370 800 6 la_data_out[91]
port 392 nsew signal output
rlabel metal2 s 434718 0 434774 800 6 la_data_out[92]
port 393 nsew signal output
rlabel metal2 s 438122 0 438178 800 6 la_data_out[93]
port 394 nsew signal output
rlabel metal2 s 441526 0 441582 800 6 la_data_out[94]
port 395 nsew signal output
rlabel metal2 s 444930 0 444986 800 6 la_data_out[95]
port 396 nsew signal output
rlabel metal2 s 448334 0 448390 800 6 la_data_out[96]
port 397 nsew signal output
rlabel metal2 s 451738 0 451794 800 6 la_data_out[97]
port 398 nsew signal output
rlabel metal2 s 455142 0 455198 800 6 la_data_out[98]
port 399 nsew signal output
rlabel metal2 s 458546 0 458602 800 6 la_data_out[99]
port 400 nsew signal output
rlabel metal2 s 152462 0 152518 800 6 la_data_out[9]
port 401 nsew signal output
rlabel metal2 s 122930 0 122986 800 6 la_oen[0]
port 402 nsew signal input
rlabel metal2 s 463054 0 463110 800 6 la_oen[100]
port 403 nsew signal input
rlabel metal2 s 466458 0 466514 800 6 la_oen[101]
port 404 nsew signal input
rlabel metal2 s 469862 0 469918 800 6 la_oen[102]
port 405 nsew signal input
rlabel metal2 s 473266 0 473322 800 6 la_oen[103]
port 406 nsew signal input
rlabel metal2 s 476670 0 476726 800 6 la_oen[104]
port 407 nsew signal input
rlabel metal2 s 480074 0 480130 800 6 la_oen[105]
port 408 nsew signal input
rlabel metal2 s 483478 0 483534 800 6 la_oen[106]
port 409 nsew signal input
rlabel metal2 s 486882 0 486938 800 6 la_oen[107]
port 410 nsew signal input
rlabel metal2 s 490286 0 490342 800 6 la_oen[108]
port 411 nsew signal input
rlabel metal2 s 493690 0 493746 800 6 la_oen[109]
port 412 nsew signal input
rlabel metal2 s 156970 0 157026 800 6 la_oen[10]
port 413 nsew signal input
rlabel metal2 s 497094 0 497150 800 6 la_oen[110]
port 414 nsew signal input
rlabel metal2 s 500498 0 500554 800 6 la_oen[111]
port 415 nsew signal input
rlabel metal2 s 503902 0 503958 800 6 la_oen[112]
port 416 nsew signal input
rlabel metal2 s 507306 0 507362 800 6 la_oen[113]
port 417 nsew signal input
rlabel metal2 s 510710 0 510766 800 6 la_oen[114]
port 418 nsew signal input
rlabel metal2 s 514114 0 514170 800 6 la_oen[115]
port 419 nsew signal input
rlabel metal2 s 517518 0 517574 800 6 la_oen[116]
port 420 nsew signal input
rlabel metal2 s 520922 0 520978 800 6 la_oen[117]
port 421 nsew signal input
rlabel metal2 s 524326 0 524382 800 6 la_oen[118]
port 422 nsew signal input
rlabel metal2 s 527730 0 527786 800 6 la_oen[119]
port 423 nsew signal input
rlabel metal2 s 160374 0 160430 800 6 la_oen[11]
port 424 nsew signal input
rlabel metal2 s 531134 0 531190 800 6 la_oen[120]
port 425 nsew signal input
rlabel metal2 s 534538 0 534594 800 6 la_oen[121]
port 426 nsew signal input
rlabel metal2 s 537942 0 537998 800 6 la_oen[122]
port 427 nsew signal input
rlabel metal2 s 541346 0 541402 800 6 la_oen[123]
port 428 nsew signal input
rlabel metal2 s 544750 0 544806 800 6 la_oen[124]
port 429 nsew signal input
rlabel metal2 s 548154 0 548210 800 6 la_oen[125]
port 430 nsew signal input
rlabel metal2 s 551558 0 551614 800 6 la_oen[126]
port 431 nsew signal input
rlabel metal2 s 554962 0 555018 800 6 la_oen[127]
port 432 nsew signal input
rlabel metal2 s 163778 0 163834 800 6 la_oen[12]
port 433 nsew signal input
rlabel metal2 s 167182 0 167238 800 6 la_oen[13]
port 434 nsew signal input
rlabel metal2 s 170586 0 170642 800 6 la_oen[14]
port 435 nsew signal input
rlabel metal2 s 173990 0 174046 800 6 la_oen[15]
port 436 nsew signal input
rlabel metal2 s 177394 0 177450 800 6 la_oen[16]
port 437 nsew signal input
rlabel metal2 s 180798 0 180854 800 6 la_oen[17]
port 438 nsew signal input
rlabel metal2 s 184202 0 184258 800 6 la_oen[18]
port 439 nsew signal input
rlabel metal2 s 187606 0 187662 800 6 la_oen[19]
port 440 nsew signal input
rlabel metal2 s 126334 0 126390 800 6 la_oen[1]
port 441 nsew signal input
rlabel metal2 s 191010 0 191066 800 6 la_oen[20]
port 442 nsew signal input
rlabel metal2 s 194414 0 194470 800 6 la_oen[21]
port 443 nsew signal input
rlabel metal2 s 197818 0 197874 800 6 la_oen[22]
port 444 nsew signal input
rlabel metal2 s 201222 0 201278 800 6 la_oen[23]
port 445 nsew signal input
rlabel metal2 s 204626 0 204682 800 6 la_oen[24]
port 446 nsew signal input
rlabel metal2 s 208030 0 208086 800 6 la_oen[25]
port 447 nsew signal input
rlabel metal2 s 211434 0 211490 800 6 la_oen[26]
port 448 nsew signal input
rlabel metal2 s 214838 0 214894 800 6 la_oen[27]
port 449 nsew signal input
rlabel metal2 s 218242 0 218298 800 6 la_oen[28]
port 450 nsew signal input
rlabel metal2 s 221646 0 221702 800 6 la_oen[29]
port 451 nsew signal input
rlabel metal2 s 129738 0 129794 800 6 la_oen[2]
port 452 nsew signal input
rlabel metal2 s 225050 0 225106 800 6 la_oen[30]
port 453 nsew signal input
rlabel metal2 s 228362 0 228418 800 6 la_oen[31]
port 454 nsew signal input
rlabel metal2 s 231766 0 231822 800 6 la_oen[32]
port 455 nsew signal input
rlabel metal2 s 235170 0 235226 800 6 la_oen[33]
port 456 nsew signal input
rlabel metal2 s 238574 0 238630 800 6 la_oen[34]
port 457 nsew signal input
rlabel metal2 s 241978 0 242034 800 6 la_oen[35]
port 458 nsew signal input
rlabel metal2 s 245382 0 245438 800 6 la_oen[36]
port 459 nsew signal input
rlabel metal2 s 248786 0 248842 800 6 la_oen[37]
port 460 nsew signal input
rlabel metal2 s 252190 0 252246 800 6 la_oen[38]
port 461 nsew signal input
rlabel metal2 s 255594 0 255650 800 6 la_oen[39]
port 462 nsew signal input
rlabel metal2 s 133142 0 133198 800 6 la_oen[3]
port 463 nsew signal input
rlabel metal2 s 258998 0 259054 800 6 la_oen[40]
port 464 nsew signal input
rlabel metal2 s 262402 0 262458 800 6 la_oen[41]
port 465 nsew signal input
rlabel metal2 s 265806 0 265862 800 6 la_oen[42]
port 466 nsew signal input
rlabel metal2 s 269210 0 269266 800 6 la_oen[43]
port 467 nsew signal input
rlabel metal2 s 272614 0 272670 800 6 la_oen[44]
port 468 nsew signal input
rlabel metal2 s 276018 0 276074 800 6 la_oen[45]
port 469 nsew signal input
rlabel metal2 s 279422 0 279478 800 6 la_oen[46]
port 470 nsew signal input
rlabel metal2 s 282826 0 282882 800 6 la_oen[47]
port 471 nsew signal input
rlabel metal2 s 286230 0 286286 800 6 la_oen[48]
port 472 nsew signal input
rlabel metal2 s 289634 0 289690 800 6 la_oen[49]
port 473 nsew signal input
rlabel metal2 s 136546 0 136602 800 6 la_oen[4]
port 474 nsew signal input
rlabel metal2 s 293038 0 293094 800 6 la_oen[50]
port 475 nsew signal input
rlabel metal2 s 296442 0 296498 800 6 la_oen[51]
port 476 nsew signal input
rlabel metal2 s 299846 0 299902 800 6 la_oen[52]
port 477 nsew signal input
rlabel metal2 s 303250 0 303306 800 6 la_oen[53]
port 478 nsew signal input
rlabel metal2 s 306654 0 306710 800 6 la_oen[54]
port 479 nsew signal input
rlabel metal2 s 310058 0 310114 800 6 la_oen[55]
port 480 nsew signal input
rlabel metal2 s 313462 0 313518 800 6 la_oen[56]
port 481 nsew signal input
rlabel metal2 s 316866 0 316922 800 6 la_oen[57]
port 482 nsew signal input
rlabel metal2 s 320270 0 320326 800 6 la_oen[58]
port 483 nsew signal input
rlabel metal2 s 323674 0 323730 800 6 la_oen[59]
port 484 nsew signal input
rlabel metal2 s 139950 0 140006 800 6 la_oen[5]
port 485 nsew signal input
rlabel metal2 s 327078 0 327134 800 6 la_oen[60]
port 486 nsew signal input
rlabel metal2 s 330482 0 330538 800 6 la_oen[61]
port 487 nsew signal input
rlabel metal2 s 333886 0 333942 800 6 la_oen[62]
port 488 nsew signal input
rlabel metal2 s 337290 0 337346 800 6 la_oen[63]
port 489 nsew signal input
rlabel metal2 s 340694 0 340750 800 6 la_oen[64]
port 490 nsew signal input
rlabel metal2 s 344006 0 344062 800 6 la_oen[65]
port 491 nsew signal input
rlabel metal2 s 347410 0 347466 800 6 la_oen[66]
port 492 nsew signal input
rlabel metal2 s 350814 0 350870 800 6 la_oen[67]
port 493 nsew signal input
rlabel metal2 s 354218 0 354274 800 6 la_oen[68]
port 494 nsew signal input
rlabel metal2 s 357622 0 357678 800 6 la_oen[69]
port 495 nsew signal input
rlabel metal2 s 143354 0 143410 800 6 la_oen[6]
port 496 nsew signal input
rlabel metal2 s 361026 0 361082 800 6 la_oen[70]
port 497 nsew signal input
rlabel metal2 s 364430 0 364486 800 6 la_oen[71]
port 498 nsew signal input
rlabel metal2 s 367834 0 367890 800 6 la_oen[72]
port 499 nsew signal input
rlabel metal2 s 371238 0 371294 800 6 la_oen[73]
port 500 nsew signal input
rlabel metal2 s 374642 0 374698 800 6 la_oen[74]
port 501 nsew signal input
rlabel metal2 s 378046 0 378102 800 6 la_oen[75]
port 502 nsew signal input
rlabel metal2 s 381450 0 381506 800 6 la_oen[76]
port 503 nsew signal input
rlabel metal2 s 384854 0 384910 800 6 la_oen[77]
port 504 nsew signal input
rlabel metal2 s 388258 0 388314 800 6 la_oen[78]
port 505 nsew signal input
rlabel metal2 s 391662 0 391718 800 6 la_oen[79]
port 506 nsew signal input
rlabel metal2 s 146758 0 146814 800 6 la_oen[7]
port 507 nsew signal input
rlabel metal2 s 395066 0 395122 800 6 la_oen[80]
port 508 nsew signal input
rlabel metal2 s 398470 0 398526 800 6 la_oen[81]
port 509 nsew signal input
rlabel metal2 s 401874 0 401930 800 6 la_oen[82]
port 510 nsew signal input
rlabel metal2 s 405278 0 405334 800 6 la_oen[83]
port 511 nsew signal input
rlabel metal2 s 408682 0 408738 800 6 la_oen[84]
port 512 nsew signal input
rlabel metal2 s 412086 0 412142 800 6 la_oen[85]
port 513 nsew signal input
rlabel metal2 s 415490 0 415546 800 6 la_oen[86]
port 514 nsew signal input
rlabel metal2 s 418894 0 418950 800 6 la_oen[87]
port 515 nsew signal input
rlabel metal2 s 422298 0 422354 800 6 la_oen[88]
port 516 nsew signal input
rlabel metal2 s 425702 0 425758 800 6 la_oen[89]
port 517 nsew signal input
rlabel metal2 s 150162 0 150218 800 6 la_oen[8]
port 518 nsew signal input
rlabel metal2 s 429106 0 429162 800 6 la_oen[90]
port 519 nsew signal input
rlabel metal2 s 432510 0 432566 800 6 la_oen[91]
port 520 nsew signal input
rlabel metal2 s 435914 0 435970 800 6 la_oen[92]
port 521 nsew signal input
rlabel metal2 s 439318 0 439374 800 6 la_oen[93]
port 522 nsew signal input
rlabel metal2 s 442722 0 442778 800 6 la_oen[94]
port 523 nsew signal input
rlabel metal2 s 446126 0 446182 800 6 la_oen[95]
port 524 nsew signal input
rlabel metal2 s 449530 0 449586 800 6 la_oen[96]
port 525 nsew signal input
rlabel metal2 s 452934 0 452990 800 6 la_oen[97]
port 526 nsew signal input
rlabel metal2 s 456246 0 456302 800 6 la_oen[98]
port 527 nsew signal input
rlabel metal2 s 459650 0 459706 800 6 la_oen[99]
port 528 nsew signal input
rlabel metal2 s 153566 0 153622 800 6 la_oen[9]
port 529 nsew signal input
rlabel metal2 s 556066 0 556122 800 6 user_clock2
port 530 nsew signal input
rlabel metal2 s 570 0 626 800 6 wb_clk_i
port 531 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wb_rst_i
port 532 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 wbs_ack_o
port 533 nsew signal output
rlabel metal2 s 7286 0 7342 800 6 wbs_adr_i[0]
port 534 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 wbs_adr_i[10]
port 535 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 wbs_adr_i[11]
port 536 nsew signal input
rlabel metal2 s 52642 0 52698 800 6 wbs_adr_i[12]
port 537 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 wbs_adr_i[13]
port 538 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 wbs_adr_i[14]
port 539 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 wbs_adr_i[15]
port 540 nsew signal input
rlabel metal2 s 66258 0 66314 800 6 wbs_adr_i[16]
port 541 nsew signal input
rlabel metal2 s 69662 0 69718 800 6 wbs_adr_i[17]
port 542 nsew signal input
rlabel metal2 s 73066 0 73122 800 6 wbs_adr_i[18]
port 543 nsew signal input
rlabel metal2 s 76470 0 76526 800 6 wbs_adr_i[19]
port 544 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 wbs_adr_i[1]
port 545 nsew signal input
rlabel metal2 s 79874 0 79930 800 6 wbs_adr_i[20]
port 546 nsew signal input
rlabel metal2 s 83278 0 83334 800 6 wbs_adr_i[21]
port 547 nsew signal input
rlabel metal2 s 86682 0 86738 800 6 wbs_adr_i[22]
port 548 nsew signal input
rlabel metal2 s 90086 0 90142 800 6 wbs_adr_i[23]
port 549 nsew signal input
rlabel metal2 s 93490 0 93546 800 6 wbs_adr_i[24]
port 550 nsew signal input
rlabel metal2 s 96894 0 96950 800 6 wbs_adr_i[25]
port 551 nsew signal input
rlabel metal2 s 100298 0 100354 800 6 wbs_adr_i[26]
port 552 nsew signal input
rlabel metal2 s 103702 0 103758 800 6 wbs_adr_i[27]
port 553 nsew signal input
rlabel metal2 s 107106 0 107162 800 6 wbs_adr_i[28]
port 554 nsew signal input
rlabel metal2 s 110510 0 110566 800 6 wbs_adr_i[29]
port 555 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 wbs_adr_i[2]
port 556 nsew signal input
rlabel metal2 s 113914 0 113970 800 6 wbs_adr_i[30]
port 557 nsew signal input
rlabel metal2 s 117318 0 117374 800 6 wbs_adr_i[31]
port 558 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 wbs_adr_i[3]
port 559 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 wbs_adr_i[4]
port 560 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 wbs_adr_i[5]
port 561 nsew signal input
rlabel metal2 s 32310 0 32366 800 6 wbs_adr_i[6]
port 562 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 wbs_adr_i[7]
port 563 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 wbs_adr_i[8]
port 564 nsew signal input
rlabel metal2 s 42430 0 42486 800 6 wbs_adr_i[9]
port 565 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 wbs_cyc_i
port 566 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_dat_i[0]
port 567 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 wbs_dat_i[10]
port 568 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 wbs_dat_i[11]
port 569 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 wbs_dat_i[12]
port 570 nsew signal input
rlabel metal2 s 57242 0 57298 800 6 wbs_dat_i[13]
port 571 nsew signal input
rlabel metal2 s 60646 0 60702 800 6 wbs_dat_i[14]
port 572 nsew signal input
rlabel metal2 s 64050 0 64106 800 6 wbs_dat_i[15]
port 573 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 wbs_dat_i[16]
port 574 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 wbs_dat_i[17]
port 575 nsew signal input
rlabel metal2 s 74262 0 74318 800 6 wbs_dat_i[18]
port 576 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 wbs_dat_i[19]
port 577 nsew signal input
rlabel metal2 s 12990 0 13046 800 6 wbs_dat_i[1]
port 578 nsew signal input
rlabel metal2 s 80978 0 81034 800 6 wbs_dat_i[20]
port 579 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 wbs_dat_i[21]
port 580 nsew signal input
rlabel metal2 s 87786 0 87842 800 6 wbs_dat_i[22]
port 581 nsew signal input
rlabel metal2 s 91190 0 91246 800 6 wbs_dat_i[23]
port 582 nsew signal input
rlabel metal2 s 94594 0 94650 800 6 wbs_dat_i[24]
port 583 nsew signal input
rlabel metal2 s 97998 0 98054 800 6 wbs_dat_i[25]
port 584 nsew signal input
rlabel metal2 s 101402 0 101458 800 6 wbs_dat_i[26]
port 585 nsew signal input
rlabel metal2 s 104806 0 104862 800 6 wbs_dat_i[27]
port 586 nsew signal input
rlabel metal2 s 108210 0 108266 800 6 wbs_dat_i[28]
port 587 nsew signal input
rlabel metal2 s 111614 0 111670 800 6 wbs_dat_i[29]
port 588 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 wbs_dat_i[2]
port 589 nsew signal input
rlabel metal2 s 115018 0 115074 800 6 wbs_dat_i[30]
port 590 nsew signal input
rlabel metal2 s 118422 0 118478 800 6 wbs_dat_i[31]
port 591 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 wbs_dat_i[3]
port 592 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 wbs_dat_i[4]
port 593 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 wbs_dat_i[5]
port 594 nsew signal input
rlabel metal2 s 33414 0 33470 800 6 wbs_dat_i[6]
port 595 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 wbs_dat_i[7]
port 596 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 wbs_dat_i[8]
port 597 nsew signal input
rlabel metal2 s 43626 0 43682 800 6 wbs_dat_i[9]
port 598 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_dat_o[0]
port 599 nsew signal output
rlabel metal2 s 48134 0 48190 800 6 wbs_dat_o[10]
port 600 nsew signal output
rlabel metal2 s 51538 0 51594 800 6 wbs_dat_o[11]
port 601 nsew signal output
rlabel metal2 s 54942 0 54998 800 6 wbs_dat_o[12]
port 602 nsew signal output
rlabel metal2 s 58346 0 58402 800 6 wbs_dat_o[13]
port 603 nsew signal output
rlabel metal2 s 61750 0 61806 800 6 wbs_dat_o[14]
port 604 nsew signal output
rlabel metal2 s 65154 0 65210 800 6 wbs_dat_o[15]
port 605 nsew signal output
rlabel metal2 s 68558 0 68614 800 6 wbs_dat_o[16]
port 606 nsew signal output
rlabel metal2 s 71962 0 72018 800 6 wbs_dat_o[17]
port 607 nsew signal output
rlabel metal2 s 75366 0 75422 800 6 wbs_dat_o[18]
port 608 nsew signal output
rlabel metal2 s 78770 0 78826 800 6 wbs_dat_o[19]
port 609 nsew signal output
rlabel metal2 s 14094 0 14150 800 6 wbs_dat_o[1]
port 610 nsew signal output
rlabel metal2 s 82174 0 82230 800 6 wbs_dat_o[20]
port 611 nsew signal output
rlabel metal2 s 85578 0 85634 800 6 wbs_dat_o[21]
port 612 nsew signal output
rlabel metal2 s 88982 0 89038 800 6 wbs_dat_o[22]
port 613 nsew signal output
rlabel metal2 s 92386 0 92442 800 6 wbs_dat_o[23]
port 614 nsew signal output
rlabel metal2 s 95790 0 95846 800 6 wbs_dat_o[24]
port 615 nsew signal output
rlabel metal2 s 99194 0 99250 800 6 wbs_dat_o[25]
port 616 nsew signal output
rlabel metal2 s 102598 0 102654 800 6 wbs_dat_o[26]
port 617 nsew signal output
rlabel metal2 s 106002 0 106058 800 6 wbs_dat_o[27]
port 618 nsew signal output
rlabel metal2 s 109406 0 109462 800 6 wbs_dat_o[28]
port 619 nsew signal output
rlabel metal2 s 112810 0 112866 800 6 wbs_dat_o[29]
port 620 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 wbs_dat_o[2]
port 621 nsew signal output
rlabel metal2 s 116122 0 116178 800 6 wbs_dat_o[30]
port 622 nsew signal output
rlabel metal2 s 119526 0 119582 800 6 wbs_dat_o[31]
port 623 nsew signal output
rlabel metal2 s 23202 0 23258 800 6 wbs_dat_o[3]
port 624 nsew signal output
rlabel metal2 s 27710 0 27766 800 6 wbs_dat_o[4]
port 625 nsew signal output
rlabel metal2 s 31114 0 31170 800 6 wbs_dat_o[5]
port 626 nsew signal output
rlabel metal2 s 34518 0 34574 800 6 wbs_dat_o[6]
port 627 nsew signal output
rlabel metal2 s 37922 0 37978 800 6 wbs_dat_o[7]
port 628 nsew signal output
rlabel metal2 s 41326 0 41382 800 6 wbs_dat_o[8]
port 629 nsew signal output
rlabel metal2 s 44730 0 44786 800 6 wbs_dat_o[9]
port 630 nsew signal output
rlabel metal2 s 10690 0 10746 800 6 wbs_sel_i[0]
port 631 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 wbs_sel_i[1]
port 632 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 wbs_sel_i[2]
port 633 nsew signal input
rlabel metal2 s 24306 0 24362 800 6 wbs_sel_i[3]
port 634 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 wbs_stb_i
port 635 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wbs_we_i
port 636 nsew signal input
rlabel metal4 s 557168 2128 557488 685488 6 VPWR
port 637 nsew power bidirectional
rlabel metal4 s 526448 2128 526768 685488 6 VPWR
port 638 nsew power bidirectional
rlabel metal4 s 495728 2128 496048 685488 6 VPWR
port 639 nsew power bidirectional
rlabel metal4 s 465008 2128 465328 685488 6 VPWR
port 640 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 685488 6 VPWR
port 641 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 685488 6 VPWR
port 642 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 685488 6 VPWR
port 643 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 685488 6 VPWR
port 644 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 685488 6 VPWR
port 645 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 685488 6 VPWR
port 646 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 685488 6 VPWR
port 647 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 685488 6 VPWR
port 648 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 685488 6 VPWR
port 649 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 685488 6 VPWR
port 650 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 685488 6 VPWR
port 651 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 685488 6 VPWR
port 652 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 685488 6 VPWR
port 653 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 685488 6 VPWR
port 654 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 685488 6 VPWR
port 655 nsew power bidirectional
rlabel metal4 s 541808 2128 542128 685488 6 VGND
port 656 nsew ground bidirectional
rlabel metal4 s 511088 2128 511408 685488 6 VGND
port 657 nsew ground bidirectional
rlabel metal4 s 480368 2128 480688 685488 6 VGND
port 658 nsew ground bidirectional
rlabel metal4 s 449648 2128 449968 685488 6 VGND
port 659 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 685488 6 VGND
port 660 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 685488 6 VGND
port 661 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 685488 6 VGND
port 662 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 685488 6 VGND
port 663 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 685488 6 VGND
port 664 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 685488 6 VGND
port 665 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 685488 6 VGND
port 666 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 685488 6 VGND
port 667 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 685488 6 VGND
port 668 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 685488 6 VGND
port 669 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 685488 6 VGND
port 670 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 685488 6 VGND
port 671 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 685488 6 VGND
port 672 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 685488 6 VGND
port 673 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 568000 688000
string LEFview TRUE
<< end >>

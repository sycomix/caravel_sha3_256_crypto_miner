magic
tech sky130A
magscale 1 2
timestamp 1608594439
<< obsli1 >>
rect 1104 2159 566812 685457
<< obsm1 >>
rect 14 1232 566812 685488
<< metal2 >>
rect 2318 687200 2374 688000
rect 7010 687200 7066 688000
rect 11702 687200 11758 688000
rect 16486 687200 16542 688000
rect 21178 687200 21234 688000
rect 25962 687200 26018 688000
rect 30654 687200 30710 688000
rect 35438 687200 35494 688000
rect 40130 687200 40186 688000
rect 44914 687200 44970 688000
rect 49606 687200 49662 688000
rect 54298 687200 54354 688000
rect 59082 687200 59138 688000
rect 63774 687200 63830 688000
rect 68558 687200 68614 688000
rect 73250 687200 73306 688000
rect 78034 687200 78090 688000
rect 82726 687200 82782 688000
rect 87510 687200 87566 688000
rect 92202 687200 92258 688000
rect 96986 687200 97042 688000
rect 101678 687200 101734 688000
rect 106370 687200 106426 688000
rect 111154 687200 111210 688000
rect 115846 687200 115902 688000
rect 120630 687200 120686 688000
rect 125322 687200 125378 688000
rect 130106 687200 130162 688000
rect 134798 687200 134854 688000
rect 139582 687200 139638 688000
rect 144274 687200 144330 688000
rect 148966 687200 149022 688000
rect 153750 687200 153806 688000
rect 158442 687200 158498 688000
rect 163226 687200 163282 688000
rect 167918 687200 167974 688000
rect 172702 687200 172758 688000
rect 177394 687200 177450 688000
rect 182178 687200 182234 688000
rect 186870 687200 186926 688000
rect 191654 687200 191710 688000
rect 196346 687200 196402 688000
rect 201038 687200 201094 688000
rect 205822 687200 205878 688000
rect 210514 687200 210570 688000
rect 215298 687200 215354 688000
rect 219990 687200 220046 688000
rect 224774 687200 224830 688000
rect 229466 687200 229522 688000
rect 234250 687200 234306 688000
rect 238942 687200 238998 688000
rect 243634 687200 243690 688000
rect 248418 687200 248474 688000
rect 253110 687200 253166 688000
rect 257894 687200 257950 688000
rect 262586 687200 262642 688000
rect 267370 687200 267426 688000
rect 272062 687200 272118 688000
rect 276846 687200 276902 688000
rect 281538 687200 281594 688000
rect 286322 687200 286378 688000
rect 291014 687200 291070 688000
rect 295706 687200 295762 688000
rect 300490 687200 300546 688000
rect 305182 687200 305238 688000
rect 309966 687200 310022 688000
rect 314658 687200 314714 688000
rect 319442 687200 319498 688000
rect 324134 687200 324190 688000
rect 328918 687200 328974 688000
rect 333610 687200 333666 688000
rect 338302 687200 338358 688000
rect 343086 687200 343142 688000
rect 347778 687200 347834 688000
rect 352562 687200 352618 688000
rect 357254 687200 357310 688000
rect 362038 687200 362094 688000
rect 366730 687200 366786 688000
rect 371514 687200 371570 688000
rect 376206 687200 376262 688000
rect 380990 687200 381046 688000
rect 385682 687200 385738 688000
rect 390374 687200 390430 688000
rect 395158 687200 395214 688000
rect 399850 687200 399906 688000
rect 404634 687200 404690 688000
rect 409326 687200 409382 688000
rect 414110 687200 414166 688000
rect 418802 687200 418858 688000
rect 423586 687200 423642 688000
rect 428278 687200 428334 688000
rect 432970 687200 433026 688000
rect 437754 687200 437810 688000
rect 442446 687200 442502 688000
rect 447230 687200 447286 688000
rect 451922 687200 451978 688000
rect 456706 687200 456762 688000
rect 461398 687200 461454 688000
rect 466182 687200 466238 688000
rect 470874 687200 470930 688000
rect 475658 687200 475714 688000
rect 480350 687200 480406 688000
rect 485042 687200 485098 688000
rect 489826 687200 489882 688000
rect 494518 687200 494574 688000
rect 499302 687200 499358 688000
rect 503994 687200 504050 688000
rect 508778 687200 508834 688000
rect 513470 687200 513526 688000
rect 518254 687200 518310 688000
rect 522946 687200 523002 688000
rect 527638 687200 527694 688000
rect 532422 687200 532478 688000
rect 537114 687200 537170 688000
rect 541898 687200 541954 688000
rect 546590 687200 546646 688000
rect 551374 687200 551430 688000
rect 556066 687200 556122 688000
rect 560850 687200 560906 688000
rect 565542 687200 565598 688000
rect 570 0 626 800
rect 1674 0 1730 800
rect 2778 0 2834 800
rect 3974 0 4030 800
rect 5078 0 5134 800
rect 6274 0 6330 800
rect 7378 0 7434 800
rect 8574 0 8630 800
rect 9678 0 9734 800
rect 10874 0 10930 800
rect 11978 0 12034 800
rect 13082 0 13138 800
rect 14278 0 14334 800
rect 15382 0 15438 800
rect 16578 0 16634 800
rect 17682 0 17738 800
rect 18878 0 18934 800
rect 19982 0 20038 800
rect 21178 0 21234 800
rect 22282 0 22338 800
rect 23386 0 23442 800
rect 24582 0 24638 800
rect 25686 0 25742 800
rect 26882 0 26938 800
rect 27986 0 28042 800
rect 29182 0 29238 800
rect 30286 0 30342 800
rect 31482 0 31538 800
rect 32586 0 32642 800
rect 33690 0 33746 800
rect 34886 0 34942 800
rect 35990 0 36046 800
rect 37186 0 37242 800
rect 38290 0 38346 800
rect 39486 0 39542 800
rect 40590 0 40646 800
rect 41786 0 41842 800
rect 42890 0 42946 800
rect 44086 0 44142 800
rect 45190 0 45246 800
rect 46294 0 46350 800
rect 47490 0 47546 800
rect 48594 0 48650 800
rect 49790 0 49846 800
rect 50894 0 50950 800
rect 52090 0 52146 800
rect 53194 0 53250 800
rect 54390 0 54446 800
rect 55494 0 55550 800
rect 56598 0 56654 800
rect 57794 0 57850 800
rect 58898 0 58954 800
rect 60094 0 60150 800
rect 61198 0 61254 800
rect 62394 0 62450 800
rect 63498 0 63554 800
rect 64694 0 64750 800
rect 65798 0 65854 800
rect 66902 0 66958 800
rect 68098 0 68154 800
rect 69202 0 69258 800
rect 70398 0 70454 800
rect 71502 0 71558 800
rect 72698 0 72754 800
rect 73802 0 73858 800
rect 74998 0 75054 800
rect 76102 0 76158 800
rect 77206 0 77262 800
rect 78402 0 78458 800
rect 79506 0 79562 800
rect 80702 0 80758 800
rect 81806 0 81862 800
rect 83002 0 83058 800
rect 84106 0 84162 800
rect 85302 0 85358 800
rect 86406 0 86462 800
rect 87602 0 87658 800
rect 88706 0 88762 800
rect 89810 0 89866 800
rect 91006 0 91062 800
rect 92110 0 92166 800
rect 93306 0 93362 800
rect 94410 0 94466 800
rect 95606 0 95662 800
rect 96710 0 96766 800
rect 97906 0 97962 800
rect 99010 0 99066 800
rect 100114 0 100170 800
rect 101310 0 101366 800
rect 102414 0 102470 800
rect 103610 0 103666 800
rect 104714 0 104770 800
rect 105910 0 105966 800
rect 107014 0 107070 800
rect 108210 0 108266 800
rect 109314 0 109370 800
rect 110418 0 110474 800
rect 111614 0 111670 800
rect 112718 0 112774 800
rect 113914 0 113970 800
rect 115018 0 115074 800
rect 116214 0 116270 800
rect 117318 0 117374 800
rect 118514 0 118570 800
rect 119618 0 119674 800
rect 120722 0 120778 800
rect 121918 0 121974 800
rect 123022 0 123078 800
rect 124218 0 124274 800
rect 125322 0 125378 800
rect 126518 0 126574 800
rect 127622 0 127678 800
rect 128818 0 128874 800
rect 129922 0 129978 800
rect 131118 0 131174 800
rect 132222 0 132278 800
rect 133326 0 133382 800
rect 134522 0 134578 800
rect 135626 0 135682 800
rect 136822 0 136878 800
rect 137926 0 137982 800
rect 139122 0 139178 800
rect 140226 0 140282 800
rect 141422 0 141478 800
rect 142526 0 142582 800
rect 143630 0 143686 800
rect 144826 0 144882 800
rect 145930 0 145986 800
rect 147126 0 147182 800
rect 148230 0 148286 800
rect 149426 0 149482 800
rect 150530 0 150586 800
rect 151726 0 151782 800
rect 152830 0 152886 800
rect 153934 0 153990 800
rect 155130 0 155186 800
rect 156234 0 156290 800
rect 157430 0 157486 800
rect 158534 0 158590 800
rect 159730 0 159786 800
rect 160834 0 160890 800
rect 162030 0 162086 800
rect 163134 0 163190 800
rect 164330 0 164386 800
rect 165434 0 165490 800
rect 166538 0 166594 800
rect 167734 0 167790 800
rect 168838 0 168894 800
rect 170034 0 170090 800
rect 171138 0 171194 800
rect 172334 0 172390 800
rect 173438 0 173494 800
rect 174634 0 174690 800
rect 175738 0 175794 800
rect 176842 0 176898 800
rect 178038 0 178094 800
rect 179142 0 179198 800
rect 180338 0 180394 800
rect 181442 0 181498 800
rect 182638 0 182694 800
rect 183742 0 183798 800
rect 184938 0 184994 800
rect 186042 0 186098 800
rect 187146 0 187202 800
rect 188342 0 188398 800
rect 189446 0 189502 800
rect 190642 0 190698 800
rect 191746 0 191802 800
rect 192942 0 192998 800
rect 194046 0 194102 800
rect 195242 0 195298 800
rect 196346 0 196402 800
rect 197450 0 197506 800
rect 198646 0 198702 800
rect 199750 0 199806 800
rect 200946 0 201002 800
rect 202050 0 202106 800
rect 203246 0 203302 800
rect 204350 0 204406 800
rect 205546 0 205602 800
rect 206650 0 206706 800
rect 207846 0 207902 800
rect 208950 0 209006 800
rect 210054 0 210110 800
rect 211250 0 211306 800
rect 212354 0 212410 800
rect 213550 0 213606 800
rect 214654 0 214710 800
rect 215850 0 215906 800
rect 216954 0 217010 800
rect 218150 0 218206 800
rect 219254 0 219310 800
rect 220358 0 220414 800
rect 221554 0 221610 800
rect 222658 0 222714 800
rect 223854 0 223910 800
rect 224958 0 225014 800
rect 226154 0 226210 800
rect 227258 0 227314 800
rect 228454 0 228510 800
rect 229558 0 229614 800
rect 230662 0 230718 800
rect 231858 0 231914 800
rect 232962 0 233018 800
rect 234158 0 234214 800
rect 235262 0 235318 800
rect 236458 0 236514 800
rect 237562 0 237618 800
rect 238758 0 238814 800
rect 239862 0 239918 800
rect 240966 0 241022 800
rect 242162 0 242218 800
rect 243266 0 243322 800
rect 244462 0 244518 800
rect 245566 0 245622 800
rect 246762 0 246818 800
rect 247866 0 247922 800
rect 249062 0 249118 800
rect 250166 0 250222 800
rect 251362 0 251418 800
rect 252466 0 252522 800
rect 253570 0 253626 800
rect 254766 0 254822 800
rect 255870 0 255926 800
rect 257066 0 257122 800
rect 258170 0 258226 800
rect 259366 0 259422 800
rect 260470 0 260526 800
rect 261666 0 261722 800
rect 262770 0 262826 800
rect 263874 0 263930 800
rect 265070 0 265126 800
rect 266174 0 266230 800
rect 267370 0 267426 800
rect 268474 0 268530 800
rect 269670 0 269726 800
rect 270774 0 270830 800
rect 271970 0 272026 800
rect 273074 0 273130 800
rect 274178 0 274234 800
rect 275374 0 275430 800
rect 276478 0 276534 800
rect 277674 0 277730 800
rect 278778 0 278834 800
rect 279974 0 280030 800
rect 281078 0 281134 800
rect 282274 0 282330 800
rect 283378 0 283434 800
rect 284574 0 284630 800
rect 285678 0 285734 800
rect 286782 0 286838 800
rect 287978 0 288034 800
rect 289082 0 289138 800
rect 290278 0 290334 800
rect 291382 0 291438 800
rect 292578 0 292634 800
rect 293682 0 293738 800
rect 294878 0 294934 800
rect 295982 0 296038 800
rect 297086 0 297142 800
rect 298282 0 298338 800
rect 299386 0 299442 800
rect 300582 0 300638 800
rect 301686 0 301742 800
rect 302882 0 302938 800
rect 303986 0 304042 800
rect 305182 0 305238 800
rect 306286 0 306342 800
rect 307390 0 307446 800
rect 308586 0 308642 800
rect 309690 0 309746 800
rect 310886 0 310942 800
rect 311990 0 312046 800
rect 313186 0 313242 800
rect 314290 0 314346 800
rect 315486 0 315542 800
rect 316590 0 316646 800
rect 317694 0 317750 800
rect 318890 0 318946 800
rect 319994 0 320050 800
rect 321190 0 321246 800
rect 322294 0 322350 800
rect 323490 0 323546 800
rect 324594 0 324650 800
rect 325790 0 325846 800
rect 326894 0 326950 800
rect 328090 0 328146 800
rect 329194 0 329250 800
rect 330298 0 330354 800
rect 331494 0 331550 800
rect 332598 0 332654 800
rect 333794 0 333850 800
rect 334898 0 334954 800
rect 336094 0 336150 800
rect 337198 0 337254 800
rect 338394 0 338450 800
rect 339498 0 339554 800
rect 340602 0 340658 800
rect 341798 0 341854 800
rect 342902 0 342958 800
rect 344098 0 344154 800
rect 345202 0 345258 800
rect 346398 0 346454 800
rect 347502 0 347558 800
rect 348698 0 348754 800
rect 349802 0 349858 800
rect 350906 0 350962 800
rect 352102 0 352158 800
rect 353206 0 353262 800
rect 354402 0 354458 800
rect 355506 0 355562 800
rect 356702 0 356758 800
rect 357806 0 357862 800
rect 359002 0 359058 800
rect 360106 0 360162 800
rect 361210 0 361266 800
rect 362406 0 362462 800
rect 363510 0 363566 800
rect 364706 0 364762 800
rect 365810 0 365866 800
rect 367006 0 367062 800
rect 368110 0 368166 800
rect 369306 0 369362 800
rect 370410 0 370466 800
rect 371606 0 371662 800
rect 372710 0 372766 800
rect 373814 0 373870 800
rect 375010 0 375066 800
rect 376114 0 376170 800
rect 377310 0 377366 800
rect 378414 0 378470 800
rect 379610 0 379666 800
rect 380714 0 380770 800
rect 381910 0 381966 800
rect 383014 0 383070 800
rect 384118 0 384174 800
rect 385314 0 385370 800
rect 386418 0 386474 800
rect 387614 0 387670 800
rect 388718 0 388774 800
rect 389914 0 389970 800
rect 391018 0 391074 800
rect 392214 0 392270 800
rect 393318 0 393374 800
rect 394422 0 394478 800
rect 395618 0 395674 800
rect 396722 0 396778 800
rect 397918 0 397974 800
rect 399022 0 399078 800
rect 400218 0 400274 800
rect 401322 0 401378 800
rect 402518 0 402574 800
rect 403622 0 403678 800
rect 404726 0 404782 800
rect 405922 0 405978 800
rect 407026 0 407082 800
rect 408222 0 408278 800
rect 409326 0 409382 800
rect 410522 0 410578 800
rect 411626 0 411682 800
rect 412822 0 412878 800
rect 413926 0 413982 800
rect 415122 0 415178 800
rect 416226 0 416282 800
rect 417330 0 417386 800
rect 418526 0 418582 800
rect 419630 0 419686 800
rect 420826 0 420882 800
rect 421930 0 421986 800
rect 423126 0 423182 800
rect 424230 0 424286 800
rect 425426 0 425482 800
rect 426530 0 426586 800
rect 427634 0 427690 800
rect 428830 0 428886 800
rect 429934 0 429990 800
rect 431130 0 431186 800
rect 432234 0 432290 800
rect 433430 0 433486 800
rect 434534 0 434590 800
rect 435730 0 435786 800
rect 436834 0 436890 800
rect 437938 0 437994 800
rect 439134 0 439190 800
rect 440238 0 440294 800
rect 441434 0 441490 800
rect 442538 0 442594 800
rect 443734 0 443790 800
rect 444838 0 444894 800
rect 446034 0 446090 800
rect 447138 0 447194 800
rect 448334 0 448390 800
rect 449438 0 449494 800
rect 450542 0 450598 800
rect 451738 0 451794 800
rect 452842 0 452898 800
rect 454038 0 454094 800
rect 455142 0 455198 800
rect 456338 0 456394 800
rect 457442 0 457498 800
rect 458638 0 458694 800
rect 459742 0 459798 800
rect 460846 0 460902 800
rect 462042 0 462098 800
rect 463146 0 463202 800
rect 464342 0 464398 800
rect 465446 0 465502 800
rect 466642 0 466698 800
rect 467746 0 467802 800
rect 468942 0 468998 800
rect 470046 0 470102 800
rect 471150 0 471206 800
rect 472346 0 472402 800
rect 473450 0 473506 800
rect 474646 0 474702 800
rect 475750 0 475806 800
rect 476946 0 477002 800
rect 478050 0 478106 800
rect 479246 0 479302 800
rect 480350 0 480406 800
rect 481454 0 481510 800
rect 482650 0 482706 800
rect 483754 0 483810 800
rect 484950 0 485006 800
rect 486054 0 486110 800
rect 487250 0 487306 800
rect 488354 0 488410 800
rect 489550 0 489606 800
rect 490654 0 490710 800
rect 491850 0 491906 800
rect 492954 0 493010 800
rect 494058 0 494114 800
rect 495254 0 495310 800
rect 496358 0 496414 800
rect 497554 0 497610 800
rect 498658 0 498714 800
rect 499854 0 499910 800
rect 500958 0 501014 800
rect 502154 0 502210 800
rect 503258 0 503314 800
rect 504362 0 504418 800
rect 505558 0 505614 800
rect 506662 0 506718 800
rect 507858 0 507914 800
rect 508962 0 509018 800
rect 510158 0 510214 800
rect 511262 0 511318 800
rect 512458 0 512514 800
rect 513562 0 513618 800
rect 514666 0 514722 800
rect 515862 0 515918 800
rect 516966 0 517022 800
rect 518162 0 518218 800
rect 519266 0 519322 800
rect 520462 0 520518 800
rect 521566 0 521622 800
rect 522762 0 522818 800
rect 523866 0 523922 800
rect 524970 0 525026 800
rect 526166 0 526222 800
rect 527270 0 527326 800
rect 528466 0 528522 800
rect 529570 0 529626 800
rect 530766 0 530822 800
rect 531870 0 531926 800
rect 533066 0 533122 800
rect 534170 0 534226 800
rect 535366 0 535422 800
rect 536470 0 536526 800
rect 537574 0 537630 800
rect 538770 0 538826 800
rect 539874 0 539930 800
rect 541070 0 541126 800
rect 542174 0 542230 800
rect 543370 0 543426 800
rect 544474 0 544530 800
rect 545670 0 545726 800
rect 546774 0 546830 800
rect 547878 0 547934 800
rect 549074 0 549130 800
rect 550178 0 550234 800
rect 551374 0 551430 800
rect 552478 0 552534 800
rect 553674 0 553730 800
rect 554778 0 554834 800
rect 555974 0 556030 800
rect 557078 0 557134 800
rect 558182 0 558238 800
rect 559378 0 559434 800
rect 560482 0 560538 800
rect 561678 0 561734 800
rect 562782 0 562838 800
rect 563978 0 564034 800
rect 565082 0 565138 800
rect 566278 0 566334 800
rect 567382 0 567438 800
<< obsm2 >>
rect 20 687144 2262 687200
rect 2430 687144 6954 687200
rect 7122 687144 11646 687200
rect 11814 687144 16430 687200
rect 16598 687144 21122 687200
rect 21290 687144 25906 687200
rect 26074 687144 30598 687200
rect 30766 687144 35382 687200
rect 35550 687144 40074 687200
rect 40242 687144 44858 687200
rect 45026 687144 49550 687200
rect 49718 687144 54242 687200
rect 54410 687144 59026 687200
rect 59194 687144 63718 687200
rect 63886 687144 68502 687200
rect 68670 687144 73194 687200
rect 73362 687144 77978 687200
rect 78146 687144 82670 687200
rect 82838 687144 87454 687200
rect 87622 687144 92146 687200
rect 92314 687144 96930 687200
rect 97098 687144 101622 687200
rect 101790 687144 106314 687200
rect 106482 687144 111098 687200
rect 111266 687144 115790 687200
rect 115958 687144 120574 687200
rect 120742 687144 125266 687200
rect 125434 687144 130050 687200
rect 130218 687144 134742 687200
rect 134910 687144 139526 687200
rect 139694 687144 144218 687200
rect 144386 687144 148910 687200
rect 149078 687144 153694 687200
rect 153862 687144 158386 687200
rect 158554 687144 163170 687200
rect 163338 687144 167862 687200
rect 168030 687144 172646 687200
rect 172814 687144 177338 687200
rect 177506 687144 182122 687200
rect 182290 687144 186814 687200
rect 186982 687144 191598 687200
rect 191766 687144 196290 687200
rect 196458 687144 200982 687200
rect 201150 687144 205766 687200
rect 205934 687144 210458 687200
rect 210626 687144 215242 687200
rect 215410 687144 219934 687200
rect 220102 687144 224718 687200
rect 224886 687144 229410 687200
rect 229578 687144 234194 687200
rect 234362 687144 238886 687200
rect 239054 687144 243578 687200
rect 243746 687144 248362 687200
rect 248530 687144 253054 687200
rect 253222 687144 257838 687200
rect 258006 687144 262530 687200
rect 262698 687144 267314 687200
rect 267482 687144 272006 687200
rect 272174 687144 276790 687200
rect 276958 687144 281482 687200
rect 281650 687144 286266 687200
rect 286434 687144 290958 687200
rect 291126 687144 295650 687200
rect 295818 687144 300434 687200
rect 300602 687144 305126 687200
rect 305294 687144 309910 687200
rect 310078 687144 314602 687200
rect 314770 687144 319386 687200
rect 319554 687144 324078 687200
rect 324246 687144 328862 687200
rect 329030 687144 333554 687200
rect 333722 687144 338246 687200
rect 338414 687144 343030 687200
rect 343198 687144 347722 687200
rect 347890 687144 352506 687200
rect 352674 687144 357198 687200
rect 357366 687144 361982 687200
rect 362150 687144 366674 687200
rect 366842 687144 371458 687200
rect 371626 687144 376150 687200
rect 376318 687144 380934 687200
rect 381102 687144 385626 687200
rect 385794 687144 390318 687200
rect 390486 687144 395102 687200
rect 395270 687144 399794 687200
rect 399962 687144 404578 687200
rect 404746 687144 409270 687200
rect 409438 687144 414054 687200
rect 414222 687144 418746 687200
rect 418914 687144 423530 687200
rect 423698 687144 428222 687200
rect 428390 687144 432914 687200
rect 433082 687144 437698 687200
rect 437866 687144 442390 687200
rect 442558 687144 447174 687200
rect 447342 687144 451866 687200
rect 452034 687144 456650 687200
rect 456818 687144 461342 687200
rect 461510 687144 466126 687200
rect 466294 687144 470818 687200
rect 470986 687144 475602 687200
rect 475770 687144 480294 687200
rect 480462 687144 484986 687200
rect 485154 687144 489770 687200
rect 489938 687144 494462 687200
rect 494630 687144 499246 687200
rect 499414 687144 503938 687200
rect 504106 687144 508722 687200
rect 508890 687144 513414 687200
rect 513582 687144 518198 687200
rect 518366 687144 522890 687200
rect 523058 687144 527582 687200
rect 527750 687144 532366 687200
rect 532534 687144 537058 687200
rect 537226 687144 541842 687200
rect 542010 687144 546534 687200
rect 546702 687144 551318 687200
rect 551486 687144 556010 687200
rect 556178 687144 560794 687200
rect 560962 687144 561734 687200
rect 20 856 561734 687144
rect 20 800 514 856
rect 682 800 1618 856
rect 1786 800 2722 856
rect 2890 800 3918 856
rect 4086 800 5022 856
rect 5190 800 6218 856
rect 6386 800 7322 856
rect 7490 800 8518 856
rect 8686 800 9622 856
rect 9790 800 10818 856
rect 10986 800 11922 856
rect 12090 800 13026 856
rect 13194 800 14222 856
rect 14390 800 15326 856
rect 15494 800 16522 856
rect 16690 800 17626 856
rect 17794 800 18822 856
rect 18990 800 19926 856
rect 20094 800 21122 856
rect 21290 800 22226 856
rect 22394 800 23330 856
rect 23498 800 24526 856
rect 24694 800 25630 856
rect 25798 800 26826 856
rect 26994 800 27930 856
rect 28098 800 29126 856
rect 29294 800 30230 856
rect 30398 800 31426 856
rect 31594 800 32530 856
rect 32698 800 33634 856
rect 33802 800 34830 856
rect 34998 800 35934 856
rect 36102 800 37130 856
rect 37298 800 38234 856
rect 38402 800 39430 856
rect 39598 800 40534 856
rect 40702 800 41730 856
rect 41898 800 42834 856
rect 43002 800 44030 856
rect 44198 800 45134 856
rect 45302 800 46238 856
rect 46406 800 47434 856
rect 47602 800 48538 856
rect 48706 800 49734 856
rect 49902 800 50838 856
rect 51006 800 52034 856
rect 52202 800 53138 856
rect 53306 800 54334 856
rect 54502 800 55438 856
rect 55606 800 56542 856
rect 56710 800 57738 856
rect 57906 800 58842 856
rect 59010 800 60038 856
rect 60206 800 61142 856
rect 61310 800 62338 856
rect 62506 800 63442 856
rect 63610 800 64638 856
rect 64806 800 65742 856
rect 65910 800 66846 856
rect 67014 800 68042 856
rect 68210 800 69146 856
rect 69314 800 70342 856
rect 70510 800 71446 856
rect 71614 800 72642 856
rect 72810 800 73746 856
rect 73914 800 74942 856
rect 75110 800 76046 856
rect 76214 800 77150 856
rect 77318 800 78346 856
rect 78514 800 79450 856
rect 79618 800 80646 856
rect 80814 800 81750 856
rect 81918 800 82946 856
rect 83114 800 84050 856
rect 84218 800 85246 856
rect 85414 800 86350 856
rect 86518 800 87546 856
rect 87714 800 88650 856
rect 88818 800 89754 856
rect 89922 800 90950 856
rect 91118 800 92054 856
rect 92222 800 93250 856
rect 93418 800 94354 856
rect 94522 800 95550 856
rect 95718 800 96654 856
rect 96822 800 97850 856
rect 98018 800 98954 856
rect 99122 800 100058 856
rect 100226 800 101254 856
rect 101422 800 102358 856
rect 102526 800 103554 856
rect 103722 800 104658 856
rect 104826 800 105854 856
rect 106022 800 106958 856
rect 107126 800 108154 856
rect 108322 800 109258 856
rect 109426 800 110362 856
rect 110530 800 111558 856
rect 111726 800 112662 856
rect 112830 800 113858 856
rect 114026 800 114962 856
rect 115130 800 116158 856
rect 116326 800 117262 856
rect 117430 800 118458 856
rect 118626 800 119562 856
rect 119730 800 120666 856
rect 120834 800 121862 856
rect 122030 800 122966 856
rect 123134 800 124162 856
rect 124330 800 125266 856
rect 125434 800 126462 856
rect 126630 800 127566 856
rect 127734 800 128762 856
rect 128930 800 129866 856
rect 130034 800 131062 856
rect 131230 800 132166 856
rect 132334 800 133270 856
rect 133438 800 134466 856
rect 134634 800 135570 856
rect 135738 800 136766 856
rect 136934 800 137870 856
rect 138038 800 139066 856
rect 139234 800 140170 856
rect 140338 800 141366 856
rect 141534 800 142470 856
rect 142638 800 143574 856
rect 143742 800 144770 856
rect 144938 800 145874 856
rect 146042 800 147070 856
rect 147238 800 148174 856
rect 148342 800 149370 856
rect 149538 800 150474 856
rect 150642 800 151670 856
rect 151838 800 152774 856
rect 152942 800 153878 856
rect 154046 800 155074 856
rect 155242 800 156178 856
rect 156346 800 157374 856
rect 157542 800 158478 856
rect 158646 800 159674 856
rect 159842 800 160778 856
rect 160946 800 161974 856
rect 162142 800 163078 856
rect 163246 800 164274 856
rect 164442 800 165378 856
rect 165546 800 166482 856
rect 166650 800 167678 856
rect 167846 800 168782 856
rect 168950 800 169978 856
rect 170146 800 171082 856
rect 171250 800 172278 856
rect 172446 800 173382 856
rect 173550 800 174578 856
rect 174746 800 175682 856
rect 175850 800 176786 856
rect 176954 800 177982 856
rect 178150 800 179086 856
rect 179254 800 180282 856
rect 180450 800 181386 856
rect 181554 800 182582 856
rect 182750 800 183686 856
rect 183854 800 184882 856
rect 185050 800 185986 856
rect 186154 800 187090 856
rect 187258 800 188286 856
rect 188454 800 189390 856
rect 189558 800 190586 856
rect 190754 800 191690 856
rect 191858 800 192886 856
rect 193054 800 193990 856
rect 194158 800 195186 856
rect 195354 800 196290 856
rect 196458 800 197394 856
rect 197562 800 198590 856
rect 198758 800 199694 856
rect 199862 800 200890 856
rect 201058 800 201994 856
rect 202162 800 203190 856
rect 203358 800 204294 856
rect 204462 800 205490 856
rect 205658 800 206594 856
rect 206762 800 207790 856
rect 207958 800 208894 856
rect 209062 800 209998 856
rect 210166 800 211194 856
rect 211362 800 212298 856
rect 212466 800 213494 856
rect 213662 800 214598 856
rect 214766 800 215794 856
rect 215962 800 216898 856
rect 217066 800 218094 856
rect 218262 800 219198 856
rect 219366 800 220302 856
rect 220470 800 221498 856
rect 221666 800 222602 856
rect 222770 800 223798 856
rect 223966 800 224902 856
rect 225070 800 226098 856
rect 226266 800 227202 856
rect 227370 800 228398 856
rect 228566 800 229502 856
rect 229670 800 230606 856
rect 230774 800 231802 856
rect 231970 800 232906 856
rect 233074 800 234102 856
rect 234270 800 235206 856
rect 235374 800 236402 856
rect 236570 800 237506 856
rect 237674 800 238702 856
rect 238870 800 239806 856
rect 239974 800 240910 856
rect 241078 800 242106 856
rect 242274 800 243210 856
rect 243378 800 244406 856
rect 244574 800 245510 856
rect 245678 800 246706 856
rect 246874 800 247810 856
rect 247978 800 249006 856
rect 249174 800 250110 856
rect 250278 800 251306 856
rect 251474 800 252410 856
rect 252578 800 253514 856
rect 253682 800 254710 856
rect 254878 800 255814 856
rect 255982 800 257010 856
rect 257178 800 258114 856
rect 258282 800 259310 856
rect 259478 800 260414 856
rect 260582 800 261610 856
rect 261778 800 262714 856
rect 262882 800 263818 856
rect 263986 800 265014 856
rect 265182 800 266118 856
rect 266286 800 267314 856
rect 267482 800 268418 856
rect 268586 800 269614 856
rect 269782 800 270718 856
rect 270886 800 271914 856
rect 272082 800 273018 856
rect 273186 800 274122 856
rect 274290 800 275318 856
rect 275486 800 276422 856
rect 276590 800 277618 856
rect 277786 800 278722 856
rect 278890 800 279918 856
rect 280086 800 281022 856
rect 281190 800 282218 856
rect 282386 800 283322 856
rect 283490 800 284518 856
rect 284686 800 285622 856
rect 285790 800 286726 856
rect 286894 800 287922 856
rect 288090 800 289026 856
rect 289194 800 290222 856
rect 290390 800 291326 856
rect 291494 800 292522 856
rect 292690 800 293626 856
rect 293794 800 294822 856
rect 294990 800 295926 856
rect 296094 800 297030 856
rect 297198 800 298226 856
rect 298394 800 299330 856
rect 299498 800 300526 856
rect 300694 800 301630 856
rect 301798 800 302826 856
rect 302994 800 303930 856
rect 304098 800 305126 856
rect 305294 800 306230 856
rect 306398 800 307334 856
rect 307502 800 308530 856
rect 308698 800 309634 856
rect 309802 800 310830 856
rect 310998 800 311934 856
rect 312102 800 313130 856
rect 313298 800 314234 856
rect 314402 800 315430 856
rect 315598 800 316534 856
rect 316702 800 317638 856
rect 317806 800 318834 856
rect 319002 800 319938 856
rect 320106 800 321134 856
rect 321302 800 322238 856
rect 322406 800 323434 856
rect 323602 800 324538 856
rect 324706 800 325734 856
rect 325902 800 326838 856
rect 327006 800 328034 856
rect 328202 800 329138 856
rect 329306 800 330242 856
rect 330410 800 331438 856
rect 331606 800 332542 856
rect 332710 800 333738 856
rect 333906 800 334842 856
rect 335010 800 336038 856
rect 336206 800 337142 856
rect 337310 800 338338 856
rect 338506 800 339442 856
rect 339610 800 340546 856
rect 340714 800 341742 856
rect 341910 800 342846 856
rect 343014 800 344042 856
rect 344210 800 345146 856
rect 345314 800 346342 856
rect 346510 800 347446 856
rect 347614 800 348642 856
rect 348810 800 349746 856
rect 349914 800 350850 856
rect 351018 800 352046 856
rect 352214 800 353150 856
rect 353318 800 354346 856
rect 354514 800 355450 856
rect 355618 800 356646 856
rect 356814 800 357750 856
rect 357918 800 358946 856
rect 359114 800 360050 856
rect 360218 800 361154 856
rect 361322 800 362350 856
rect 362518 800 363454 856
rect 363622 800 364650 856
rect 364818 800 365754 856
rect 365922 800 366950 856
rect 367118 800 368054 856
rect 368222 800 369250 856
rect 369418 800 370354 856
rect 370522 800 371550 856
rect 371718 800 372654 856
rect 372822 800 373758 856
rect 373926 800 374954 856
rect 375122 800 376058 856
rect 376226 800 377254 856
rect 377422 800 378358 856
rect 378526 800 379554 856
rect 379722 800 380658 856
rect 380826 800 381854 856
rect 382022 800 382958 856
rect 383126 800 384062 856
rect 384230 800 385258 856
rect 385426 800 386362 856
rect 386530 800 387558 856
rect 387726 800 388662 856
rect 388830 800 389858 856
rect 390026 800 390962 856
rect 391130 800 392158 856
rect 392326 800 393262 856
rect 393430 800 394366 856
rect 394534 800 395562 856
rect 395730 800 396666 856
rect 396834 800 397862 856
rect 398030 800 398966 856
rect 399134 800 400162 856
rect 400330 800 401266 856
rect 401434 800 402462 856
rect 402630 800 403566 856
rect 403734 800 404670 856
rect 404838 800 405866 856
rect 406034 800 406970 856
rect 407138 800 408166 856
rect 408334 800 409270 856
rect 409438 800 410466 856
rect 410634 800 411570 856
rect 411738 800 412766 856
rect 412934 800 413870 856
rect 414038 800 415066 856
rect 415234 800 416170 856
rect 416338 800 417274 856
rect 417442 800 418470 856
rect 418638 800 419574 856
rect 419742 800 420770 856
rect 420938 800 421874 856
rect 422042 800 423070 856
rect 423238 800 424174 856
rect 424342 800 425370 856
rect 425538 800 426474 856
rect 426642 800 427578 856
rect 427746 800 428774 856
rect 428942 800 429878 856
rect 430046 800 431074 856
rect 431242 800 432178 856
rect 432346 800 433374 856
rect 433542 800 434478 856
rect 434646 800 435674 856
rect 435842 800 436778 856
rect 436946 800 437882 856
rect 438050 800 439078 856
rect 439246 800 440182 856
rect 440350 800 441378 856
rect 441546 800 442482 856
rect 442650 800 443678 856
rect 443846 800 444782 856
rect 444950 800 445978 856
rect 446146 800 447082 856
rect 447250 800 448278 856
rect 448446 800 449382 856
rect 449550 800 450486 856
rect 450654 800 451682 856
rect 451850 800 452786 856
rect 452954 800 453982 856
rect 454150 800 455086 856
rect 455254 800 456282 856
rect 456450 800 457386 856
rect 457554 800 458582 856
rect 458750 800 459686 856
rect 459854 800 460790 856
rect 460958 800 461986 856
rect 462154 800 463090 856
rect 463258 800 464286 856
rect 464454 800 465390 856
rect 465558 800 466586 856
rect 466754 800 467690 856
rect 467858 800 468886 856
rect 469054 800 469990 856
rect 470158 800 471094 856
rect 471262 800 472290 856
rect 472458 800 473394 856
rect 473562 800 474590 856
rect 474758 800 475694 856
rect 475862 800 476890 856
rect 477058 800 477994 856
rect 478162 800 479190 856
rect 479358 800 480294 856
rect 480462 800 481398 856
rect 481566 800 482594 856
rect 482762 800 483698 856
rect 483866 800 484894 856
rect 485062 800 485998 856
rect 486166 800 487194 856
rect 487362 800 488298 856
rect 488466 800 489494 856
rect 489662 800 490598 856
rect 490766 800 491794 856
rect 491962 800 492898 856
rect 493066 800 494002 856
rect 494170 800 495198 856
rect 495366 800 496302 856
rect 496470 800 497498 856
rect 497666 800 498602 856
rect 498770 800 499798 856
rect 499966 800 500902 856
rect 501070 800 502098 856
rect 502266 800 503202 856
rect 503370 800 504306 856
rect 504474 800 505502 856
rect 505670 800 506606 856
rect 506774 800 507802 856
rect 507970 800 508906 856
rect 509074 800 510102 856
rect 510270 800 511206 856
rect 511374 800 512402 856
rect 512570 800 513506 856
rect 513674 800 514610 856
rect 514778 800 515806 856
rect 515974 800 516910 856
rect 517078 800 518106 856
rect 518274 800 519210 856
rect 519378 800 520406 856
rect 520574 800 521510 856
rect 521678 800 522706 856
rect 522874 800 523810 856
rect 523978 800 524914 856
rect 525082 800 526110 856
rect 526278 800 527214 856
rect 527382 800 528410 856
rect 528578 800 529514 856
rect 529682 800 530710 856
rect 530878 800 531814 856
rect 531982 800 533010 856
rect 533178 800 534114 856
rect 534282 800 535310 856
rect 535478 800 536414 856
rect 536582 800 537518 856
rect 537686 800 538714 856
rect 538882 800 539818 856
rect 539986 800 541014 856
rect 541182 800 542118 856
rect 542286 800 543314 856
rect 543482 800 544418 856
rect 544586 800 545614 856
rect 545782 800 546718 856
rect 546886 800 547822 856
rect 547990 800 549018 856
rect 549186 800 550122 856
rect 550290 800 551318 856
rect 551486 800 552422 856
rect 552590 800 553618 856
rect 553786 800 554722 856
rect 554890 800 555918 856
rect 556086 800 557022 856
rect 557190 800 558126 856
rect 558294 800 559322 856
rect 559490 800 560426 856
rect 560594 800 561622 856
<< metal3 >>
rect 0 649680 800 649800
rect 0 573248 800 573368
rect 0 496816 800 496936
rect 0 420384 800 420504
rect 0 343952 800 344072
rect 0 267520 800 267640
rect 0 191088 800 191208
rect 0 114656 800 114776
rect 0 38224 800 38344
rect 567200 656616 568000 656736
rect 567200 594056 568000 594176
rect 567200 531496 568000 531616
rect 567200 468936 568000 469056
rect 567200 406376 568000 406496
rect 567200 343816 568000 343936
rect 567200 281256 568000 281376
rect 567200 218696 568000 218816
rect 567200 156136 568000 156256
rect 567200 93576 568000 93696
rect 567200 31152 568000 31272
<< obsm3 >>
rect 2405 2143 561739 685473
<< metal4 >>
rect 4208 2128 4528 685488
rect 19568 2128 19888 685488
rect 34928 2128 35248 685488
rect 50288 2128 50608 685488
rect 65648 2128 65968 685488
rect 81008 2128 81328 685488
rect 96368 2128 96688 685488
rect 111728 2128 112048 685488
rect 127088 2128 127408 685488
rect 142448 2128 142768 685488
rect 157808 2128 158128 685488
rect 173168 2128 173488 685488
rect 188528 2128 188848 685488
rect 203888 2128 204208 685488
rect 219248 2128 219568 685488
rect 234608 2128 234928 685488
rect 249968 2128 250288 685488
rect 265328 2128 265648 685488
rect 280688 2128 281008 685488
rect 296048 2128 296368 685488
rect 311408 2128 311728 685488
rect 326768 2128 327088 685488
rect 342128 2128 342448 685488
rect 357488 2128 357808 685488
rect 372848 2128 373168 685488
rect 388208 2128 388528 685488
rect 403568 2128 403888 685488
rect 418928 2128 419248 685488
rect 434288 2128 434608 685488
rect 449648 2128 449968 685488
rect 465008 2128 465328 685488
rect 480368 2128 480688 685488
rect 495728 2128 496048 685488
rect 511088 2128 511408 685488
rect 526448 2128 526768 685488
rect 541808 2128 542128 685488
rect 557168 2128 557488 685488
<< obsm4 >>
rect 3003 2483 4128 683637
rect 4608 2483 19488 683637
rect 19968 2483 34848 683637
rect 35328 2483 50208 683637
rect 50688 2483 65568 683637
rect 66048 2483 80928 683637
rect 81408 2483 96288 683637
rect 96768 2483 111648 683637
rect 112128 2483 127008 683637
rect 127488 2483 142368 683637
rect 142848 2483 157728 683637
rect 158208 2483 173088 683637
rect 173568 2483 188448 683637
rect 188928 2483 203808 683637
rect 204288 2483 219168 683637
rect 219648 2483 234528 683637
rect 235008 2483 249888 683637
rect 250368 2483 265248 683637
rect 265728 2483 280608 683637
rect 281088 2483 295968 683637
rect 296448 2483 311328 683637
rect 311808 2483 326688 683637
rect 327168 2483 342048 683637
rect 342528 2483 357408 683637
rect 357888 2483 372768 683637
rect 373248 2483 388128 683637
rect 388608 2483 403488 683637
rect 403968 2483 418848 683637
rect 419328 2483 434208 683637
rect 434688 2483 449568 683637
rect 450048 2483 464928 683637
rect 465408 2483 480288 683637
rect 480768 2483 495648 683637
rect 496128 2483 511008 683637
rect 511488 2483 526368 683637
rect 526848 2483 541728 683637
rect 542208 2483 549733 683637
<< labels >>
rlabel metal3 s 567200 31152 568000 31272 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 546590 687200 546646 688000 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 551374 687200 551430 688000 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal3 s 0 343952 800 344072 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal3 s 567200 281256 568000 281376 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 563978 0 564034 800 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal3 s 0 420384 800 420504 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal3 s 567200 343816 568000 343936 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s 567200 406376 568000 406496 6 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s 0 496816 800 496936 6 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s 567200 468936 568000 469056 6 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal2 s 541898 687200 541954 688000 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal2 s 556066 687200 556122 688000 6 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s 0 573248 800 573368 6 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal2 s 565082 0 565138 800 6 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal2 s 560850 687200 560906 688000 6 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal2 s 565542 687200 565598 688000 6 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s 0 649680 800 649800 6 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal2 s 566278 0 566334 800 6 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s 567200 531496 568000 531616 6 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal2 s 567382 0 567438 800 6 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 567200 594056 568000 594176 6 analog_io[29]
port 22 nsew signal bidirectional
rlabel metal3 s 0 38224 800 38344 6 analog_io[2]
port 23 nsew signal bidirectional
rlabel metal3 s 567200 656616 568000 656736 6 analog_io[30]
port 24 nsew signal bidirectional
rlabel metal3 s 567200 93576 568000 93696 6 analog_io[3]
port 25 nsew signal bidirectional
rlabel metal3 s 0 114656 800 114776 6 analog_io[4]
port 26 nsew signal bidirectional
rlabel metal3 s 0 191088 800 191208 6 analog_io[5]
port 27 nsew signal bidirectional
rlabel metal3 s 567200 156136 568000 156256 6 analog_io[6]
port 28 nsew signal bidirectional
rlabel metal3 s 0 267520 800 267640 6 analog_io[7]
port 29 nsew signal bidirectional
rlabel metal3 s 567200 218696 568000 218816 6 analog_io[8]
port 30 nsew signal bidirectional
rlabel metal2 s 562782 0 562838 800 6 analog_io[9]
port 31 nsew signal bidirectional
rlabel metal2 s 2318 687200 2374 688000 6 io_in[0]
port 32 nsew signal input
rlabel metal2 s 144274 687200 144330 688000 6 io_in[10]
port 33 nsew signal input
rlabel metal2 s 158442 687200 158498 688000 6 io_in[11]
port 34 nsew signal input
rlabel metal2 s 172702 687200 172758 688000 6 io_in[12]
port 35 nsew signal input
rlabel metal2 s 186870 687200 186926 688000 6 io_in[13]
port 36 nsew signal input
rlabel metal2 s 201038 687200 201094 688000 6 io_in[14]
port 37 nsew signal input
rlabel metal2 s 215298 687200 215354 688000 6 io_in[15]
port 38 nsew signal input
rlabel metal2 s 229466 687200 229522 688000 6 io_in[16]
port 39 nsew signal input
rlabel metal2 s 243634 687200 243690 688000 6 io_in[17]
port 40 nsew signal input
rlabel metal2 s 257894 687200 257950 688000 6 io_in[18]
port 41 nsew signal input
rlabel metal2 s 272062 687200 272118 688000 6 io_in[19]
port 42 nsew signal input
rlabel metal2 s 16486 687200 16542 688000 6 io_in[1]
port 43 nsew signal input
rlabel metal2 s 286322 687200 286378 688000 6 io_in[20]
port 44 nsew signal input
rlabel metal2 s 300490 687200 300546 688000 6 io_in[21]
port 45 nsew signal input
rlabel metal2 s 314658 687200 314714 688000 6 io_in[22]
port 46 nsew signal input
rlabel metal2 s 328918 687200 328974 688000 6 io_in[23]
port 47 nsew signal input
rlabel metal2 s 343086 687200 343142 688000 6 io_in[24]
port 48 nsew signal input
rlabel metal2 s 357254 687200 357310 688000 6 io_in[25]
port 49 nsew signal input
rlabel metal2 s 371514 687200 371570 688000 6 io_in[26]
port 50 nsew signal input
rlabel metal2 s 385682 687200 385738 688000 6 io_in[27]
port 51 nsew signal input
rlabel metal2 s 399850 687200 399906 688000 6 io_in[28]
port 52 nsew signal input
rlabel metal2 s 414110 687200 414166 688000 6 io_in[29]
port 53 nsew signal input
rlabel metal2 s 30654 687200 30710 688000 6 io_in[2]
port 54 nsew signal input
rlabel metal2 s 428278 687200 428334 688000 6 io_in[30]
port 55 nsew signal input
rlabel metal2 s 442446 687200 442502 688000 6 io_in[31]
port 56 nsew signal input
rlabel metal2 s 456706 687200 456762 688000 6 io_in[32]
port 57 nsew signal input
rlabel metal2 s 470874 687200 470930 688000 6 io_in[33]
port 58 nsew signal input
rlabel metal2 s 485042 687200 485098 688000 6 io_in[34]
port 59 nsew signal input
rlabel metal2 s 499302 687200 499358 688000 6 io_in[35]
port 60 nsew signal input
rlabel metal2 s 513470 687200 513526 688000 6 io_in[36]
port 61 nsew signal input
rlabel metal2 s 527638 687200 527694 688000 6 io_in[37]
port 62 nsew signal input
rlabel metal2 s 44914 687200 44970 688000 6 io_in[3]
port 63 nsew signal input
rlabel metal2 s 59082 687200 59138 688000 6 io_in[4]
port 64 nsew signal input
rlabel metal2 s 73250 687200 73306 688000 6 io_in[5]
port 65 nsew signal input
rlabel metal2 s 87510 687200 87566 688000 6 io_in[6]
port 66 nsew signal input
rlabel metal2 s 101678 687200 101734 688000 6 io_in[7]
port 67 nsew signal input
rlabel metal2 s 115846 687200 115902 688000 6 io_in[8]
port 68 nsew signal input
rlabel metal2 s 130106 687200 130162 688000 6 io_in[9]
port 69 nsew signal input
rlabel metal2 s 7010 687200 7066 688000 6 io_oeb[0]
port 70 nsew signal output
rlabel metal2 s 148966 687200 149022 688000 6 io_oeb[10]
port 71 nsew signal output
rlabel metal2 s 163226 687200 163282 688000 6 io_oeb[11]
port 72 nsew signal output
rlabel metal2 s 177394 687200 177450 688000 6 io_oeb[12]
port 73 nsew signal output
rlabel metal2 s 191654 687200 191710 688000 6 io_oeb[13]
port 74 nsew signal output
rlabel metal2 s 205822 687200 205878 688000 6 io_oeb[14]
port 75 nsew signal output
rlabel metal2 s 219990 687200 220046 688000 6 io_oeb[15]
port 76 nsew signal output
rlabel metal2 s 234250 687200 234306 688000 6 io_oeb[16]
port 77 nsew signal output
rlabel metal2 s 248418 687200 248474 688000 6 io_oeb[17]
port 78 nsew signal output
rlabel metal2 s 262586 687200 262642 688000 6 io_oeb[18]
port 79 nsew signal output
rlabel metal2 s 276846 687200 276902 688000 6 io_oeb[19]
port 80 nsew signal output
rlabel metal2 s 21178 687200 21234 688000 6 io_oeb[1]
port 81 nsew signal output
rlabel metal2 s 291014 687200 291070 688000 6 io_oeb[20]
port 82 nsew signal output
rlabel metal2 s 305182 687200 305238 688000 6 io_oeb[21]
port 83 nsew signal output
rlabel metal2 s 319442 687200 319498 688000 6 io_oeb[22]
port 84 nsew signal output
rlabel metal2 s 333610 687200 333666 688000 6 io_oeb[23]
port 85 nsew signal output
rlabel metal2 s 347778 687200 347834 688000 6 io_oeb[24]
port 86 nsew signal output
rlabel metal2 s 362038 687200 362094 688000 6 io_oeb[25]
port 87 nsew signal output
rlabel metal2 s 376206 687200 376262 688000 6 io_oeb[26]
port 88 nsew signal output
rlabel metal2 s 390374 687200 390430 688000 6 io_oeb[27]
port 89 nsew signal output
rlabel metal2 s 404634 687200 404690 688000 6 io_oeb[28]
port 90 nsew signal output
rlabel metal2 s 418802 687200 418858 688000 6 io_oeb[29]
port 91 nsew signal output
rlabel metal2 s 35438 687200 35494 688000 6 io_oeb[2]
port 92 nsew signal output
rlabel metal2 s 432970 687200 433026 688000 6 io_oeb[30]
port 93 nsew signal output
rlabel metal2 s 447230 687200 447286 688000 6 io_oeb[31]
port 94 nsew signal output
rlabel metal2 s 461398 687200 461454 688000 6 io_oeb[32]
port 95 nsew signal output
rlabel metal2 s 475658 687200 475714 688000 6 io_oeb[33]
port 96 nsew signal output
rlabel metal2 s 489826 687200 489882 688000 6 io_oeb[34]
port 97 nsew signal output
rlabel metal2 s 503994 687200 504050 688000 6 io_oeb[35]
port 98 nsew signal output
rlabel metal2 s 518254 687200 518310 688000 6 io_oeb[36]
port 99 nsew signal output
rlabel metal2 s 532422 687200 532478 688000 6 io_oeb[37]
port 100 nsew signal output
rlabel metal2 s 49606 687200 49662 688000 6 io_oeb[3]
port 101 nsew signal output
rlabel metal2 s 63774 687200 63830 688000 6 io_oeb[4]
port 102 nsew signal output
rlabel metal2 s 78034 687200 78090 688000 6 io_oeb[5]
port 103 nsew signal output
rlabel metal2 s 92202 687200 92258 688000 6 io_oeb[6]
port 104 nsew signal output
rlabel metal2 s 106370 687200 106426 688000 6 io_oeb[7]
port 105 nsew signal output
rlabel metal2 s 120630 687200 120686 688000 6 io_oeb[8]
port 106 nsew signal output
rlabel metal2 s 134798 687200 134854 688000 6 io_oeb[9]
port 107 nsew signal output
rlabel metal2 s 11702 687200 11758 688000 6 io_out[0]
port 108 nsew signal output
rlabel metal2 s 153750 687200 153806 688000 6 io_out[10]
port 109 nsew signal output
rlabel metal2 s 167918 687200 167974 688000 6 io_out[11]
port 110 nsew signal output
rlabel metal2 s 182178 687200 182234 688000 6 io_out[12]
port 111 nsew signal output
rlabel metal2 s 196346 687200 196402 688000 6 io_out[13]
port 112 nsew signal output
rlabel metal2 s 210514 687200 210570 688000 6 io_out[14]
port 113 nsew signal output
rlabel metal2 s 224774 687200 224830 688000 6 io_out[15]
port 114 nsew signal output
rlabel metal2 s 238942 687200 238998 688000 6 io_out[16]
port 115 nsew signal output
rlabel metal2 s 253110 687200 253166 688000 6 io_out[17]
port 116 nsew signal output
rlabel metal2 s 267370 687200 267426 688000 6 io_out[18]
port 117 nsew signal output
rlabel metal2 s 281538 687200 281594 688000 6 io_out[19]
port 118 nsew signal output
rlabel metal2 s 25962 687200 26018 688000 6 io_out[1]
port 119 nsew signal output
rlabel metal2 s 295706 687200 295762 688000 6 io_out[20]
port 120 nsew signal output
rlabel metal2 s 309966 687200 310022 688000 6 io_out[21]
port 121 nsew signal output
rlabel metal2 s 324134 687200 324190 688000 6 io_out[22]
port 122 nsew signal output
rlabel metal2 s 338302 687200 338358 688000 6 io_out[23]
port 123 nsew signal output
rlabel metal2 s 352562 687200 352618 688000 6 io_out[24]
port 124 nsew signal output
rlabel metal2 s 366730 687200 366786 688000 6 io_out[25]
port 125 nsew signal output
rlabel metal2 s 380990 687200 381046 688000 6 io_out[26]
port 126 nsew signal output
rlabel metal2 s 395158 687200 395214 688000 6 io_out[27]
port 127 nsew signal output
rlabel metal2 s 409326 687200 409382 688000 6 io_out[28]
port 128 nsew signal output
rlabel metal2 s 423586 687200 423642 688000 6 io_out[29]
port 129 nsew signal output
rlabel metal2 s 40130 687200 40186 688000 6 io_out[2]
port 130 nsew signal output
rlabel metal2 s 437754 687200 437810 688000 6 io_out[30]
port 131 nsew signal output
rlabel metal2 s 451922 687200 451978 688000 6 io_out[31]
port 132 nsew signal output
rlabel metal2 s 466182 687200 466238 688000 6 io_out[32]
port 133 nsew signal output
rlabel metal2 s 480350 687200 480406 688000 6 io_out[33]
port 134 nsew signal output
rlabel metal2 s 494518 687200 494574 688000 6 io_out[34]
port 135 nsew signal output
rlabel metal2 s 508778 687200 508834 688000 6 io_out[35]
port 136 nsew signal output
rlabel metal2 s 522946 687200 523002 688000 6 io_out[36]
port 137 nsew signal output
rlabel metal2 s 537114 687200 537170 688000 6 io_out[37]
port 138 nsew signal output
rlabel metal2 s 54298 687200 54354 688000 6 io_out[3]
port 139 nsew signal output
rlabel metal2 s 68558 687200 68614 688000 6 io_out[4]
port 140 nsew signal output
rlabel metal2 s 82726 687200 82782 688000 6 io_out[5]
port 141 nsew signal output
rlabel metal2 s 96986 687200 97042 688000 6 io_out[6]
port 142 nsew signal output
rlabel metal2 s 111154 687200 111210 688000 6 io_out[7]
port 143 nsew signal output
rlabel metal2 s 125322 687200 125378 688000 6 io_out[8]
port 144 nsew signal output
rlabel metal2 s 139582 687200 139638 688000 6 io_out[9]
port 145 nsew signal output
rlabel metal2 s 121918 0 121974 800 6 la_data_in[0]
port 146 nsew signal input
rlabel metal2 s 465446 0 465502 800 6 la_data_in[100]
port 147 nsew signal input
rlabel metal2 s 468942 0 468998 800 6 la_data_in[101]
port 148 nsew signal input
rlabel metal2 s 472346 0 472402 800 6 la_data_in[102]
port 149 nsew signal input
rlabel metal2 s 475750 0 475806 800 6 la_data_in[103]
port 150 nsew signal input
rlabel metal2 s 479246 0 479302 800 6 la_data_in[104]
port 151 nsew signal input
rlabel metal2 s 482650 0 482706 800 6 la_data_in[105]
port 152 nsew signal input
rlabel metal2 s 486054 0 486110 800 6 la_data_in[106]
port 153 nsew signal input
rlabel metal2 s 489550 0 489606 800 6 la_data_in[107]
port 154 nsew signal input
rlabel metal2 s 492954 0 493010 800 6 la_data_in[108]
port 155 nsew signal input
rlabel metal2 s 496358 0 496414 800 6 la_data_in[109]
port 156 nsew signal input
rlabel metal2 s 156234 0 156290 800 6 la_data_in[10]
port 157 nsew signal input
rlabel metal2 s 499854 0 499910 800 6 la_data_in[110]
port 158 nsew signal input
rlabel metal2 s 503258 0 503314 800 6 la_data_in[111]
port 159 nsew signal input
rlabel metal2 s 506662 0 506718 800 6 la_data_in[112]
port 160 nsew signal input
rlabel metal2 s 510158 0 510214 800 6 la_data_in[113]
port 161 nsew signal input
rlabel metal2 s 513562 0 513618 800 6 la_data_in[114]
port 162 nsew signal input
rlabel metal2 s 516966 0 517022 800 6 la_data_in[115]
port 163 nsew signal input
rlabel metal2 s 520462 0 520518 800 6 la_data_in[116]
port 164 nsew signal input
rlabel metal2 s 523866 0 523922 800 6 la_data_in[117]
port 165 nsew signal input
rlabel metal2 s 527270 0 527326 800 6 la_data_in[118]
port 166 nsew signal input
rlabel metal2 s 530766 0 530822 800 6 la_data_in[119]
port 167 nsew signal input
rlabel metal2 s 159730 0 159786 800 6 la_data_in[11]
port 168 nsew signal input
rlabel metal2 s 534170 0 534226 800 6 la_data_in[120]
port 169 nsew signal input
rlabel metal2 s 537574 0 537630 800 6 la_data_in[121]
port 170 nsew signal input
rlabel metal2 s 541070 0 541126 800 6 la_data_in[122]
port 171 nsew signal input
rlabel metal2 s 544474 0 544530 800 6 la_data_in[123]
port 172 nsew signal input
rlabel metal2 s 547878 0 547934 800 6 la_data_in[124]
port 173 nsew signal input
rlabel metal2 s 551374 0 551430 800 6 la_data_in[125]
port 174 nsew signal input
rlabel metal2 s 554778 0 554834 800 6 la_data_in[126]
port 175 nsew signal input
rlabel metal2 s 558182 0 558238 800 6 la_data_in[127]
port 176 nsew signal input
rlabel metal2 s 163134 0 163190 800 6 la_data_in[12]
port 177 nsew signal input
rlabel metal2 s 166538 0 166594 800 6 la_data_in[13]
port 178 nsew signal input
rlabel metal2 s 170034 0 170090 800 6 la_data_in[14]
port 179 nsew signal input
rlabel metal2 s 173438 0 173494 800 6 la_data_in[15]
port 180 nsew signal input
rlabel metal2 s 176842 0 176898 800 6 la_data_in[16]
port 181 nsew signal input
rlabel metal2 s 180338 0 180394 800 6 la_data_in[17]
port 182 nsew signal input
rlabel metal2 s 183742 0 183798 800 6 la_data_in[18]
port 183 nsew signal input
rlabel metal2 s 187146 0 187202 800 6 la_data_in[19]
port 184 nsew signal input
rlabel metal2 s 125322 0 125378 800 6 la_data_in[1]
port 185 nsew signal input
rlabel metal2 s 190642 0 190698 800 6 la_data_in[20]
port 186 nsew signal input
rlabel metal2 s 194046 0 194102 800 6 la_data_in[21]
port 187 nsew signal input
rlabel metal2 s 197450 0 197506 800 6 la_data_in[22]
port 188 nsew signal input
rlabel metal2 s 200946 0 201002 800 6 la_data_in[23]
port 189 nsew signal input
rlabel metal2 s 204350 0 204406 800 6 la_data_in[24]
port 190 nsew signal input
rlabel metal2 s 207846 0 207902 800 6 la_data_in[25]
port 191 nsew signal input
rlabel metal2 s 211250 0 211306 800 6 la_data_in[26]
port 192 nsew signal input
rlabel metal2 s 214654 0 214710 800 6 la_data_in[27]
port 193 nsew signal input
rlabel metal2 s 218150 0 218206 800 6 la_data_in[28]
port 194 nsew signal input
rlabel metal2 s 221554 0 221610 800 6 la_data_in[29]
port 195 nsew signal input
rlabel metal2 s 128818 0 128874 800 6 la_data_in[2]
port 196 nsew signal input
rlabel metal2 s 224958 0 225014 800 6 la_data_in[30]
port 197 nsew signal input
rlabel metal2 s 228454 0 228510 800 6 la_data_in[31]
port 198 nsew signal input
rlabel metal2 s 231858 0 231914 800 6 la_data_in[32]
port 199 nsew signal input
rlabel metal2 s 235262 0 235318 800 6 la_data_in[33]
port 200 nsew signal input
rlabel metal2 s 238758 0 238814 800 6 la_data_in[34]
port 201 nsew signal input
rlabel metal2 s 242162 0 242218 800 6 la_data_in[35]
port 202 nsew signal input
rlabel metal2 s 245566 0 245622 800 6 la_data_in[36]
port 203 nsew signal input
rlabel metal2 s 249062 0 249118 800 6 la_data_in[37]
port 204 nsew signal input
rlabel metal2 s 252466 0 252522 800 6 la_data_in[38]
port 205 nsew signal input
rlabel metal2 s 255870 0 255926 800 6 la_data_in[39]
port 206 nsew signal input
rlabel metal2 s 132222 0 132278 800 6 la_data_in[3]
port 207 nsew signal input
rlabel metal2 s 259366 0 259422 800 6 la_data_in[40]
port 208 nsew signal input
rlabel metal2 s 262770 0 262826 800 6 la_data_in[41]
port 209 nsew signal input
rlabel metal2 s 266174 0 266230 800 6 la_data_in[42]
port 210 nsew signal input
rlabel metal2 s 269670 0 269726 800 6 la_data_in[43]
port 211 nsew signal input
rlabel metal2 s 273074 0 273130 800 6 la_data_in[44]
port 212 nsew signal input
rlabel metal2 s 276478 0 276534 800 6 la_data_in[45]
port 213 nsew signal input
rlabel metal2 s 279974 0 280030 800 6 la_data_in[46]
port 214 nsew signal input
rlabel metal2 s 283378 0 283434 800 6 la_data_in[47]
port 215 nsew signal input
rlabel metal2 s 286782 0 286838 800 6 la_data_in[48]
port 216 nsew signal input
rlabel metal2 s 290278 0 290334 800 6 la_data_in[49]
port 217 nsew signal input
rlabel metal2 s 135626 0 135682 800 6 la_data_in[4]
port 218 nsew signal input
rlabel metal2 s 293682 0 293738 800 6 la_data_in[50]
port 219 nsew signal input
rlabel metal2 s 297086 0 297142 800 6 la_data_in[51]
port 220 nsew signal input
rlabel metal2 s 300582 0 300638 800 6 la_data_in[52]
port 221 nsew signal input
rlabel metal2 s 303986 0 304042 800 6 la_data_in[53]
port 222 nsew signal input
rlabel metal2 s 307390 0 307446 800 6 la_data_in[54]
port 223 nsew signal input
rlabel metal2 s 310886 0 310942 800 6 la_data_in[55]
port 224 nsew signal input
rlabel metal2 s 314290 0 314346 800 6 la_data_in[56]
port 225 nsew signal input
rlabel metal2 s 317694 0 317750 800 6 la_data_in[57]
port 226 nsew signal input
rlabel metal2 s 321190 0 321246 800 6 la_data_in[58]
port 227 nsew signal input
rlabel metal2 s 324594 0 324650 800 6 la_data_in[59]
port 228 nsew signal input
rlabel metal2 s 139122 0 139178 800 6 la_data_in[5]
port 229 nsew signal input
rlabel metal2 s 328090 0 328146 800 6 la_data_in[60]
port 230 nsew signal input
rlabel metal2 s 331494 0 331550 800 6 la_data_in[61]
port 231 nsew signal input
rlabel metal2 s 334898 0 334954 800 6 la_data_in[62]
port 232 nsew signal input
rlabel metal2 s 338394 0 338450 800 6 la_data_in[63]
port 233 nsew signal input
rlabel metal2 s 341798 0 341854 800 6 la_data_in[64]
port 234 nsew signal input
rlabel metal2 s 345202 0 345258 800 6 la_data_in[65]
port 235 nsew signal input
rlabel metal2 s 348698 0 348754 800 6 la_data_in[66]
port 236 nsew signal input
rlabel metal2 s 352102 0 352158 800 6 la_data_in[67]
port 237 nsew signal input
rlabel metal2 s 355506 0 355562 800 6 la_data_in[68]
port 238 nsew signal input
rlabel metal2 s 359002 0 359058 800 6 la_data_in[69]
port 239 nsew signal input
rlabel metal2 s 142526 0 142582 800 6 la_data_in[6]
port 240 nsew signal input
rlabel metal2 s 362406 0 362462 800 6 la_data_in[70]
port 241 nsew signal input
rlabel metal2 s 365810 0 365866 800 6 la_data_in[71]
port 242 nsew signal input
rlabel metal2 s 369306 0 369362 800 6 la_data_in[72]
port 243 nsew signal input
rlabel metal2 s 372710 0 372766 800 6 la_data_in[73]
port 244 nsew signal input
rlabel metal2 s 376114 0 376170 800 6 la_data_in[74]
port 245 nsew signal input
rlabel metal2 s 379610 0 379666 800 6 la_data_in[75]
port 246 nsew signal input
rlabel metal2 s 383014 0 383070 800 6 la_data_in[76]
port 247 nsew signal input
rlabel metal2 s 386418 0 386474 800 6 la_data_in[77]
port 248 nsew signal input
rlabel metal2 s 389914 0 389970 800 6 la_data_in[78]
port 249 nsew signal input
rlabel metal2 s 393318 0 393374 800 6 la_data_in[79]
port 250 nsew signal input
rlabel metal2 s 145930 0 145986 800 6 la_data_in[7]
port 251 nsew signal input
rlabel metal2 s 396722 0 396778 800 6 la_data_in[80]
port 252 nsew signal input
rlabel metal2 s 400218 0 400274 800 6 la_data_in[81]
port 253 nsew signal input
rlabel metal2 s 403622 0 403678 800 6 la_data_in[82]
port 254 nsew signal input
rlabel metal2 s 407026 0 407082 800 6 la_data_in[83]
port 255 nsew signal input
rlabel metal2 s 410522 0 410578 800 6 la_data_in[84]
port 256 nsew signal input
rlabel metal2 s 413926 0 413982 800 6 la_data_in[85]
port 257 nsew signal input
rlabel metal2 s 417330 0 417386 800 6 la_data_in[86]
port 258 nsew signal input
rlabel metal2 s 420826 0 420882 800 6 la_data_in[87]
port 259 nsew signal input
rlabel metal2 s 424230 0 424286 800 6 la_data_in[88]
port 260 nsew signal input
rlabel metal2 s 427634 0 427690 800 6 la_data_in[89]
port 261 nsew signal input
rlabel metal2 s 149426 0 149482 800 6 la_data_in[8]
port 262 nsew signal input
rlabel metal2 s 431130 0 431186 800 6 la_data_in[90]
port 263 nsew signal input
rlabel metal2 s 434534 0 434590 800 6 la_data_in[91]
port 264 nsew signal input
rlabel metal2 s 437938 0 437994 800 6 la_data_in[92]
port 265 nsew signal input
rlabel metal2 s 441434 0 441490 800 6 la_data_in[93]
port 266 nsew signal input
rlabel metal2 s 444838 0 444894 800 6 la_data_in[94]
port 267 nsew signal input
rlabel metal2 s 448334 0 448390 800 6 la_data_in[95]
port 268 nsew signal input
rlabel metal2 s 451738 0 451794 800 6 la_data_in[96]
port 269 nsew signal input
rlabel metal2 s 455142 0 455198 800 6 la_data_in[97]
port 270 nsew signal input
rlabel metal2 s 458638 0 458694 800 6 la_data_in[98]
port 271 nsew signal input
rlabel metal2 s 462042 0 462098 800 6 la_data_in[99]
port 272 nsew signal input
rlabel metal2 s 152830 0 152886 800 6 la_data_in[9]
port 273 nsew signal input
rlabel metal2 s 123022 0 123078 800 6 la_data_out[0]
port 274 nsew signal output
rlabel metal2 s 466642 0 466698 800 6 la_data_out[100]
port 275 nsew signal output
rlabel metal2 s 470046 0 470102 800 6 la_data_out[101]
port 276 nsew signal output
rlabel metal2 s 473450 0 473506 800 6 la_data_out[102]
port 277 nsew signal output
rlabel metal2 s 476946 0 477002 800 6 la_data_out[103]
port 278 nsew signal output
rlabel metal2 s 480350 0 480406 800 6 la_data_out[104]
port 279 nsew signal output
rlabel metal2 s 483754 0 483810 800 6 la_data_out[105]
port 280 nsew signal output
rlabel metal2 s 487250 0 487306 800 6 la_data_out[106]
port 281 nsew signal output
rlabel metal2 s 490654 0 490710 800 6 la_data_out[107]
port 282 nsew signal output
rlabel metal2 s 494058 0 494114 800 6 la_data_out[108]
port 283 nsew signal output
rlabel metal2 s 497554 0 497610 800 6 la_data_out[109]
port 284 nsew signal output
rlabel metal2 s 157430 0 157486 800 6 la_data_out[10]
port 285 nsew signal output
rlabel metal2 s 500958 0 501014 800 6 la_data_out[110]
port 286 nsew signal output
rlabel metal2 s 504362 0 504418 800 6 la_data_out[111]
port 287 nsew signal output
rlabel metal2 s 507858 0 507914 800 6 la_data_out[112]
port 288 nsew signal output
rlabel metal2 s 511262 0 511318 800 6 la_data_out[113]
port 289 nsew signal output
rlabel metal2 s 514666 0 514722 800 6 la_data_out[114]
port 290 nsew signal output
rlabel metal2 s 518162 0 518218 800 6 la_data_out[115]
port 291 nsew signal output
rlabel metal2 s 521566 0 521622 800 6 la_data_out[116]
port 292 nsew signal output
rlabel metal2 s 524970 0 525026 800 6 la_data_out[117]
port 293 nsew signal output
rlabel metal2 s 528466 0 528522 800 6 la_data_out[118]
port 294 nsew signal output
rlabel metal2 s 531870 0 531926 800 6 la_data_out[119]
port 295 nsew signal output
rlabel metal2 s 160834 0 160890 800 6 la_data_out[11]
port 296 nsew signal output
rlabel metal2 s 535366 0 535422 800 6 la_data_out[120]
port 297 nsew signal output
rlabel metal2 s 538770 0 538826 800 6 la_data_out[121]
port 298 nsew signal output
rlabel metal2 s 542174 0 542230 800 6 la_data_out[122]
port 299 nsew signal output
rlabel metal2 s 545670 0 545726 800 6 la_data_out[123]
port 300 nsew signal output
rlabel metal2 s 549074 0 549130 800 6 la_data_out[124]
port 301 nsew signal output
rlabel metal2 s 552478 0 552534 800 6 la_data_out[125]
port 302 nsew signal output
rlabel metal2 s 555974 0 556030 800 6 la_data_out[126]
port 303 nsew signal output
rlabel metal2 s 559378 0 559434 800 6 la_data_out[127]
port 304 nsew signal output
rlabel metal2 s 164330 0 164386 800 6 la_data_out[12]
port 305 nsew signal output
rlabel metal2 s 167734 0 167790 800 6 la_data_out[13]
port 306 nsew signal output
rlabel metal2 s 171138 0 171194 800 6 la_data_out[14]
port 307 nsew signal output
rlabel metal2 s 174634 0 174690 800 6 la_data_out[15]
port 308 nsew signal output
rlabel metal2 s 178038 0 178094 800 6 la_data_out[16]
port 309 nsew signal output
rlabel metal2 s 181442 0 181498 800 6 la_data_out[17]
port 310 nsew signal output
rlabel metal2 s 184938 0 184994 800 6 la_data_out[18]
port 311 nsew signal output
rlabel metal2 s 188342 0 188398 800 6 la_data_out[19]
port 312 nsew signal output
rlabel metal2 s 126518 0 126574 800 6 la_data_out[1]
port 313 nsew signal output
rlabel metal2 s 191746 0 191802 800 6 la_data_out[20]
port 314 nsew signal output
rlabel metal2 s 195242 0 195298 800 6 la_data_out[21]
port 315 nsew signal output
rlabel metal2 s 198646 0 198702 800 6 la_data_out[22]
port 316 nsew signal output
rlabel metal2 s 202050 0 202106 800 6 la_data_out[23]
port 317 nsew signal output
rlabel metal2 s 205546 0 205602 800 6 la_data_out[24]
port 318 nsew signal output
rlabel metal2 s 208950 0 209006 800 6 la_data_out[25]
port 319 nsew signal output
rlabel metal2 s 212354 0 212410 800 6 la_data_out[26]
port 320 nsew signal output
rlabel metal2 s 215850 0 215906 800 6 la_data_out[27]
port 321 nsew signal output
rlabel metal2 s 219254 0 219310 800 6 la_data_out[28]
port 322 nsew signal output
rlabel metal2 s 222658 0 222714 800 6 la_data_out[29]
port 323 nsew signal output
rlabel metal2 s 129922 0 129978 800 6 la_data_out[2]
port 324 nsew signal output
rlabel metal2 s 226154 0 226210 800 6 la_data_out[30]
port 325 nsew signal output
rlabel metal2 s 229558 0 229614 800 6 la_data_out[31]
port 326 nsew signal output
rlabel metal2 s 232962 0 233018 800 6 la_data_out[32]
port 327 nsew signal output
rlabel metal2 s 236458 0 236514 800 6 la_data_out[33]
port 328 nsew signal output
rlabel metal2 s 239862 0 239918 800 6 la_data_out[34]
port 329 nsew signal output
rlabel metal2 s 243266 0 243322 800 6 la_data_out[35]
port 330 nsew signal output
rlabel metal2 s 246762 0 246818 800 6 la_data_out[36]
port 331 nsew signal output
rlabel metal2 s 250166 0 250222 800 6 la_data_out[37]
port 332 nsew signal output
rlabel metal2 s 253570 0 253626 800 6 la_data_out[38]
port 333 nsew signal output
rlabel metal2 s 257066 0 257122 800 6 la_data_out[39]
port 334 nsew signal output
rlabel metal2 s 133326 0 133382 800 6 la_data_out[3]
port 335 nsew signal output
rlabel metal2 s 260470 0 260526 800 6 la_data_out[40]
port 336 nsew signal output
rlabel metal2 s 263874 0 263930 800 6 la_data_out[41]
port 337 nsew signal output
rlabel metal2 s 267370 0 267426 800 6 la_data_out[42]
port 338 nsew signal output
rlabel metal2 s 270774 0 270830 800 6 la_data_out[43]
port 339 nsew signal output
rlabel metal2 s 274178 0 274234 800 6 la_data_out[44]
port 340 nsew signal output
rlabel metal2 s 277674 0 277730 800 6 la_data_out[45]
port 341 nsew signal output
rlabel metal2 s 281078 0 281134 800 6 la_data_out[46]
port 342 nsew signal output
rlabel metal2 s 284574 0 284630 800 6 la_data_out[47]
port 343 nsew signal output
rlabel metal2 s 287978 0 288034 800 6 la_data_out[48]
port 344 nsew signal output
rlabel metal2 s 291382 0 291438 800 6 la_data_out[49]
port 345 nsew signal output
rlabel metal2 s 136822 0 136878 800 6 la_data_out[4]
port 346 nsew signal output
rlabel metal2 s 294878 0 294934 800 6 la_data_out[50]
port 347 nsew signal output
rlabel metal2 s 298282 0 298338 800 6 la_data_out[51]
port 348 nsew signal output
rlabel metal2 s 301686 0 301742 800 6 la_data_out[52]
port 349 nsew signal output
rlabel metal2 s 305182 0 305238 800 6 la_data_out[53]
port 350 nsew signal output
rlabel metal2 s 308586 0 308642 800 6 la_data_out[54]
port 351 nsew signal output
rlabel metal2 s 311990 0 312046 800 6 la_data_out[55]
port 352 nsew signal output
rlabel metal2 s 315486 0 315542 800 6 la_data_out[56]
port 353 nsew signal output
rlabel metal2 s 318890 0 318946 800 6 la_data_out[57]
port 354 nsew signal output
rlabel metal2 s 322294 0 322350 800 6 la_data_out[58]
port 355 nsew signal output
rlabel metal2 s 325790 0 325846 800 6 la_data_out[59]
port 356 nsew signal output
rlabel metal2 s 140226 0 140282 800 6 la_data_out[5]
port 357 nsew signal output
rlabel metal2 s 329194 0 329250 800 6 la_data_out[60]
port 358 nsew signal output
rlabel metal2 s 332598 0 332654 800 6 la_data_out[61]
port 359 nsew signal output
rlabel metal2 s 336094 0 336150 800 6 la_data_out[62]
port 360 nsew signal output
rlabel metal2 s 339498 0 339554 800 6 la_data_out[63]
port 361 nsew signal output
rlabel metal2 s 342902 0 342958 800 6 la_data_out[64]
port 362 nsew signal output
rlabel metal2 s 346398 0 346454 800 6 la_data_out[65]
port 363 nsew signal output
rlabel metal2 s 349802 0 349858 800 6 la_data_out[66]
port 364 nsew signal output
rlabel metal2 s 353206 0 353262 800 6 la_data_out[67]
port 365 nsew signal output
rlabel metal2 s 356702 0 356758 800 6 la_data_out[68]
port 366 nsew signal output
rlabel metal2 s 360106 0 360162 800 6 la_data_out[69]
port 367 nsew signal output
rlabel metal2 s 143630 0 143686 800 6 la_data_out[6]
port 368 nsew signal output
rlabel metal2 s 363510 0 363566 800 6 la_data_out[70]
port 369 nsew signal output
rlabel metal2 s 367006 0 367062 800 6 la_data_out[71]
port 370 nsew signal output
rlabel metal2 s 370410 0 370466 800 6 la_data_out[72]
port 371 nsew signal output
rlabel metal2 s 373814 0 373870 800 6 la_data_out[73]
port 372 nsew signal output
rlabel metal2 s 377310 0 377366 800 6 la_data_out[74]
port 373 nsew signal output
rlabel metal2 s 380714 0 380770 800 6 la_data_out[75]
port 374 nsew signal output
rlabel metal2 s 384118 0 384174 800 6 la_data_out[76]
port 375 nsew signal output
rlabel metal2 s 387614 0 387670 800 6 la_data_out[77]
port 376 nsew signal output
rlabel metal2 s 391018 0 391074 800 6 la_data_out[78]
port 377 nsew signal output
rlabel metal2 s 394422 0 394478 800 6 la_data_out[79]
port 378 nsew signal output
rlabel metal2 s 147126 0 147182 800 6 la_data_out[7]
port 379 nsew signal output
rlabel metal2 s 397918 0 397974 800 6 la_data_out[80]
port 380 nsew signal output
rlabel metal2 s 401322 0 401378 800 6 la_data_out[81]
port 381 nsew signal output
rlabel metal2 s 404726 0 404782 800 6 la_data_out[82]
port 382 nsew signal output
rlabel metal2 s 408222 0 408278 800 6 la_data_out[83]
port 383 nsew signal output
rlabel metal2 s 411626 0 411682 800 6 la_data_out[84]
port 384 nsew signal output
rlabel metal2 s 415122 0 415178 800 6 la_data_out[85]
port 385 nsew signal output
rlabel metal2 s 418526 0 418582 800 6 la_data_out[86]
port 386 nsew signal output
rlabel metal2 s 421930 0 421986 800 6 la_data_out[87]
port 387 nsew signal output
rlabel metal2 s 425426 0 425482 800 6 la_data_out[88]
port 388 nsew signal output
rlabel metal2 s 428830 0 428886 800 6 la_data_out[89]
port 389 nsew signal output
rlabel metal2 s 150530 0 150586 800 6 la_data_out[8]
port 390 nsew signal output
rlabel metal2 s 432234 0 432290 800 6 la_data_out[90]
port 391 nsew signal output
rlabel metal2 s 435730 0 435786 800 6 la_data_out[91]
port 392 nsew signal output
rlabel metal2 s 439134 0 439190 800 6 la_data_out[92]
port 393 nsew signal output
rlabel metal2 s 442538 0 442594 800 6 la_data_out[93]
port 394 nsew signal output
rlabel metal2 s 446034 0 446090 800 6 la_data_out[94]
port 395 nsew signal output
rlabel metal2 s 449438 0 449494 800 6 la_data_out[95]
port 396 nsew signal output
rlabel metal2 s 452842 0 452898 800 6 la_data_out[96]
port 397 nsew signal output
rlabel metal2 s 456338 0 456394 800 6 la_data_out[97]
port 398 nsew signal output
rlabel metal2 s 459742 0 459798 800 6 la_data_out[98]
port 399 nsew signal output
rlabel metal2 s 463146 0 463202 800 6 la_data_out[99]
port 400 nsew signal output
rlabel metal2 s 153934 0 153990 800 6 la_data_out[9]
port 401 nsew signal output
rlabel metal2 s 124218 0 124274 800 6 la_oen[0]
port 402 nsew signal input
rlabel metal2 s 467746 0 467802 800 6 la_oen[100]
port 403 nsew signal input
rlabel metal2 s 471150 0 471206 800 6 la_oen[101]
port 404 nsew signal input
rlabel metal2 s 474646 0 474702 800 6 la_oen[102]
port 405 nsew signal input
rlabel metal2 s 478050 0 478106 800 6 la_oen[103]
port 406 nsew signal input
rlabel metal2 s 481454 0 481510 800 6 la_oen[104]
port 407 nsew signal input
rlabel metal2 s 484950 0 485006 800 6 la_oen[105]
port 408 nsew signal input
rlabel metal2 s 488354 0 488410 800 6 la_oen[106]
port 409 nsew signal input
rlabel metal2 s 491850 0 491906 800 6 la_oen[107]
port 410 nsew signal input
rlabel metal2 s 495254 0 495310 800 6 la_oen[108]
port 411 nsew signal input
rlabel metal2 s 498658 0 498714 800 6 la_oen[109]
port 412 nsew signal input
rlabel metal2 s 158534 0 158590 800 6 la_oen[10]
port 413 nsew signal input
rlabel metal2 s 502154 0 502210 800 6 la_oen[110]
port 414 nsew signal input
rlabel metal2 s 505558 0 505614 800 6 la_oen[111]
port 415 nsew signal input
rlabel metal2 s 508962 0 509018 800 6 la_oen[112]
port 416 nsew signal input
rlabel metal2 s 512458 0 512514 800 6 la_oen[113]
port 417 nsew signal input
rlabel metal2 s 515862 0 515918 800 6 la_oen[114]
port 418 nsew signal input
rlabel metal2 s 519266 0 519322 800 6 la_oen[115]
port 419 nsew signal input
rlabel metal2 s 522762 0 522818 800 6 la_oen[116]
port 420 nsew signal input
rlabel metal2 s 526166 0 526222 800 6 la_oen[117]
port 421 nsew signal input
rlabel metal2 s 529570 0 529626 800 6 la_oen[118]
port 422 nsew signal input
rlabel metal2 s 533066 0 533122 800 6 la_oen[119]
port 423 nsew signal input
rlabel metal2 s 162030 0 162086 800 6 la_oen[11]
port 424 nsew signal input
rlabel metal2 s 536470 0 536526 800 6 la_oen[120]
port 425 nsew signal input
rlabel metal2 s 539874 0 539930 800 6 la_oen[121]
port 426 nsew signal input
rlabel metal2 s 543370 0 543426 800 6 la_oen[122]
port 427 nsew signal input
rlabel metal2 s 546774 0 546830 800 6 la_oen[123]
port 428 nsew signal input
rlabel metal2 s 550178 0 550234 800 6 la_oen[124]
port 429 nsew signal input
rlabel metal2 s 553674 0 553730 800 6 la_oen[125]
port 430 nsew signal input
rlabel metal2 s 557078 0 557134 800 6 la_oen[126]
port 431 nsew signal input
rlabel metal2 s 560482 0 560538 800 6 la_oen[127]
port 432 nsew signal input
rlabel metal2 s 165434 0 165490 800 6 la_oen[12]
port 433 nsew signal input
rlabel metal2 s 168838 0 168894 800 6 la_oen[13]
port 434 nsew signal input
rlabel metal2 s 172334 0 172390 800 6 la_oen[14]
port 435 nsew signal input
rlabel metal2 s 175738 0 175794 800 6 la_oen[15]
port 436 nsew signal input
rlabel metal2 s 179142 0 179198 800 6 la_oen[16]
port 437 nsew signal input
rlabel metal2 s 182638 0 182694 800 6 la_oen[17]
port 438 nsew signal input
rlabel metal2 s 186042 0 186098 800 6 la_oen[18]
port 439 nsew signal input
rlabel metal2 s 189446 0 189502 800 6 la_oen[19]
port 440 nsew signal input
rlabel metal2 s 127622 0 127678 800 6 la_oen[1]
port 441 nsew signal input
rlabel metal2 s 192942 0 192998 800 6 la_oen[20]
port 442 nsew signal input
rlabel metal2 s 196346 0 196402 800 6 la_oen[21]
port 443 nsew signal input
rlabel metal2 s 199750 0 199806 800 6 la_oen[22]
port 444 nsew signal input
rlabel metal2 s 203246 0 203302 800 6 la_oen[23]
port 445 nsew signal input
rlabel metal2 s 206650 0 206706 800 6 la_oen[24]
port 446 nsew signal input
rlabel metal2 s 210054 0 210110 800 6 la_oen[25]
port 447 nsew signal input
rlabel metal2 s 213550 0 213606 800 6 la_oen[26]
port 448 nsew signal input
rlabel metal2 s 216954 0 217010 800 6 la_oen[27]
port 449 nsew signal input
rlabel metal2 s 220358 0 220414 800 6 la_oen[28]
port 450 nsew signal input
rlabel metal2 s 223854 0 223910 800 6 la_oen[29]
port 451 nsew signal input
rlabel metal2 s 131118 0 131174 800 6 la_oen[2]
port 452 nsew signal input
rlabel metal2 s 227258 0 227314 800 6 la_oen[30]
port 453 nsew signal input
rlabel metal2 s 230662 0 230718 800 6 la_oen[31]
port 454 nsew signal input
rlabel metal2 s 234158 0 234214 800 6 la_oen[32]
port 455 nsew signal input
rlabel metal2 s 237562 0 237618 800 6 la_oen[33]
port 456 nsew signal input
rlabel metal2 s 240966 0 241022 800 6 la_oen[34]
port 457 nsew signal input
rlabel metal2 s 244462 0 244518 800 6 la_oen[35]
port 458 nsew signal input
rlabel metal2 s 247866 0 247922 800 6 la_oen[36]
port 459 nsew signal input
rlabel metal2 s 251362 0 251418 800 6 la_oen[37]
port 460 nsew signal input
rlabel metal2 s 254766 0 254822 800 6 la_oen[38]
port 461 nsew signal input
rlabel metal2 s 258170 0 258226 800 6 la_oen[39]
port 462 nsew signal input
rlabel metal2 s 134522 0 134578 800 6 la_oen[3]
port 463 nsew signal input
rlabel metal2 s 261666 0 261722 800 6 la_oen[40]
port 464 nsew signal input
rlabel metal2 s 265070 0 265126 800 6 la_oen[41]
port 465 nsew signal input
rlabel metal2 s 268474 0 268530 800 6 la_oen[42]
port 466 nsew signal input
rlabel metal2 s 271970 0 272026 800 6 la_oen[43]
port 467 nsew signal input
rlabel metal2 s 275374 0 275430 800 6 la_oen[44]
port 468 nsew signal input
rlabel metal2 s 278778 0 278834 800 6 la_oen[45]
port 469 nsew signal input
rlabel metal2 s 282274 0 282330 800 6 la_oen[46]
port 470 nsew signal input
rlabel metal2 s 285678 0 285734 800 6 la_oen[47]
port 471 nsew signal input
rlabel metal2 s 289082 0 289138 800 6 la_oen[48]
port 472 nsew signal input
rlabel metal2 s 292578 0 292634 800 6 la_oen[49]
port 473 nsew signal input
rlabel metal2 s 137926 0 137982 800 6 la_oen[4]
port 474 nsew signal input
rlabel metal2 s 295982 0 296038 800 6 la_oen[50]
port 475 nsew signal input
rlabel metal2 s 299386 0 299442 800 6 la_oen[51]
port 476 nsew signal input
rlabel metal2 s 302882 0 302938 800 6 la_oen[52]
port 477 nsew signal input
rlabel metal2 s 306286 0 306342 800 6 la_oen[53]
port 478 nsew signal input
rlabel metal2 s 309690 0 309746 800 6 la_oen[54]
port 479 nsew signal input
rlabel metal2 s 313186 0 313242 800 6 la_oen[55]
port 480 nsew signal input
rlabel metal2 s 316590 0 316646 800 6 la_oen[56]
port 481 nsew signal input
rlabel metal2 s 319994 0 320050 800 6 la_oen[57]
port 482 nsew signal input
rlabel metal2 s 323490 0 323546 800 6 la_oen[58]
port 483 nsew signal input
rlabel metal2 s 326894 0 326950 800 6 la_oen[59]
port 484 nsew signal input
rlabel metal2 s 141422 0 141478 800 6 la_oen[5]
port 485 nsew signal input
rlabel metal2 s 330298 0 330354 800 6 la_oen[60]
port 486 nsew signal input
rlabel metal2 s 333794 0 333850 800 6 la_oen[61]
port 487 nsew signal input
rlabel metal2 s 337198 0 337254 800 6 la_oen[62]
port 488 nsew signal input
rlabel metal2 s 340602 0 340658 800 6 la_oen[63]
port 489 nsew signal input
rlabel metal2 s 344098 0 344154 800 6 la_oen[64]
port 490 nsew signal input
rlabel metal2 s 347502 0 347558 800 6 la_oen[65]
port 491 nsew signal input
rlabel metal2 s 350906 0 350962 800 6 la_oen[66]
port 492 nsew signal input
rlabel metal2 s 354402 0 354458 800 6 la_oen[67]
port 493 nsew signal input
rlabel metal2 s 357806 0 357862 800 6 la_oen[68]
port 494 nsew signal input
rlabel metal2 s 361210 0 361266 800 6 la_oen[69]
port 495 nsew signal input
rlabel metal2 s 144826 0 144882 800 6 la_oen[6]
port 496 nsew signal input
rlabel metal2 s 364706 0 364762 800 6 la_oen[70]
port 497 nsew signal input
rlabel metal2 s 368110 0 368166 800 6 la_oen[71]
port 498 nsew signal input
rlabel metal2 s 371606 0 371662 800 6 la_oen[72]
port 499 nsew signal input
rlabel metal2 s 375010 0 375066 800 6 la_oen[73]
port 500 nsew signal input
rlabel metal2 s 378414 0 378470 800 6 la_oen[74]
port 501 nsew signal input
rlabel metal2 s 381910 0 381966 800 6 la_oen[75]
port 502 nsew signal input
rlabel metal2 s 385314 0 385370 800 6 la_oen[76]
port 503 nsew signal input
rlabel metal2 s 388718 0 388774 800 6 la_oen[77]
port 504 nsew signal input
rlabel metal2 s 392214 0 392270 800 6 la_oen[78]
port 505 nsew signal input
rlabel metal2 s 395618 0 395674 800 6 la_oen[79]
port 506 nsew signal input
rlabel metal2 s 148230 0 148286 800 6 la_oen[7]
port 507 nsew signal input
rlabel metal2 s 399022 0 399078 800 6 la_oen[80]
port 508 nsew signal input
rlabel metal2 s 402518 0 402574 800 6 la_oen[81]
port 509 nsew signal input
rlabel metal2 s 405922 0 405978 800 6 la_oen[82]
port 510 nsew signal input
rlabel metal2 s 409326 0 409382 800 6 la_oen[83]
port 511 nsew signal input
rlabel metal2 s 412822 0 412878 800 6 la_oen[84]
port 512 nsew signal input
rlabel metal2 s 416226 0 416282 800 6 la_oen[85]
port 513 nsew signal input
rlabel metal2 s 419630 0 419686 800 6 la_oen[86]
port 514 nsew signal input
rlabel metal2 s 423126 0 423182 800 6 la_oen[87]
port 515 nsew signal input
rlabel metal2 s 426530 0 426586 800 6 la_oen[88]
port 516 nsew signal input
rlabel metal2 s 429934 0 429990 800 6 la_oen[89]
port 517 nsew signal input
rlabel metal2 s 151726 0 151782 800 6 la_oen[8]
port 518 nsew signal input
rlabel metal2 s 433430 0 433486 800 6 la_oen[90]
port 519 nsew signal input
rlabel metal2 s 436834 0 436890 800 6 la_oen[91]
port 520 nsew signal input
rlabel metal2 s 440238 0 440294 800 6 la_oen[92]
port 521 nsew signal input
rlabel metal2 s 443734 0 443790 800 6 la_oen[93]
port 522 nsew signal input
rlabel metal2 s 447138 0 447194 800 6 la_oen[94]
port 523 nsew signal input
rlabel metal2 s 450542 0 450598 800 6 la_oen[95]
port 524 nsew signal input
rlabel metal2 s 454038 0 454094 800 6 la_oen[96]
port 525 nsew signal input
rlabel metal2 s 457442 0 457498 800 6 la_oen[97]
port 526 nsew signal input
rlabel metal2 s 460846 0 460902 800 6 la_oen[98]
port 527 nsew signal input
rlabel metal2 s 464342 0 464398 800 6 la_oen[99]
port 528 nsew signal input
rlabel metal2 s 155130 0 155186 800 6 la_oen[9]
port 529 nsew signal input
rlabel metal2 s 561678 0 561734 800 6 user_clock2
port 530 nsew signal input
rlabel metal2 s 570 0 626 800 6 wb_clk_i
port 531 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wb_rst_i
port 532 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 wbs_ack_o
port 533 nsew signal output
rlabel metal2 s 7378 0 7434 800 6 wbs_adr_i[0]
port 534 nsew signal input
rlabel metal2 s 46294 0 46350 800 6 wbs_adr_i[10]
port 535 nsew signal input
rlabel metal2 s 49790 0 49846 800 6 wbs_adr_i[11]
port 536 nsew signal input
rlabel metal2 s 53194 0 53250 800 6 wbs_adr_i[12]
port 537 nsew signal input
rlabel metal2 s 56598 0 56654 800 6 wbs_adr_i[13]
port 538 nsew signal input
rlabel metal2 s 60094 0 60150 800 6 wbs_adr_i[14]
port 539 nsew signal input
rlabel metal2 s 63498 0 63554 800 6 wbs_adr_i[15]
port 540 nsew signal input
rlabel metal2 s 66902 0 66958 800 6 wbs_adr_i[16]
port 541 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 wbs_adr_i[17]
port 542 nsew signal input
rlabel metal2 s 73802 0 73858 800 6 wbs_adr_i[18]
port 543 nsew signal input
rlabel metal2 s 77206 0 77262 800 6 wbs_adr_i[19]
port 544 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 wbs_adr_i[1]
port 545 nsew signal input
rlabel metal2 s 80702 0 80758 800 6 wbs_adr_i[20]
port 546 nsew signal input
rlabel metal2 s 84106 0 84162 800 6 wbs_adr_i[21]
port 547 nsew signal input
rlabel metal2 s 87602 0 87658 800 6 wbs_adr_i[22]
port 548 nsew signal input
rlabel metal2 s 91006 0 91062 800 6 wbs_adr_i[23]
port 549 nsew signal input
rlabel metal2 s 94410 0 94466 800 6 wbs_adr_i[24]
port 550 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 wbs_adr_i[25]
port 551 nsew signal input
rlabel metal2 s 101310 0 101366 800 6 wbs_adr_i[26]
port 552 nsew signal input
rlabel metal2 s 104714 0 104770 800 6 wbs_adr_i[27]
port 553 nsew signal input
rlabel metal2 s 108210 0 108266 800 6 wbs_adr_i[28]
port 554 nsew signal input
rlabel metal2 s 111614 0 111670 800 6 wbs_adr_i[29]
port 555 nsew signal input
rlabel metal2 s 16578 0 16634 800 6 wbs_adr_i[2]
port 556 nsew signal input
rlabel metal2 s 115018 0 115074 800 6 wbs_adr_i[30]
port 557 nsew signal input
rlabel metal2 s 118514 0 118570 800 6 wbs_adr_i[31]
port 558 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 wbs_adr_i[3]
port 559 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 wbs_adr_i[4]
port 560 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 wbs_adr_i[5]
port 561 nsew signal input
rlabel metal2 s 32586 0 32642 800 6 wbs_adr_i[6]
port 562 nsew signal input
rlabel metal2 s 35990 0 36046 800 6 wbs_adr_i[7]
port 563 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 wbs_adr_i[8]
port 564 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 wbs_adr_i[9]
port 565 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 wbs_cyc_i
port 566 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 wbs_dat_i[0]
port 567 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 wbs_dat_i[10]
port 568 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 wbs_dat_i[11]
port 569 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 wbs_dat_i[12]
port 570 nsew signal input
rlabel metal2 s 57794 0 57850 800 6 wbs_dat_i[13]
port 571 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 wbs_dat_i[14]
port 572 nsew signal input
rlabel metal2 s 64694 0 64750 800 6 wbs_dat_i[15]
port 573 nsew signal input
rlabel metal2 s 68098 0 68154 800 6 wbs_dat_i[16]
port 574 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 wbs_dat_i[17]
port 575 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 wbs_dat_i[18]
port 576 nsew signal input
rlabel metal2 s 78402 0 78458 800 6 wbs_dat_i[19]
port 577 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 wbs_dat_i[1]
port 578 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 wbs_dat_i[20]
port 579 nsew signal input
rlabel metal2 s 85302 0 85358 800 6 wbs_dat_i[21]
port 580 nsew signal input
rlabel metal2 s 88706 0 88762 800 6 wbs_dat_i[22]
port 581 nsew signal input
rlabel metal2 s 92110 0 92166 800 6 wbs_dat_i[23]
port 582 nsew signal input
rlabel metal2 s 95606 0 95662 800 6 wbs_dat_i[24]
port 583 nsew signal input
rlabel metal2 s 99010 0 99066 800 6 wbs_dat_i[25]
port 584 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 wbs_dat_i[26]
port 585 nsew signal input
rlabel metal2 s 105910 0 105966 800 6 wbs_dat_i[27]
port 586 nsew signal input
rlabel metal2 s 109314 0 109370 800 6 wbs_dat_i[28]
port 587 nsew signal input
rlabel metal2 s 112718 0 112774 800 6 wbs_dat_i[29]
port 588 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 wbs_dat_i[2]
port 589 nsew signal input
rlabel metal2 s 116214 0 116270 800 6 wbs_dat_i[30]
port 590 nsew signal input
rlabel metal2 s 119618 0 119674 800 6 wbs_dat_i[31]
port 591 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 wbs_dat_i[3]
port 592 nsew signal input
rlabel metal2 s 26882 0 26938 800 6 wbs_dat_i[4]
port 593 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 wbs_dat_i[5]
port 594 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 wbs_dat_i[6]
port 595 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 wbs_dat_i[7]
port 596 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 wbs_dat_i[8]
port 597 nsew signal input
rlabel metal2 s 44086 0 44142 800 6 wbs_dat_i[9]
port 598 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 wbs_dat_o[0]
port 599 nsew signal output
rlabel metal2 s 48594 0 48650 800 6 wbs_dat_o[10]
port 600 nsew signal output
rlabel metal2 s 52090 0 52146 800 6 wbs_dat_o[11]
port 601 nsew signal output
rlabel metal2 s 55494 0 55550 800 6 wbs_dat_o[12]
port 602 nsew signal output
rlabel metal2 s 58898 0 58954 800 6 wbs_dat_o[13]
port 603 nsew signal output
rlabel metal2 s 62394 0 62450 800 6 wbs_dat_o[14]
port 604 nsew signal output
rlabel metal2 s 65798 0 65854 800 6 wbs_dat_o[15]
port 605 nsew signal output
rlabel metal2 s 69202 0 69258 800 6 wbs_dat_o[16]
port 606 nsew signal output
rlabel metal2 s 72698 0 72754 800 6 wbs_dat_o[17]
port 607 nsew signal output
rlabel metal2 s 76102 0 76158 800 6 wbs_dat_o[18]
port 608 nsew signal output
rlabel metal2 s 79506 0 79562 800 6 wbs_dat_o[19]
port 609 nsew signal output
rlabel metal2 s 14278 0 14334 800 6 wbs_dat_o[1]
port 610 nsew signal output
rlabel metal2 s 83002 0 83058 800 6 wbs_dat_o[20]
port 611 nsew signal output
rlabel metal2 s 86406 0 86462 800 6 wbs_dat_o[21]
port 612 nsew signal output
rlabel metal2 s 89810 0 89866 800 6 wbs_dat_o[22]
port 613 nsew signal output
rlabel metal2 s 93306 0 93362 800 6 wbs_dat_o[23]
port 614 nsew signal output
rlabel metal2 s 96710 0 96766 800 6 wbs_dat_o[24]
port 615 nsew signal output
rlabel metal2 s 100114 0 100170 800 6 wbs_dat_o[25]
port 616 nsew signal output
rlabel metal2 s 103610 0 103666 800 6 wbs_dat_o[26]
port 617 nsew signal output
rlabel metal2 s 107014 0 107070 800 6 wbs_dat_o[27]
port 618 nsew signal output
rlabel metal2 s 110418 0 110474 800 6 wbs_dat_o[28]
port 619 nsew signal output
rlabel metal2 s 113914 0 113970 800 6 wbs_dat_o[29]
port 620 nsew signal output
rlabel metal2 s 18878 0 18934 800 6 wbs_dat_o[2]
port 621 nsew signal output
rlabel metal2 s 117318 0 117374 800 6 wbs_dat_o[30]
port 622 nsew signal output
rlabel metal2 s 120722 0 120778 800 6 wbs_dat_o[31]
port 623 nsew signal output
rlabel metal2 s 23386 0 23442 800 6 wbs_dat_o[3]
port 624 nsew signal output
rlabel metal2 s 27986 0 28042 800 6 wbs_dat_o[4]
port 625 nsew signal output
rlabel metal2 s 31482 0 31538 800 6 wbs_dat_o[5]
port 626 nsew signal output
rlabel metal2 s 34886 0 34942 800 6 wbs_dat_o[6]
port 627 nsew signal output
rlabel metal2 s 38290 0 38346 800 6 wbs_dat_o[7]
port 628 nsew signal output
rlabel metal2 s 41786 0 41842 800 6 wbs_dat_o[8]
port 629 nsew signal output
rlabel metal2 s 45190 0 45246 800 6 wbs_dat_o[9]
port 630 nsew signal output
rlabel metal2 s 10874 0 10930 800 6 wbs_sel_i[0]
port 631 nsew signal input
rlabel metal2 s 15382 0 15438 800 6 wbs_sel_i[1]
port 632 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 wbs_sel_i[2]
port 633 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 wbs_sel_i[3]
port 634 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 wbs_stb_i
port 635 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 wbs_we_i
port 636 nsew signal input
rlabel metal4 s 557168 2128 557488 685488 6 VPWR
port 637 nsew power bidirectional
rlabel metal4 s 526448 2128 526768 685488 6 VPWR
port 638 nsew power bidirectional
rlabel metal4 s 495728 2128 496048 685488 6 VPWR
port 639 nsew power bidirectional
rlabel metal4 s 465008 2128 465328 685488 6 VPWR
port 640 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 685488 6 VPWR
port 641 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 685488 6 VPWR
port 642 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 685488 6 VPWR
port 643 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 685488 6 VPWR
port 644 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 685488 6 VPWR
port 645 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 685488 6 VPWR
port 646 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 685488 6 VPWR
port 647 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 685488 6 VPWR
port 648 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 685488 6 VPWR
port 649 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 685488 6 VPWR
port 650 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 685488 6 VPWR
port 651 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 685488 6 VPWR
port 652 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 685488 6 VPWR
port 653 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 685488 6 VPWR
port 654 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 685488 6 VPWR
port 655 nsew power bidirectional
rlabel metal4 s 541808 2128 542128 685488 6 VGND
port 656 nsew ground bidirectional
rlabel metal4 s 511088 2128 511408 685488 6 VGND
port 657 nsew ground bidirectional
rlabel metal4 s 480368 2128 480688 685488 6 VGND
port 658 nsew ground bidirectional
rlabel metal4 s 449648 2128 449968 685488 6 VGND
port 659 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 685488 6 VGND
port 660 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 685488 6 VGND
port 661 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 685488 6 VGND
port 662 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 685488 6 VGND
port 663 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 685488 6 VGND
port 664 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 685488 6 VGND
port 665 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 685488 6 VGND
port 666 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 685488 6 VGND
port 667 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 685488 6 VGND
port 668 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 685488 6 VGND
port 669 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 685488 6 VGND
port 670 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 685488 6 VGND
port 671 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 685488 6 VGND
port 672 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 685488 6 VGND
port 673 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 568000 688000
string LEFview TRUE
<< end >>

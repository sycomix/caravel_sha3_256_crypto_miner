magic
tech sky130A
magscale 1 2
timestamp 1610260563
<< locali >>
rect 249717 699703 249751 701641
rect 260791 699873 260849 699907
rect 269129 699703 269163 699805
rect 136557 698071 136591 698173
rect 153209 697935 153243 698173
rect 157993 697935 158027 698105
rect 6101 696711 6135 696813
rect 19349 696779 19383 696881
rect 28917 696711 28951 696881
rect 165629 696779 165663 696881
rect 128369 696711 128403 696745
rect 128311 696677 128403 696711
rect 113097 696439 113131 696541
rect 116593 696439 116627 696541
rect 143733 696303 143767 696405
rect 160109 696371 160143 696405
rect 160051 696337 160143 696371
rect 8033 694943 8067 695045
rect 14013 694943 14047 695181
rect 15025 695181 15243 695215
rect 15025 695079 15059 695181
rect 15209 695079 15243 695181
rect 29561 694195 29595 695249
rect 43729 694263 43763 695249
rect 67465 694399 67499 695249
rect 81265 694467 81299 696201
rect 86417 694535 86451 695249
rect 95801 694671 95835 695249
rect 103471 695181 103563 695215
rect 103529 695147 103563 695181
rect 109969 694807 110003 695249
rect 124137 694875 124171 695249
rect 128921 694943 128955 695249
rect 138489 695011 138523 695249
rect 125609 694739 125643 694909
rect 140605 694739 140639 695249
rect 144963 695181 145021 695215
rect 152473 694739 152507 695249
rect 171517 695215 171551 699669
rect 186237 699227 186271 699669
rect 267565 699227 267599 699669
rect 269037 699635 269071 699669
rect 269221 699635 269255 699805
rect 273269 699703 273303 701029
rect 269037 699601 269255 699635
rect 273361 699363 273395 699669
rect 273303 699329 273395 699363
rect 237515 698377 237573 698411
rect 218195 698309 218345 698343
rect 237423 698309 237665 698343
rect 237515 698241 237757 698275
rect 215159 698173 215217 698207
rect 186329 698139 186363 698173
rect 172529 697935 172563 698105
rect 186271 698105 186363 698139
rect 193263 698105 193321 698139
rect 218103 698105 218253 698139
rect 237515 698105 237757 698139
rect 182097 697935 182131 698105
rect 237423 698037 237665 698071
rect 277593 696915 277627 701029
rect 296821 699771 296855 699873
rect 302249 699669 302433 699703
rect 282963 699329 283055 699363
rect 283021 698955 283055 699329
rect 302249 699227 302283 699669
rect 311817 699227 311851 699737
rect 316233 699703 316267 700009
rect 303353 699193 303571 699227
rect 303353 698955 303387 699193
rect 303537 699159 303571 699193
rect 305285 699193 305469 699227
rect 305285 699159 305319 699193
rect 321569 699159 321603 699873
rect 326353 699703 326387 700009
rect 331229 699771 331263 699873
rect 331229 699737 331321 699771
rect 335277 699703 335311 700009
rect 335921 699193 336139 699227
rect 303445 698955 303479 699125
rect 335921 698955 335955 699193
rect 336105 699159 336139 699193
rect 340797 699159 340831 699737
rect 344661 699227 344695 699737
rect 344753 699159 344787 699805
rect 344937 699227 344971 699873
rect 345029 699703 345063 699873
rect 345121 699703 345155 699805
rect 354781 699431 354815 699669
rect 364165 699431 364199 699669
rect 364257 699431 364291 699805
rect 336013 698955 336047 699125
rect 344845 698955 344879 699125
rect 354689 698207 354723 699397
rect 364441 699227 364475 699669
rect 373825 699227 373859 699669
rect 374101 699227 374135 699669
rect 383485 699227 383519 699669
rect 383761 699363 383795 699669
rect 383669 698275 383703 699329
rect 175197 696711 175231 696881
rect 224969 696779 225003 696881
rect 207063 696745 207155 696779
rect 253949 696779 253983 696881
rect 263609 696779 263643 696881
rect 271429 696779 271463 696881
rect 284953 696779 284987 696881
rect 289829 696779 289863 696881
rect 207121 696711 207155 696745
rect 208535 696609 208685 696643
rect 208443 696541 208777 696575
rect 302249 696371 302283 696881
rect 205683 696337 205741 696371
rect 311817 696371 311851 696881
rect 321569 696371 321603 696881
rect 331137 696371 331171 696881
rect 340889 696371 340923 696881
rect 350457 696371 350491 696881
rect 355333 696371 355367 696813
rect 364993 696371 365027 696813
rect 371157 696371 371191 696745
rect 563437 696167 563471 696269
rect 164249 695181 164341 695215
rect 164249 695147 164283 695181
rect 355609 694739 355643 695453
rect 364993 694739 365027 695453
rect 374653 694739 374687 695385
rect 384313 694739 384347 695385
rect 393973 694739 394007 695317
rect 403633 694739 403667 695317
rect 413293 694739 413327 695317
rect 422953 694739 422987 695317
rect 432613 694739 432647 695385
rect 440709 695079 440743 695317
rect 442273 694739 442307 695385
rect 483397 695079 483431 695317
rect 450277 694739 450311 695045
rect 459937 694739 459971 695045
rect 469597 694739 469631 695045
rect 497565 694603 497599 695317
rect 511917 694331 511951 695317
rect 412557 6443 412591 6613
rect 489469 6103 489503 6341
rect 538505 3383 538539 4029
rect 538999 3485 539241 3519
rect 541817 2975 541851 3553
rect 545405 3519 545439 4029
rect 547705 3927 547739 4165
rect 547797 3587 547831 3893
rect 547981 3655 548015 4165
rect 552707 3689 552799 3723
rect 547739 3553 547831 3587
rect 544209 3111 544243 3417
rect 547889 3111 547923 3621
rect 552765 3519 552799 3689
rect 547981 2635 548015 3009
rect 552673 2907 552707 3485
rect 558193 3111 558227 4029
rect 558285 3927 558319 4029
rect 559665 3383 559699 3417
rect 562057 3383 562091 3893
rect 563253 3587 563287 4165
rect 558285 3349 558469 3383
rect 559665 3349 559849 3383
rect 558101 3043 558135 3077
rect 558285 3043 558319 3349
rect 558101 3009 558319 3043
rect 560861 2975 560895 3077
rect 564449 2975 564483 3553
rect 567117 3179 567151 3553
rect 560861 2941 561137 2975
rect 560769 2635 560803 2941
rect 566841 2907 566875 3077
rect 565645 2635 565679 2873
<< viali >>
rect 249717 701641 249751 701675
rect 273269 701029 273303 701063
rect 260757 699873 260791 699907
rect 260849 699873 260883 699907
rect 269129 699805 269163 699839
rect 171517 699669 171551 699703
rect 136557 698173 136591 698207
rect 136557 698037 136591 698071
rect 153209 698173 153243 698207
rect 153209 697901 153243 697935
rect 157993 698105 158027 698139
rect 157993 697901 158027 697935
rect 19349 696881 19383 696915
rect 6101 696813 6135 696847
rect 19349 696745 19383 696779
rect 28917 696881 28951 696915
rect 6101 696677 6135 696711
rect 165629 696881 165663 696915
rect 128369 696745 128403 696779
rect 165629 696745 165663 696779
rect 28917 696677 28951 696711
rect 128277 696677 128311 696711
rect 113097 696541 113131 696575
rect 113097 696405 113131 696439
rect 116593 696541 116627 696575
rect 116593 696405 116627 696439
rect 143733 696405 143767 696439
rect 160109 696405 160143 696439
rect 160017 696337 160051 696371
rect 143733 696269 143767 696303
rect 81265 696201 81299 696235
rect 29561 695249 29595 695283
rect 14013 695181 14047 695215
rect 8033 695045 8067 695079
rect 8033 694909 8067 694943
rect 15025 695045 15059 695079
rect 15209 695045 15243 695079
rect 14013 694909 14047 694943
rect 43729 695249 43763 695283
rect 67465 695249 67499 695283
rect 86417 695249 86451 695283
rect 95801 695249 95835 695283
rect 109969 695249 110003 695283
rect 103437 695181 103471 695215
rect 103529 695113 103563 695147
rect 124137 695249 124171 695283
rect 128921 695249 128955 695283
rect 138489 695249 138523 695283
rect 138489 694977 138523 695011
rect 140605 695249 140639 695283
rect 124137 694841 124171 694875
rect 125609 694909 125643 694943
rect 128921 694909 128955 694943
rect 109969 694773 110003 694807
rect 125609 694705 125643 694739
rect 152473 695249 152507 695283
rect 144929 695181 144963 695215
rect 145021 695181 145055 695215
rect 140605 694705 140639 694739
rect 186237 699669 186271 699703
rect 249717 699669 249751 699703
rect 267565 699669 267599 699703
rect 186237 699193 186271 699227
rect 269037 699669 269071 699703
rect 269129 699669 269163 699703
rect 269221 699805 269255 699839
rect 277593 701029 277627 701063
rect 273269 699669 273303 699703
rect 273361 699669 273395 699703
rect 273269 699329 273303 699363
rect 267565 699193 267599 699227
rect 237481 698377 237515 698411
rect 237573 698377 237607 698411
rect 218161 698309 218195 698343
rect 218345 698309 218379 698343
rect 237389 698309 237423 698343
rect 237665 698309 237699 698343
rect 237481 698241 237515 698275
rect 237757 698241 237791 698275
rect 186329 698173 186363 698207
rect 215125 698173 215159 698207
rect 215217 698173 215251 698207
rect 172529 698105 172563 698139
rect 172529 697901 172563 697935
rect 182097 698105 182131 698139
rect 186237 698105 186271 698139
rect 193229 698105 193263 698139
rect 193321 698105 193355 698139
rect 218069 698105 218103 698139
rect 218253 698105 218287 698139
rect 237481 698105 237515 698139
rect 237757 698105 237791 698139
rect 237389 698037 237423 698071
rect 237665 698037 237699 698071
rect 182097 697901 182131 697935
rect 316233 700009 316267 700043
rect 296821 699873 296855 699907
rect 296821 699737 296855 699771
rect 311817 699737 311851 699771
rect 302433 699669 302467 699703
rect 282929 699329 282963 699363
rect 326353 700009 326387 700043
rect 316233 699669 316267 699703
rect 321569 699873 321603 699907
rect 302249 699193 302283 699227
rect 283021 698921 283055 698955
rect 303353 698921 303387 698955
rect 303445 699125 303479 699159
rect 303537 699125 303571 699159
rect 305469 699193 305503 699227
rect 311817 699193 311851 699227
rect 305285 699125 305319 699159
rect 335277 700009 335311 700043
rect 331229 699873 331263 699907
rect 331321 699737 331355 699771
rect 326353 699669 326387 699703
rect 344937 699873 344971 699907
rect 344753 699805 344787 699839
rect 335277 699669 335311 699703
rect 340797 699737 340831 699771
rect 321569 699125 321603 699159
rect 303445 698921 303479 698955
rect 335921 698921 335955 698955
rect 336013 699125 336047 699159
rect 336105 699125 336139 699159
rect 344661 699737 344695 699771
rect 344661 699193 344695 699227
rect 340797 699125 340831 699159
rect 345029 699873 345063 699907
rect 345029 699669 345063 699703
rect 345121 699805 345155 699839
rect 364257 699805 364291 699839
rect 345121 699669 345155 699703
rect 354781 699669 354815 699703
rect 344937 699193 344971 699227
rect 354689 699397 354723 699431
rect 354781 699397 354815 699431
rect 364165 699669 364199 699703
rect 364165 699397 364199 699431
rect 364257 699397 364291 699431
rect 364441 699669 364475 699703
rect 344753 699125 344787 699159
rect 344845 699125 344879 699159
rect 336013 698921 336047 698955
rect 344845 698921 344879 698955
rect 364441 699193 364475 699227
rect 373825 699669 373859 699703
rect 373825 699193 373859 699227
rect 374101 699669 374135 699703
rect 374101 699193 374135 699227
rect 383485 699669 383519 699703
rect 383761 699669 383795 699703
rect 383485 699193 383519 699227
rect 383669 699329 383703 699363
rect 383761 699329 383795 699363
rect 383669 698241 383703 698275
rect 354689 698173 354723 698207
rect 175197 696881 175231 696915
rect 224969 696881 225003 696915
rect 207029 696745 207063 696779
rect 224969 696745 225003 696779
rect 253949 696881 253983 696915
rect 253949 696745 253983 696779
rect 263609 696881 263643 696915
rect 263609 696745 263643 696779
rect 271429 696881 271463 696915
rect 277593 696881 277627 696915
rect 284953 696881 284987 696915
rect 271429 696745 271463 696779
rect 284953 696745 284987 696779
rect 289829 696881 289863 696915
rect 289829 696745 289863 696779
rect 302249 696881 302283 696915
rect 175197 696677 175231 696711
rect 207121 696677 207155 696711
rect 208501 696609 208535 696643
rect 208685 696609 208719 696643
rect 208409 696541 208443 696575
rect 208777 696541 208811 696575
rect 205649 696337 205683 696371
rect 205741 696337 205775 696371
rect 302249 696337 302283 696371
rect 311817 696881 311851 696915
rect 311817 696337 311851 696371
rect 321569 696881 321603 696915
rect 321569 696337 321603 696371
rect 331137 696881 331171 696915
rect 331137 696337 331171 696371
rect 340889 696881 340923 696915
rect 340889 696337 340923 696371
rect 350457 696881 350491 696915
rect 350457 696337 350491 696371
rect 355333 696813 355367 696847
rect 355333 696337 355367 696371
rect 364993 696813 365027 696847
rect 364993 696337 365027 696371
rect 371157 696745 371191 696779
rect 371157 696337 371191 696371
rect 563437 696269 563471 696303
rect 563437 696133 563471 696167
rect 164341 695181 164375 695215
rect 171517 695181 171551 695215
rect 355609 695453 355643 695487
rect 164249 695113 164283 695147
rect 152473 694705 152507 694739
rect 355609 694705 355643 694739
rect 364993 695453 365027 695487
rect 364993 694705 365027 694739
rect 374653 695385 374687 695419
rect 374653 694705 374687 694739
rect 384313 695385 384347 695419
rect 432613 695385 432647 695419
rect 384313 694705 384347 694739
rect 393973 695317 394007 695351
rect 393973 694705 394007 694739
rect 403633 695317 403667 695351
rect 403633 694705 403667 694739
rect 413293 695317 413327 695351
rect 413293 694705 413327 694739
rect 422953 695317 422987 695351
rect 422953 694705 422987 694739
rect 442273 695385 442307 695419
rect 440709 695317 440743 695351
rect 440709 695045 440743 695079
rect 432613 694705 432647 694739
rect 483397 695317 483431 695351
rect 442273 694705 442307 694739
rect 450277 695045 450311 695079
rect 450277 694705 450311 694739
rect 459937 695045 459971 695079
rect 459937 694705 459971 694739
rect 469597 695045 469631 695079
rect 483397 695045 483431 695079
rect 497565 695317 497599 695351
rect 469597 694705 469631 694739
rect 95801 694637 95835 694671
rect 497565 694569 497599 694603
rect 511917 695317 511951 695351
rect 86417 694501 86451 694535
rect 81265 694433 81299 694467
rect 67465 694365 67499 694399
rect 511917 694297 511951 694331
rect 43729 694229 43763 694263
rect 29561 694161 29595 694195
rect 412557 6613 412591 6647
rect 412557 6409 412591 6443
rect 489469 6341 489503 6375
rect 489469 6069 489503 6103
rect 547705 4165 547739 4199
rect 538505 4029 538539 4063
rect 545405 4029 545439 4063
rect 541817 3553 541851 3587
rect 538965 3485 538999 3519
rect 539241 3485 539275 3519
rect 538505 3349 538539 3383
rect 547981 4165 548015 4199
rect 547705 3893 547739 3927
rect 547797 3893 547831 3927
rect 563253 4165 563287 4199
rect 558193 4029 558227 4063
rect 552673 3689 552707 3723
rect 547705 3553 547739 3587
rect 547889 3621 547923 3655
rect 547981 3621 548015 3655
rect 545405 3485 545439 3519
rect 544209 3417 544243 3451
rect 544209 3077 544243 3111
rect 547889 3077 547923 3111
rect 552673 3485 552707 3519
rect 552765 3485 552799 3519
rect 541817 2941 541851 2975
rect 547981 3009 548015 3043
rect 558285 4029 558319 4063
rect 558285 3893 558319 3927
rect 562057 3893 562091 3927
rect 559665 3417 559699 3451
rect 563253 3553 563287 3587
rect 564449 3553 564483 3587
rect 558101 3077 558135 3111
rect 558193 3077 558227 3111
rect 558469 3349 558503 3383
rect 559849 3349 559883 3383
rect 562057 3349 562091 3383
rect 560861 3077 560895 3111
rect 567117 3553 567151 3587
rect 567117 3145 567151 3179
rect 552673 2873 552707 2907
rect 560769 2941 560803 2975
rect 561137 2941 561171 2975
rect 564449 2941 564483 2975
rect 566841 3077 566875 3111
rect 547981 2601 548015 2635
rect 560769 2601 560803 2635
rect 565645 2873 565679 2907
rect 566841 2873 566875 2907
rect 565645 2601 565679 2635
<< metal1 >>
rect 251634 701972 251640 702024
rect 251692 702012 251698 702024
rect 429838 702012 429844 702024
rect 251692 701984 429844 702012
rect 251692 701972 251698 701984
rect 429838 701972 429844 701984
rect 429896 701972 429902 702024
rect 237466 701904 237472 701956
rect 237524 701944 237530 701956
rect 494790 701944 494796 701956
rect 237524 701916 494796 701944
rect 237524 701904 237530 701916
rect 494790 701904 494796 701916
rect 494848 701904 494854 701956
rect 223298 701836 223304 701888
rect 223356 701876 223362 701888
rect 559650 701876 559656 701888
rect 223356 701848 559656 701876
rect 223356 701836 223362 701848
rect 559650 701836 559656 701848
rect 559708 701836 559714 701888
rect 1104 701786 582820 701808
rect 1104 701734 36822 701786
rect 36874 701734 36886 701786
rect 36938 701734 36950 701786
rect 37002 701734 37014 701786
rect 37066 701734 37078 701786
rect 37130 701734 37142 701786
rect 37194 701734 37206 701786
rect 37258 701734 37270 701786
rect 37322 701734 37334 701786
rect 37386 701734 72822 701786
rect 72874 701734 72886 701786
rect 72938 701734 72950 701786
rect 73002 701734 73014 701786
rect 73066 701734 73078 701786
rect 73130 701734 73142 701786
rect 73194 701734 73206 701786
rect 73258 701734 73270 701786
rect 73322 701734 73334 701786
rect 73386 701734 108822 701786
rect 108874 701734 108886 701786
rect 108938 701734 108950 701786
rect 109002 701734 109014 701786
rect 109066 701734 109078 701786
rect 109130 701734 109142 701786
rect 109194 701734 109206 701786
rect 109258 701734 109270 701786
rect 109322 701734 109334 701786
rect 109386 701734 144822 701786
rect 144874 701734 144886 701786
rect 144938 701734 144950 701786
rect 145002 701734 145014 701786
rect 145066 701734 145078 701786
rect 145130 701734 145142 701786
rect 145194 701734 145206 701786
rect 145258 701734 145270 701786
rect 145322 701734 145334 701786
rect 145386 701734 180822 701786
rect 180874 701734 180886 701786
rect 180938 701734 180950 701786
rect 181002 701734 181014 701786
rect 181066 701734 181078 701786
rect 181130 701734 181142 701786
rect 181194 701734 181206 701786
rect 181258 701734 181270 701786
rect 181322 701734 181334 701786
rect 181386 701734 216822 701786
rect 216874 701734 216886 701786
rect 216938 701734 216950 701786
rect 217002 701734 217014 701786
rect 217066 701734 217078 701786
rect 217130 701734 217142 701786
rect 217194 701734 217206 701786
rect 217258 701734 217270 701786
rect 217322 701734 217334 701786
rect 217386 701734 252822 701786
rect 252874 701734 252886 701786
rect 252938 701734 252950 701786
rect 253002 701734 253014 701786
rect 253066 701734 253078 701786
rect 253130 701734 253142 701786
rect 253194 701734 253206 701786
rect 253258 701734 253270 701786
rect 253322 701734 253334 701786
rect 253386 701734 288822 701786
rect 288874 701734 288886 701786
rect 288938 701734 288950 701786
rect 289002 701734 289014 701786
rect 289066 701734 289078 701786
rect 289130 701734 289142 701786
rect 289194 701734 289206 701786
rect 289258 701734 289270 701786
rect 289322 701734 289334 701786
rect 289386 701734 324822 701786
rect 324874 701734 324886 701786
rect 324938 701734 324950 701786
rect 325002 701734 325014 701786
rect 325066 701734 325078 701786
rect 325130 701734 325142 701786
rect 325194 701734 325206 701786
rect 325258 701734 325270 701786
rect 325322 701734 325334 701786
rect 325386 701734 360822 701786
rect 360874 701734 360886 701786
rect 360938 701734 360950 701786
rect 361002 701734 361014 701786
rect 361066 701734 361078 701786
rect 361130 701734 361142 701786
rect 361194 701734 361206 701786
rect 361258 701734 361270 701786
rect 361322 701734 361334 701786
rect 361386 701734 396822 701786
rect 396874 701734 396886 701786
rect 396938 701734 396950 701786
rect 397002 701734 397014 701786
rect 397066 701734 397078 701786
rect 397130 701734 397142 701786
rect 397194 701734 397206 701786
rect 397258 701734 397270 701786
rect 397322 701734 397334 701786
rect 397386 701734 432822 701786
rect 432874 701734 432886 701786
rect 432938 701734 432950 701786
rect 433002 701734 433014 701786
rect 433066 701734 433078 701786
rect 433130 701734 433142 701786
rect 433194 701734 433206 701786
rect 433258 701734 433270 701786
rect 433322 701734 433334 701786
rect 433386 701734 468822 701786
rect 468874 701734 468886 701786
rect 468938 701734 468950 701786
rect 469002 701734 469014 701786
rect 469066 701734 469078 701786
rect 469130 701734 469142 701786
rect 469194 701734 469206 701786
rect 469258 701734 469270 701786
rect 469322 701734 469334 701786
rect 469386 701734 504822 701786
rect 504874 701734 504886 701786
rect 504938 701734 504950 701786
rect 505002 701734 505014 701786
rect 505066 701734 505078 701786
rect 505130 701734 505142 701786
rect 505194 701734 505206 701786
rect 505258 701734 505270 701786
rect 505322 701734 505334 701786
rect 505386 701734 540822 701786
rect 540874 701734 540886 701786
rect 540938 701734 540950 701786
rect 541002 701734 541014 701786
rect 541066 701734 541078 701786
rect 541130 701734 541142 701786
rect 541194 701734 541206 701786
rect 541258 701734 541270 701786
rect 541322 701734 541334 701786
rect 541386 701734 576822 701786
rect 576874 701734 576886 701786
rect 576938 701734 576950 701786
rect 577002 701734 577014 701786
rect 577066 701734 577078 701786
rect 577130 701734 577142 701786
rect 577194 701734 577206 701786
rect 577258 701734 577270 701786
rect 577322 701734 577334 701786
rect 577386 701734 582820 701786
rect 1104 701712 582820 701734
rect 235166 701632 235172 701684
rect 235224 701672 235230 701684
rect 249705 701675 249763 701681
rect 249705 701672 249717 701675
rect 235224 701644 249717 701672
rect 235224 701632 235230 701644
rect 249705 701641 249717 701644
rect 249751 701641 249763 701675
rect 249705 701635 249763 701641
rect 1104 701242 582820 701264
rect 1104 701190 18822 701242
rect 18874 701190 18886 701242
rect 18938 701190 18950 701242
rect 19002 701190 19014 701242
rect 19066 701190 19078 701242
rect 19130 701190 19142 701242
rect 19194 701190 19206 701242
rect 19258 701190 19270 701242
rect 19322 701190 19334 701242
rect 19386 701190 54822 701242
rect 54874 701190 54886 701242
rect 54938 701190 54950 701242
rect 55002 701190 55014 701242
rect 55066 701190 55078 701242
rect 55130 701190 55142 701242
rect 55194 701190 55206 701242
rect 55258 701190 55270 701242
rect 55322 701190 55334 701242
rect 55386 701190 90822 701242
rect 90874 701190 90886 701242
rect 90938 701190 90950 701242
rect 91002 701190 91014 701242
rect 91066 701190 91078 701242
rect 91130 701190 91142 701242
rect 91194 701190 91206 701242
rect 91258 701190 91270 701242
rect 91322 701190 91334 701242
rect 91386 701190 126822 701242
rect 126874 701190 126886 701242
rect 126938 701190 126950 701242
rect 127002 701190 127014 701242
rect 127066 701190 127078 701242
rect 127130 701190 127142 701242
rect 127194 701190 127206 701242
rect 127258 701190 127270 701242
rect 127322 701190 127334 701242
rect 127386 701190 162822 701242
rect 162874 701190 162886 701242
rect 162938 701190 162950 701242
rect 163002 701190 163014 701242
rect 163066 701190 163078 701242
rect 163130 701190 163142 701242
rect 163194 701190 163206 701242
rect 163258 701190 163270 701242
rect 163322 701190 163334 701242
rect 163386 701190 198822 701242
rect 198874 701190 198886 701242
rect 198938 701190 198950 701242
rect 199002 701190 199014 701242
rect 199066 701190 199078 701242
rect 199130 701190 199142 701242
rect 199194 701190 199206 701242
rect 199258 701190 199270 701242
rect 199322 701190 199334 701242
rect 199386 701190 234822 701242
rect 234874 701190 234886 701242
rect 234938 701190 234950 701242
rect 235002 701190 235014 701242
rect 235066 701190 235078 701242
rect 235130 701190 235142 701242
rect 235194 701190 235206 701242
rect 235258 701190 235270 701242
rect 235322 701190 235334 701242
rect 235386 701190 270822 701242
rect 270874 701190 270886 701242
rect 270938 701190 270950 701242
rect 271002 701190 271014 701242
rect 271066 701190 271078 701242
rect 271130 701190 271142 701242
rect 271194 701190 271206 701242
rect 271258 701190 271270 701242
rect 271322 701190 271334 701242
rect 271386 701190 306822 701242
rect 306874 701190 306886 701242
rect 306938 701190 306950 701242
rect 307002 701190 307014 701242
rect 307066 701190 307078 701242
rect 307130 701190 307142 701242
rect 307194 701190 307206 701242
rect 307258 701190 307270 701242
rect 307322 701190 307334 701242
rect 307386 701190 342822 701242
rect 342874 701190 342886 701242
rect 342938 701190 342950 701242
rect 343002 701190 343014 701242
rect 343066 701190 343078 701242
rect 343130 701190 343142 701242
rect 343194 701190 343206 701242
rect 343258 701190 343270 701242
rect 343322 701190 343334 701242
rect 343386 701190 378822 701242
rect 378874 701190 378886 701242
rect 378938 701190 378950 701242
rect 379002 701190 379014 701242
rect 379066 701190 379078 701242
rect 379130 701190 379142 701242
rect 379194 701190 379206 701242
rect 379258 701190 379270 701242
rect 379322 701190 379334 701242
rect 379386 701190 414822 701242
rect 414874 701190 414886 701242
rect 414938 701190 414950 701242
rect 415002 701190 415014 701242
rect 415066 701190 415078 701242
rect 415130 701190 415142 701242
rect 415194 701190 415206 701242
rect 415258 701190 415270 701242
rect 415322 701190 415334 701242
rect 415386 701190 450822 701242
rect 450874 701190 450886 701242
rect 450938 701190 450950 701242
rect 451002 701190 451014 701242
rect 451066 701190 451078 701242
rect 451130 701190 451142 701242
rect 451194 701190 451206 701242
rect 451258 701190 451270 701242
rect 451322 701190 451334 701242
rect 451386 701190 486822 701242
rect 486874 701190 486886 701242
rect 486938 701190 486950 701242
rect 487002 701190 487014 701242
rect 487066 701190 487078 701242
rect 487130 701190 487142 701242
rect 487194 701190 487206 701242
rect 487258 701190 487270 701242
rect 487322 701190 487334 701242
rect 487386 701190 522822 701242
rect 522874 701190 522886 701242
rect 522938 701190 522950 701242
rect 523002 701190 523014 701242
rect 523066 701190 523078 701242
rect 523130 701190 523142 701242
rect 523194 701190 523206 701242
rect 523258 701190 523270 701242
rect 523322 701190 523334 701242
rect 523386 701190 558822 701242
rect 558874 701190 558886 701242
rect 558938 701190 558950 701242
rect 559002 701190 559014 701242
rect 559066 701190 559078 701242
rect 559130 701190 559142 701242
rect 559194 701190 559206 701242
rect 559258 701190 559270 701242
rect 559322 701190 559334 701242
rect 559386 701190 582820 701242
rect 1104 701168 582820 701190
rect 273257 701063 273315 701069
rect 273257 701029 273269 701063
rect 273303 701060 273315 701063
rect 277581 701063 277639 701069
rect 277581 701060 277593 701063
rect 273303 701032 277593 701060
rect 273303 701029 273315 701032
rect 273257 701023 273315 701029
rect 277581 701029 277593 701032
rect 277627 701029 277639 701063
rect 277581 701023 277639 701029
rect 261110 700952 261116 701004
rect 261168 700992 261174 701004
rect 413646 700992 413652 701004
rect 261168 700964 413652 700992
rect 261168 700952 261174 700964
rect 413646 700952 413652 700964
rect 413704 700952 413710 701004
rect 154114 700884 154120 700936
rect 154172 700924 154178 700936
rect 317966 700924 317972 700936
rect 154172 700896 317972 700924
rect 154172 700884 154178 700896
rect 317966 700884 317972 700896
rect 318024 700884 318030 700936
rect 137830 700816 137836 700868
rect 137888 700856 137894 700868
rect 313182 700856 313188 700868
rect 137888 700828 313188 700856
rect 137888 700816 137894 700828
rect 313182 700816 313188 700828
rect 313240 700816 313246 700868
rect 105446 700748 105452 700800
rect 105504 700788 105510 700800
rect 322658 700788 322664 700800
rect 105504 700760 322664 700788
rect 105504 700748 105510 700760
rect 322658 700748 322664 700760
rect 322716 700748 322722 700800
rect 1104 700698 582820 700720
rect 1104 700646 36822 700698
rect 36874 700646 36886 700698
rect 36938 700646 36950 700698
rect 37002 700646 37014 700698
rect 37066 700646 37078 700698
rect 37130 700646 37142 700698
rect 37194 700646 37206 700698
rect 37258 700646 37270 700698
rect 37322 700646 37334 700698
rect 37386 700646 72822 700698
rect 72874 700646 72886 700698
rect 72938 700646 72950 700698
rect 73002 700646 73014 700698
rect 73066 700646 73078 700698
rect 73130 700646 73142 700698
rect 73194 700646 73206 700698
rect 73258 700646 73270 700698
rect 73322 700646 73334 700698
rect 73386 700646 108822 700698
rect 108874 700646 108886 700698
rect 108938 700646 108950 700698
rect 109002 700646 109014 700698
rect 109066 700646 109078 700698
rect 109130 700646 109142 700698
rect 109194 700646 109206 700698
rect 109258 700646 109270 700698
rect 109322 700646 109334 700698
rect 109386 700646 144822 700698
rect 144874 700646 144886 700698
rect 144938 700646 144950 700698
rect 145002 700646 145014 700698
rect 145066 700646 145078 700698
rect 145130 700646 145142 700698
rect 145194 700646 145206 700698
rect 145258 700646 145270 700698
rect 145322 700646 145334 700698
rect 145386 700646 180822 700698
rect 180874 700646 180886 700698
rect 180938 700646 180950 700698
rect 181002 700646 181014 700698
rect 181066 700646 181078 700698
rect 181130 700646 181142 700698
rect 181194 700646 181206 700698
rect 181258 700646 181270 700698
rect 181322 700646 181334 700698
rect 181386 700646 216822 700698
rect 216874 700646 216886 700698
rect 216938 700646 216950 700698
rect 217002 700646 217014 700698
rect 217066 700646 217078 700698
rect 217130 700646 217142 700698
rect 217194 700646 217206 700698
rect 217258 700646 217270 700698
rect 217322 700646 217334 700698
rect 217386 700646 252822 700698
rect 252874 700646 252886 700698
rect 252938 700646 252950 700698
rect 253002 700646 253014 700698
rect 253066 700646 253078 700698
rect 253130 700646 253142 700698
rect 253194 700646 253206 700698
rect 253258 700646 253270 700698
rect 253322 700646 253334 700698
rect 253386 700646 288822 700698
rect 288874 700646 288886 700698
rect 288938 700646 288950 700698
rect 289002 700646 289014 700698
rect 289066 700646 289078 700698
rect 289130 700646 289142 700698
rect 289194 700646 289206 700698
rect 289258 700646 289270 700698
rect 289322 700646 289334 700698
rect 289386 700646 324822 700698
rect 324874 700646 324886 700698
rect 324938 700646 324950 700698
rect 325002 700646 325014 700698
rect 325066 700646 325078 700698
rect 325130 700646 325142 700698
rect 325194 700646 325206 700698
rect 325258 700646 325270 700698
rect 325322 700646 325334 700698
rect 325386 700646 360822 700698
rect 360874 700646 360886 700698
rect 360938 700646 360950 700698
rect 361002 700646 361014 700698
rect 361066 700646 361078 700698
rect 361130 700646 361142 700698
rect 361194 700646 361206 700698
rect 361258 700646 361270 700698
rect 361322 700646 361334 700698
rect 361386 700646 396822 700698
rect 396874 700646 396886 700698
rect 396938 700646 396950 700698
rect 397002 700646 397014 700698
rect 397066 700646 397078 700698
rect 397130 700646 397142 700698
rect 397194 700646 397206 700698
rect 397258 700646 397270 700698
rect 397322 700646 397334 700698
rect 397386 700646 432822 700698
rect 432874 700646 432886 700698
rect 432938 700646 432950 700698
rect 433002 700646 433014 700698
rect 433066 700646 433078 700698
rect 433130 700646 433142 700698
rect 433194 700646 433206 700698
rect 433258 700646 433270 700698
rect 433322 700646 433334 700698
rect 433386 700646 468822 700698
rect 468874 700646 468886 700698
rect 468938 700646 468950 700698
rect 469002 700646 469014 700698
rect 469066 700646 469078 700698
rect 469130 700646 469142 700698
rect 469194 700646 469206 700698
rect 469258 700646 469270 700698
rect 469322 700646 469334 700698
rect 469386 700646 504822 700698
rect 504874 700646 504886 700698
rect 504938 700646 504950 700698
rect 505002 700646 505014 700698
rect 505066 700646 505078 700698
rect 505130 700646 505142 700698
rect 505194 700646 505206 700698
rect 505258 700646 505270 700698
rect 505322 700646 505334 700698
rect 505386 700646 540822 700698
rect 540874 700646 540886 700698
rect 540938 700646 540950 700698
rect 541002 700646 541014 700698
rect 541066 700646 541078 700698
rect 541130 700646 541142 700698
rect 541194 700646 541206 700698
rect 541258 700646 541270 700698
rect 541322 700646 541334 700698
rect 541386 700646 576822 700698
rect 576874 700646 576886 700698
rect 576938 700646 576950 700698
rect 577002 700646 577014 700698
rect 577066 700646 577078 700698
rect 577130 700646 577142 700698
rect 577194 700646 577206 700698
rect 577258 700646 577270 700698
rect 577322 700646 577334 700698
rect 577386 700646 582820 700698
rect 1104 700624 582820 700646
rect 242250 700544 242256 700596
rect 242308 700584 242314 700596
rect 462314 700584 462320 700596
rect 242308 700556 462320 700584
rect 242308 700544 242314 700556
rect 462314 700544 462320 700556
rect 462372 700544 462378 700596
rect 246942 700476 246948 700528
rect 247000 700516 247006 700528
rect 478506 700516 478512 700528
rect 247000 700488 478512 700516
rect 247000 700476 247006 700488
rect 478506 700476 478512 700488
rect 478564 700476 478570 700528
rect 89162 700408 89168 700460
rect 89220 700448 89226 700460
rect 332134 700448 332140 700460
rect 89220 700420 332140 700448
rect 89220 700408 89226 700420
rect 332134 700408 332140 700420
rect 332192 700408 332198 700460
rect 202782 700340 202788 700392
rect 202840 700380 202846 700392
rect 296530 700380 296536 700392
rect 202840 700352 296536 700380
rect 202840 700340 202846 700352
rect 296530 700340 296536 700352
rect 296588 700340 296594 700392
rect 296622 700340 296628 700392
rect 296680 700380 296686 700392
rect 543458 700380 543464 700392
rect 296680 700352 543464 700380
rect 296680 700340 296686 700352
rect 543458 700340 543464 700352
rect 543516 700340 543522 700392
rect 72694 700272 72700 700324
rect 72752 700312 72758 700324
rect 327442 700312 327448 700324
rect 72752 700284 327448 700312
rect 72752 700272 72758 700284
rect 327442 700272 327448 700284
rect 327500 700272 327506 700324
rect 256418 700204 256424 700256
rect 256476 700244 256482 700256
rect 397454 700244 397460 700256
rect 256476 700216 397460 700244
rect 256476 700204 256482 700216
rect 397454 700204 397460 700216
rect 397512 700204 397518 700256
rect 1104 700154 582820 700176
rect 1104 700102 18822 700154
rect 18874 700102 18886 700154
rect 18938 700102 18950 700154
rect 19002 700102 19014 700154
rect 19066 700102 19078 700154
rect 19130 700102 19142 700154
rect 19194 700102 19206 700154
rect 19258 700102 19270 700154
rect 19322 700102 19334 700154
rect 19386 700102 54822 700154
rect 54874 700102 54886 700154
rect 54938 700102 54950 700154
rect 55002 700102 55014 700154
rect 55066 700102 55078 700154
rect 55130 700102 55142 700154
rect 55194 700102 55206 700154
rect 55258 700102 55270 700154
rect 55322 700102 55334 700154
rect 55386 700102 90822 700154
rect 90874 700102 90886 700154
rect 90938 700102 90950 700154
rect 91002 700102 91014 700154
rect 91066 700102 91078 700154
rect 91130 700102 91142 700154
rect 91194 700102 91206 700154
rect 91258 700102 91270 700154
rect 91322 700102 91334 700154
rect 91386 700102 126822 700154
rect 126874 700102 126886 700154
rect 126938 700102 126950 700154
rect 127002 700102 127014 700154
rect 127066 700102 127078 700154
rect 127130 700102 127142 700154
rect 127194 700102 127206 700154
rect 127258 700102 127270 700154
rect 127322 700102 127334 700154
rect 127386 700102 162822 700154
rect 162874 700102 162886 700154
rect 162938 700102 162950 700154
rect 163002 700102 163014 700154
rect 163066 700102 163078 700154
rect 163130 700102 163142 700154
rect 163194 700102 163206 700154
rect 163258 700102 163270 700154
rect 163322 700102 163334 700154
rect 163386 700102 198822 700154
rect 198874 700102 198886 700154
rect 198938 700102 198950 700154
rect 199002 700102 199014 700154
rect 199066 700102 199078 700154
rect 199130 700102 199142 700154
rect 199194 700102 199206 700154
rect 199258 700102 199270 700154
rect 199322 700102 199334 700154
rect 199386 700102 234822 700154
rect 234874 700102 234886 700154
rect 234938 700102 234950 700154
rect 235002 700102 235014 700154
rect 235066 700102 235078 700154
rect 235130 700102 235142 700154
rect 235194 700102 235206 700154
rect 235258 700102 235270 700154
rect 235322 700102 235334 700154
rect 235386 700102 270822 700154
rect 270874 700102 270886 700154
rect 270938 700102 270950 700154
rect 271002 700102 271014 700154
rect 271066 700102 271078 700154
rect 271130 700102 271142 700154
rect 271194 700102 271206 700154
rect 271258 700102 271270 700154
rect 271322 700102 271334 700154
rect 271386 700102 306822 700154
rect 306874 700102 306886 700154
rect 306938 700102 306950 700154
rect 307002 700102 307014 700154
rect 307066 700102 307078 700154
rect 307130 700102 307142 700154
rect 307194 700102 307206 700154
rect 307258 700102 307270 700154
rect 307322 700102 307334 700154
rect 307386 700102 342822 700154
rect 342874 700102 342886 700154
rect 342938 700102 342950 700154
rect 343002 700102 343014 700154
rect 343066 700102 343078 700154
rect 343130 700102 343142 700154
rect 343194 700102 343206 700154
rect 343258 700102 343270 700154
rect 343322 700102 343334 700154
rect 343386 700102 378822 700154
rect 378874 700102 378886 700154
rect 378938 700102 378950 700154
rect 379002 700102 379014 700154
rect 379066 700102 379078 700154
rect 379130 700102 379142 700154
rect 379194 700102 379206 700154
rect 379258 700102 379270 700154
rect 379322 700102 379334 700154
rect 379386 700102 414822 700154
rect 414874 700102 414886 700154
rect 414938 700102 414950 700154
rect 415002 700102 415014 700154
rect 415066 700102 415078 700154
rect 415130 700102 415142 700154
rect 415194 700102 415206 700154
rect 415258 700102 415270 700154
rect 415322 700102 415334 700154
rect 415386 700102 450822 700154
rect 450874 700102 450886 700154
rect 450938 700102 450950 700154
rect 451002 700102 451014 700154
rect 451066 700102 451078 700154
rect 451130 700102 451142 700154
rect 451194 700102 451206 700154
rect 451258 700102 451270 700154
rect 451322 700102 451334 700154
rect 451386 700102 486822 700154
rect 486874 700102 486886 700154
rect 486938 700102 486950 700154
rect 487002 700102 487014 700154
rect 487066 700102 487078 700154
rect 487130 700102 487142 700154
rect 487194 700102 487206 700154
rect 487258 700102 487270 700154
rect 487322 700102 487334 700154
rect 487386 700102 522822 700154
rect 522874 700102 522886 700154
rect 522938 700102 522950 700154
rect 523002 700102 523014 700154
rect 523066 700102 523078 700154
rect 523130 700102 523142 700154
rect 523194 700102 523206 700154
rect 523258 700102 523270 700154
rect 523322 700102 523334 700154
rect 523386 700102 558822 700154
rect 558874 700102 558886 700154
rect 558938 700102 558950 700154
rect 559002 700102 559014 700154
rect 559066 700102 559078 700154
rect 559130 700102 559142 700154
rect 559194 700102 559206 700154
rect 559258 700102 559270 700154
rect 559322 700102 559334 700154
rect 559386 700102 582820 700154
rect 1104 700080 582820 700102
rect 170306 700000 170312 700052
rect 170364 700040 170370 700052
rect 308490 700040 308496 700052
rect 170364 700012 308496 700040
rect 170364 700000 170370 700012
rect 308490 700000 308496 700012
rect 308548 700000 308554 700052
rect 308582 700000 308588 700052
rect 308640 700040 308646 700052
rect 316221 700043 316279 700049
rect 316221 700040 316233 700043
rect 308640 700012 316233 700040
rect 308640 700000 308646 700012
rect 316221 700009 316233 700012
rect 316267 700009 316279 700043
rect 316221 700003 316279 700009
rect 326341 700043 326399 700049
rect 326341 700009 326353 700043
rect 326387 700040 326399 700043
rect 335265 700043 335323 700049
rect 335265 700040 335277 700043
rect 326387 700012 335277 700040
rect 326387 700009 326399 700012
rect 326341 700003 326399 700009
rect 335265 700009 335277 700012
rect 335311 700009 335323 700043
rect 335265 700003 335323 700009
rect 265894 699932 265900 699984
rect 265952 699972 265958 699984
rect 364978 699972 364984 699984
rect 265952 699944 364984 699972
rect 265952 699932 265958 699944
rect 364978 699932 364984 699944
rect 365036 699932 365042 699984
rect 218974 699864 218980 699916
rect 219032 699904 219038 699916
rect 260745 699907 260803 699913
rect 260745 699904 260757 699907
rect 219032 699876 260757 699904
rect 219032 699864 219038 699876
rect 260745 699873 260757 699876
rect 260791 699873 260803 699907
rect 260745 699867 260803 699873
rect 260837 699907 260895 699913
rect 260837 699873 260849 699907
rect 260883 699904 260895 699907
rect 296714 699904 296720 699916
rect 260883 699876 296720 699904
rect 260883 699873 260895 699876
rect 260837 699867 260895 699873
rect 296714 699864 296720 699876
rect 296772 699864 296778 699916
rect 296809 699907 296867 699913
rect 296809 699873 296821 699907
rect 296855 699904 296867 699907
rect 298002 699904 298008 699916
rect 296855 699876 298008 699904
rect 296855 699873 296867 699876
rect 296809 699867 296867 699873
rect 298002 699864 298008 699876
rect 298060 699864 298066 699916
rect 321557 699907 321615 699913
rect 298756 699876 311940 699904
rect 251082 699796 251088 699848
rect 251140 699836 251146 699848
rect 251140 699808 259500 699836
rect 251140 699796 251146 699808
rect 259472 699780 259500 699808
rect 267642 699796 267648 699848
rect 267700 699836 267706 699848
rect 269117 699839 269175 699845
rect 269117 699836 269129 699839
rect 267700 699808 269129 699836
rect 267700 699796 267706 699808
rect 269117 699805 269129 699808
rect 269163 699805 269175 699839
rect 269117 699799 269175 699805
rect 269209 699839 269267 699845
rect 269209 699805 269221 699839
rect 269255 699836 269267 699839
rect 273254 699836 273260 699848
rect 269255 699808 273260 699836
rect 269255 699805 269267 699808
rect 269209 699799 269267 699805
rect 273254 699796 273260 699808
rect 273312 699796 273318 699848
rect 298756 699836 298784 699876
rect 273364 699808 298784 699836
rect 311912 699836 311940 699876
rect 321557 699873 321569 699907
rect 321603 699904 321615 699907
rect 331217 699907 331275 699913
rect 331217 699904 331229 699907
rect 321603 699876 331229 699904
rect 321603 699873 321615 699876
rect 321557 699867 321615 699873
rect 331217 699873 331229 699876
rect 331263 699873 331275 699907
rect 331217 699867 331275 699873
rect 331306 699864 331312 699916
rect 331364 699904 331370 699916
rect 344925 699907 344983 699913
rect 344925 699904 344937 699907
rect 331364 699876 344937 699904
rect 331364 699864 331370 699876
rect 344925 699873 344937 699876
rect 344971 699873 344983 699907
rect 344925 699867 344983 699873
rect 345017 699907 345075 699913
rect 345017 699873 345029 699907
rect 345063 699904 345075 699907
rect 348786 699904 348792 699916
rect 345063 699876 348792 699904
rect 345063 699873 345075 699876
rect 345017 699867 345075 699873
rect 348786 699864 348792 699876
rect 348844 699864 348850 699916
rect 332502 699836 332508 699848
rect 311912 699808 332508 699836
rect 259454 699728 259460 699780
rect 259512 699728 259518 699780
rect 270586 699728 270592 699780
rect 270644 699768 270650 699780
rect 273364 699768 273392 699808
rect 332502 699796 332508 699808
rect 332560 699796 332566 699848
rect 344741 699839 344799 699845
rect 344741 699805 344753 699839
rect 344787 699836 344799 699839
rect 345109 699839 345167 699845
rect 345109 699836 345121 699839
rect 344787 699808 345121 699836
rect 344787 699805 344799 699808
rect 344741 699799 344799 699805
rect 345109 699805 345121 699808
rect 345155 699805 345167 699839
rect 364245 699839 364303 699845
rect 364245 699836 364257 699839
rect 345109 699799 345167 699805
rect 345216 699808 364257 699836
rect 270644 699740 273392 699768
rect 270644 699728 270650 699740
rect 273898 699728 273904 699780
rect 273956 699768 273962 699780
rect 283742 699768 283748 699780
rect 273956 699740 283748 699768
rect 273956 699728 273962 699740
rect 283742 699728 283748 699740
rect 283800 699728 283806 699780
rect 283834 699728 283840 699780
rect 283892 699768 283898 699780
rect 288526 699768 288532 699780
rect 283892 699740 288532 699768
rect 283892 699728 283898 699740
rect 288526 699728 288532 699740
rect 288584 699728 288590 699780
rect 296809 699771 296867 699777
rect 296809 699768 296821 699771
rect 288636 699740 296821 699768
rect 171505 699703 171563 699709
rect 171505 699669 171517 699703
rect 171551 699700 171563 699703
rect 186225 699703 186283 699709
rect 186225 699700 186237 699703
rect 171551 699672 186237 699700
rect 171551 699669 171563 699672
rect 171505 699663 171563 699669
rect 186225 699669 186237 699672
rect 186271 699669 186283 699703
rect 186225 699663 186283 699669
rect 249705 699703 249763 699709
rect 249705 699669 249717 699703
rect 249751 699700 249763 699703
rect 251082 699700 251088 699712
rect 249751 699672 251088 699700
rect 249751 699669 249763 699672
rect 249705 699663 249763 699669
rect 251082 699660 251088 699672
rect 251140 699660 251146 699712
rect 267553 699703 267611 699709
rect 267553 699669 267565 699703
rect 267599 699700 267611 699703
rect 269025 699703 269083 699709
rect 269025 699700 269037 699703
rect 267599 699672 269037 699700
rect 267599 699669 267611 699672
rect 267553 699663 267611 699669
rect 269025 699669 269037 699672
rect 269071 699669 269083 699703
rect 269025 699663 269083 699669
rect 269117 699703 269175 699709
rect 269117 699669 269129 699703
rect 269163 699700 269175 699703
rect 273257 699703 273315 699709
rect 273257 699700 273269 699703
rect 269163 699672 273269 699700
rect 269163 699669 269175 699672
rect 269117 699663 269175 699669
rect 273257 699669 273269 699672
rect 273303 699669 273315 699703
rect 273257 699663 273315 699669
rect 273349 699703 273407 699709
rect 273349 699669 273361 699703
rect 273395 699700 273407 699703
rect 282914 699700 282920 699712
rect 273395 699672 282920 699700
rect 273395 699669 273407 699672
rect 273349 699663 273407 699669
rect 282914 699660 282920 699672
rect 282972 699660 282978 699712
rect 283006 699660 283012 699712
rect 283064 699700 283070 699712
rect 288636 699700 288664 699740
rect 296809 699737 296821 699740
rect 296855 699737 296867 699771
rect 296809 699731 296867 699737
rect 296898 699728 296904 699780
rect 296956 699768 296962 699780
rect 311805 699771 311863 699777
rect 311805 699768 311817 699771
rect 296956 699740 311817 699768
rect 296956 699728 296962 699740
rect 311805 699737 311817 699740
rect 311851 699737 311863 699771
rect 311805 699731 311863 699737
rect 331309 699771 331367 699777
rect 331309 699737 331321 699771
rect 331355 699768 331367 699771
rect 340785 699771 340843 699777
rect 340785 699768 340797 699771
rect 331355 699740 340797 699768
rect 331355 699737 331367 699740
rect 331309 699731 331367 699737
rect 340785 699737 340797 699740
rect 340831 699737 340843 699771
rect 340785 699731 340843 699737
rect 344649 699771 344707 699777
rect 344649 699737 344661 699771
rect 344695 699768 344707 699771
rect 345216 699768 345244 699808
rect 364245 699805 364257 699808
rect 364291 699805 364303 699839
rect 364245 699799 364303 699805
rect 344695 699740 345244 699768
rect 344695 699737 344707 699740
rect 344649 699731 344707 699737
rect 283064 699672 288664 699700
rect 283064 699660 283070 699672
rect 288710 699660 288716 699712
rect 288768 699700 288774 699712
rect 292390 699700 292396 699712
rect 288768 699672 292396 699700
rect 288768 699660 288774 699672
rect 292390 699660 292396 699672
rect 292448 699660 292454 699712
rect 292482 699660 292488 699712
rect 292540 699700 292546 699712
rect 302326 699700 302332 699712
rect 292540 699672 302332 699700
rect 292540 699660 292546 699672
rect 302326 699660 302332 699672
rect 302384 699660 302390 699712
rect 302421 699703 302479 699709
rect 302421 699669 302433 699703
rect 302467 699700 302479 699703
rect 311986 699700 311992 699712
rect 302467 699672 311992 699700
rect 302467 699669 302479 699672
rect 302421 699663 302479 699669
rect 311986 699660 311992 699672
rect 312044 699660 312050 699712
rect 316221 699703 316279 699709
rect 316221 699669 316233 699703
rect 316267 699700 316279 699703
rect 326341 699703 326399 699709
rect 326341 699700 326353 699703
rect 316267 699672 326353 699700
rect 316267 699669 316279 699672
rect 316221 699663 316279 699669
rect 326341 699669 326353 699672
rect 326387 699669 326399 699703
rect 326341 699663 326399 699669
rect 335265 699703 335323 699709
rect 335265 699669 335277 699703
rect 335311 699700 335323 699703
rect 345017 699703 345075 699709
rect 345017 699700 345029 699703
rect 335311 699672 345029 699700
rect 335311 699669 335323 699672
rect 335265 699663 335323 699669
rect 345017 699669 345029 699672
rect 345063 699669 345075 699703
rect 345017 699663 345075 699669
rect 345109 699703 345167 699709
rect 345109 699669 345121 699703
rect 345155 699700 345167 699703
rect 354769 699703 354827 699709
rect 354769 699700 354781 699703
rect 345155 699672 354781 699700
rect 345155 699669 345167 699672
rect 345109 699663 345167 699669
rect 354769 699669 354781 699672
rect 354815 699669 354827 699703
rect 354769 699663 354827 699669
rect 364153 699703 364211 699709
rect 364153 699669 364165 699703
rect 364199 699700 364211 699703
rect 364429 699703 364487 699709
rect 364429 699700 364441 699703
rect 364199 699672 364441 699700
rect 364199 699669 364211 699672
rect 364153 699663 364211 699669
rect 364429 699669 364441 699672
rect 364475 699669 364487 699703
rect 364429 699663 364487 699669
rect 373813 699703 373871 699709
rect 373813 699669 373825 699703
rect 373859 699700 373871 699703
rect 374089 699703 374147 699709
rect 374089 699700 374101 699703
rect 373859 699672 374101 699700
rect 373859 699669 373871 699672
rect 373813 699663 373871 699669
rect 374089 699669 374101 699672
rect 374135 699669 374147 699703
rect 374089 699663 374147 699669
rect 383473 699703 383531 699709
rect 383473 699669 383485 699703
rect 383519 699700 383531 699703
rect 383749 699703 383807 699709
rect 383749 699700 383761 699703
rect 383519 699672 383761 699700
rect 383519 699669 383531 699672
rect 383473 699663 383531 699669
rect 383749 699669 383761 699672
rect 383795 699669 383807 699703
rect 383749 699663 383807 699669
rect 1104 699610 582820 699632
rect 1104 699558 36822 699610
rect 36874 699558 36886 699610
rect 36938 699558 36950 699610
rect 37002 699558 37014 699610
rect 37066 699558 37078 699610
rect 37130 699558 37142 699610
rect 37194 699558 37206 699610
rect 37258 699558 37270 699610
rect 37322 699558 37334 699610
rect 37386 699558 72822 699610
rect 72874 699558 72886 699610
rect 72938 699558 72950 699610
rect 73002 699558 73014 699610
rect 73066 699558 73078 699610
rect 73130 699558 73142 699610
rect 73194 699558 73206 699610
rect 73258 699558 73270 699610
rect 73322 699558 73334 699610
rect 73386 699558 108822 699610
rect 108874 699558 108886 699610
rect 108938 699558 108950 699610
rect 109002 699558 109014 699610
rect 109066 699558 109078 699610
rect 109130 699558 109142 699610
rect 109194 699558 109206 699610
rect 109258 699558 109270 699610
rect 109322 699558 109334 699610
rect 109386 699558 144822 699610
rect 144874 699558 144886 699610
rect 144938 699558 144950 699610
rect 145002 699558 145014 699610
rect 145066 699558 145078 699610
rect 145130 699558 145142 699610
rect 145194 699558 145206 699610
rect 145258 699558 145270 699610
rect 145322 699558 145334 699610
rect 145386 699558 180822 699610
rect 180874 699558 180886 699610
rect 180938 699558 180950 699610
rect 181002 699558 181014 699610
rect 181066 699558 181078 699610
rect 181130 699558 181142 699610
rect 181194 699558 181206 699610
rect 181258 699558 181270 699610
rect 181322 699558 181334 699610
rect 181386 699558 216822 699610
rect 216874 699558 216886 699610
rect 216938 699558 216950 699610
rect 217002 699558 217014 699610
rect 217066 699558 217078 699610
rect 217130 699558 217142 699610
rect 217194 699558 217206 699610
rect 217258 699558 217270 699610
rect 217322 699558 217334 699610
rect 217386 699558 252822 699610
rect 252874 699558 252886 699610
rect 252938 699558 252950 699610
rect 253002 699558 253014 699610
rect 253066 699558 253078 699610
rect 253130 699558 253142 699610
rect 253194 699558 253206 699610
rect 253258 699558 253270 699610
rect 253322 699558 253334 699610
rect 253386 699558 288822 699610
rect 288874 699558 288886 699610
rect 288938 699558 288950 699610
rect 289002 699558 289014 699610
rect 289066 699558 289078 699610
rect 289130 699558 289142 699610
rect 289194 699558 289206 699610
rect 289258 699558 289270 699610
rect 289322 699558 289334 699610
rect 289386 699558 324822 699610
rect 324874 699558 324886 699610
rect 324938 699558 324950 699610
rect 325002 699558 325014 699610
rect 325066 699558 325078 699610
rect 325130 699558 325142 699610
rect 325194 699558 325206 699610
rect 325258 699558 325270 699610
rect 325322 699558 325334 699610
rect 325386 699558 360822 699610
rect 360874 699558 360886 699610
rect 360938 699558 360950 699610
rect 361002 699558 361014 699610
rect 361066 699558 361078 699610
rect 361130 699558 361142 699610
rect 361194 699558 361206 699610
rect 361258 699558 361270 699610
rect 361322 699558 361334 699610
rect 361386 699558 396822 699610
rect 396874 699558 396886 699610
rect 396938 699558 396950 699610
rect 397002 699558 397014 699610
rect 397066 699558 397078 699610
rect 397130 699558 397142 699610
rect 397194 699558 397206 699610
rect 397258 699558 397270 699610
rect 397322 699558 397334 699610
rect 397386 699558 432822 699610
rect 432874 699558 432886 699610
rect 432938 699558 432950 699610
rect 433002 699558 433014 699610
rect 433066 699558 433078 699610
rect 433130 699558 433142 699610
rect 433194 699558 433206 699610
rect 433258 699558 433270 699610
rect 433322 699558 433334 699610
rect 433386 699558 468822 699610
rect 468874 699558 468886 699610
rect 468938 699558 468950 699610
rect 469002 699558 469014 699610
rect 469066 699558 469078 699610
rect 469130 699558 469142 699610
rect 469194 699558 469206 699610
rect 469258 699558 469270 699610
rect 469322 699558 469334 699610
rect 469386 699558 504822 699610
rect 504874 699558 504886 699610
rect 504938 699558 504950 699610
rect 505002 699558 505014 699610
rect 505066 699558 505078 699610
rect 505130 699558 505142 699610
rect 505194 699558 505206 699610
rect 505258 699558 505270 699610
rect 505322 699558 505334 699610
rect 505386 699558 540822 699610
rect 540874 699558 540886 699610
rect 540938 699558 540950 699610
rect 541002 699558 541014 699610
rect 541066 699558 541078 699610
rect 541130 699558 541142 699610
rect 541194 699558 541206 699610
rect 541258 699558 541270 699610
rect 541322 699558 541334 699610
rect 541386 699558 576822 699610
rect 576874 699558 576886 699610
rect 576938 699558 576950 699610
rect 577002 699558 577014 699610
rect 577066 699558 577078 699610
rect 577130 699558 577142 699610
rect 577194 699558 577206 699610
rect 577258 699558 577270 699610
rect 577322 699558 577334 699610
rect 577386 699558 582820 699610
rect 1104 699536 582820 699558
rect 142798 699456 142804 699508
rect 142856 699496 142862 699508
rect 403342 699496 403348 699508
rect 142856 699468 403348 699496
rect 142856 699456 142862 699468
rect 403342 699456 403348 699468
rect 403400 699456 403406 699508
rect 71774 699388 71780 699440
rect 71832 699428 71838 699440
rect 354677 699431 354735 699437
rect 354677 699428 354689 699431
rect 71832 699400 354689 699428
rect 71832 699388 71838 699400
rect 354677 699397 354689 699400
rect 354723 699397 354735 699431
rect 354677 699391 354735 699397
rect 354769 699431 354827 699437
rect 354769 699397 354781 699431
rect 354815 699428 354827 699431
rect 364153 699431 364211 699437
rect 364153 699428 364165 699431
rect 354815 699400 364165 699428
rect 354815 699397 354827 699400
rect 354769 699391 354827 699397
rect 364153 699397 364165 699400
rect 364199 699397 364211 699431
rect 364153 699391 364211 699397
rect 364245 699431 364303 699437
rect 364245 699397 364257 699431
rect 364291 699428 364303 699431
rect 417326 699428 417332 699440
rect 364291 699400 417332 699428
rect 364291 699397 364303 699400
rect 364245 699391 364303 699397
rect 417326 699388 417332 699400
rect 417384 699388 417390 699440
rect 100202 699320 100208 699372
rect 100260 699360 100266 699372
rect 273257 699363 273315 699369
rect 273257 699360 273269 699363
rect 100260 699332 273269 699360
rect 100260 699320 100266 699332
rect 273257 699329 273269 699332
rect 273303 699329 273315 699363
rect 273257 699323 273315 699329
rect 273346 699320 273352 699372
rect 273404 699360 273410 699372
rect 282917 699363 282975 699369
rect 282917 699360 282929 699363
rect 273404 699332 282929 699360
rect 273404 699320 273410 699332
rect 282917 699329 282929 699332
rect 282963 699329 282975 699363
rect 282917 699323 282975 699329
rect 283006 699320 283012 699372
rect 283064 699360 283070 699372
rect 296530 699360 296536 699372
rect 283064 699332 296536 699360
rect 283064 699320 283070 699332
rect 296530 699320 296536 699332
rect 296588 699320 296594 699372
rect 296622 699320 296628 699372
rect 296680 699360 296686 699372
rect 383657 699363 383715 699369
rect 383657 699360 383669 699363
rect 296680 699332 383669 699360
rect 296680 699320 296686 699332
rect 383657 699329 383669 699332
rect 383703 699329 383715 699363
rect 383657 699323 383715 699329
rect 383749 699363 383807 699369
rect 383749 699329 383761 699363
rect 383795 699360 383807 699363
rect 445754 699360 445760 699372
rect 383795 699332 445760 699360
rect 383795 699329 383807 699332
rect 383749 699323 383807 699329
rect 445754 699320 445760 699332
rect 445812 699320 445818 699372
rect 133322 699252 133328 699304
rect 133380 699292 133386 699304
rect 146938 699292 146944 699304
rect 133380 699264 146944 699292
rect 133380 699252 133386 699264
rect 146938 699252 146944 699264
rect 146996 699252 147002 699304
rect 161750 699252 161756 699304
rect 161808 699292 161814 699304
rect 579338 699292 579344 699304
rect 161808 699264 579344 699292
rect 161808 699252 161814 699264
rect 579338 699252 579344 699264
rect 579396 699252 579402 699304
rect 48130 699184 48136 699236
rect 48188 699224 48194 699236
rect 142706 699224 142712 699236
rect 48188 699196 142712 699224
rect 48188 699184 48194 699196
rect 142706 699184 142712 699196
rect 142764 699184 142770 699236
rect 147582 699184 147588 699236
rect 147640 699224 147646 699236
rect 186130 699224 186136 699236
rect 147640 699196 186136 699224
rect 147640 699184 147646 699196
rect 186130 699184 186136 699196
rect 186188 699184 186194 699236
rect 186225 699227 186283 699233
rect 186225 699193 186237 699227
rect 186271 699224 186283 699227
rect 267553 699227 267611 699233
rect 267553 699224 267565 699227
rect 186271 699196 267565 699224
rect 186271 699193 186283 699196
rect 186225 699187 186283 699193
rect 267553 699193 267565 699196
rect 267599 699193 267611 699227
rect 267553 699187 267611 699193
rect 267642 699184 267648 699236
rect 267700 699224 267706 699236
rect 302237 699227 302295 699233
rect 302237 699224 302249 699227
rect 267700 699196 302249 699224
rect 267700 699184 267706 699196
rect 302237 699193 302249 699196
rect 302283 699193 302295 699227
rect 302237 699187 302295 699193
rect 302326 699184 302332 699236
rect 302384 699224 302390 699236
rect 305457 699227 305515 699233
rect 302384 699196 305408 699224
rect 302384 699184 302390 699196
rect 5074 699116 5080 699168
rect 5132 699156 5138 699168
rect 303433 699159 303491 699165
rect 303433 699156 303445 699159
rect 5132 699128 303445 699156
rect 5132 699116 5138 699128
rect 303433 699125 303445 699128
rect 303479 699125 303491 699159
rect 303433 699119 303491 699125
rect 303525 699159 303583 699165
rect 303525 699125 303537 699159
rect 303571 699156 303583 699159
rect 305273 699159 305331 699165
rect 305273 699156 305285 699159
rect 303571 699128 305285 699156
rect 303571 699125 303583 699128
rect 303525 699119 303583 699125
rect 305273 699125 305285 699128
rect 305319 699125 305331 699159
rect 305380 699156 305408 699196
rect 305457 699193 305469 699227
rect 305503 699224 305515 699227
rect 311710 699224 311716 699236
rect 305503 699196 311716 699224
rect 305503 699193 305515 699196
rect 305457 699187 305515 699193
rect 311710 699184 311716 699196
rect 311768 699184 311774 699236
rect 311805 699227 311863 699233
rect 311805 699193 311817 699227
rect 311851 699224 311863 699227
rect 344649 699227 344707 699233
rect 344649 699224 344661 699227
rect 311851 699196 344661 699224
rect 311851 699193 311863 699196
rect 311805 699187 311863 699193
rect 344649 699193 344661 699196
rect 344695 699193 344707 699227
rect 344649 699187 344707 699193
rect 344925 699227 344983 699233
rect 344925 699193 344937 699227
rect 344971 699224 344983 699227
rect 364334 699224 364340 699236
rect 344971 699196 364340 699224
rect 344971 699193 344983 699196
rect 344925 699187 344983 699193
rect 364334 699184 364340 699196
rect 364392 699184 364398 699236
rect 364429 699227 364487 699233
rect 364429 699193 364441 699227
rect 364475 699224 364487 699227
rect 373813 699227 373871 699233
rect 373813 699224 373825 699227
rect 364475 699196 373825 699224
rect 364475 699193 364487 699196
rect 364429 699187 364487 699193
rect 373813 699193 373825 699196
rect 373859 699193 373871 699227
rect 373813 699187 373871 699193
rect 373902 699184 373908 699236
rect 373960 699224 373966 699236
rect 373994 699224 374000 699236
rect 373960 699196 374000 699224
rect 373960 699184 373966 699196
rect 373994 699184 374000 699196
rect 374052 699184 374058 699236
rect 374089 699227 374147 699233
rect 374089 699193 374101 699227
rect 374135 699224 374147 699227
rect 383473 699227 383531 699233
rect 383473 699224 383485 699227
rect 374135 699196 383485 699224
rect 374135 699193 374147 699196
rect 374089 699187 374147 699193
rect 383473 699193 383485 699196
rect 383519 699193 383531 699227
rect 383473 699187 383531 699193
rect 383562 699184 383568 699236
rect 383620 699224 383626 699236
rect 579246 699224 579252 699236
rect 383620 699196 579252 699224
rect 383620 699184 383626 699196
rect 579246 699184 579252 699196
rect 579304 699184 579310 699236
rect 321557 699159 321615 699165
rect 321557 699156 321569 699159
rect 305380 699128 321569 699156
rect 305273 699119 305331 699125
rect 321557 699125 321569 699128
rect 321603 699125 321615 699159
rect 321557 699119 321615 699125
rect 321646 699116 321652 699168
rect 321704 699156 321710 699168
rect 331030 699156 331036 699168
rect 321704 699128 331036 699156
rect 321704 699116 321710 699128
rect 331030 699116 331036 699128
rect 331088 699116 331094 699168
rect 331122 699116 331128 699168
rect 331180 699156 331186 699168
rect 336001 699159 336059 699165
rect 336001 699156 336013 699159
rect 331180 699128 336013 699156
rect 331180 699116 331186 699128
rect 336001 699125 336013 699128
rect 336047 699125 336059 699159
rect 336001 699119 336059 699125
rect 336093 699159 336151 699165
rect 336093 699125 336105 699159
rect 336139 699156 336151 699159
rect 340690 699156 340696 699168
rect 336139 699128 340696 699156
rect 336139 699125 336151 699128
rect 336093 699119 336151 699125
rect 340690 699116 340696 699128
rect 340748 699116 340754 699168
rect 340785 699159 340843 699165
rect 340785 699125 340797 699159
rect 340831 699156 340843 699159
rect 344741 699159 344799 699165
rect 344741 699156 344753 699159
rect 340831 699128 344753 699156
rect 340831 699125 340843 699128
rect 340785 699119 340843 699125
rect 344741 699125 344753 699128
rect 344787 699125 344799 699159
rect 344741 699119 344799 699125
rect 344833 699159 344891 699165
rect 344833 699125 344845 699159
rect 344879 699156 344891 699159
rect 459922 699156 459928 699168
rect 344879 699128 459928 699156
rect 344879 699125 344891 699128
rect 344833 699119 344891 699125
rect 459922 699116 459928 699128
rect 459980 699116 459986 699168
rect 1104 699066 582820 699088
rect 1104 699014 18822 699066
rect 18874 699014 18886 699066
rect 18938 699014 18950 699066
rect 19002 699014 19014 699066
rect 19066 699014 19078 699066
rect 19130 699014 19142 699066
rect 19194 699014 19206 699066
rect 19258 699014 19270 699066
rect 19322 699014 19334 699066
rect 19386 699014 54822 699066
rect 54874 699014 54886 699066
rect 54938 699014 54950 699066
rect 55002 699014 55014 699066
rect 55066 699014 55078 699066
rect 55130 699014 55142 699066
rect 55194 699014 55206 699066
rect 55258 699014 55270 699066
rect 55322 699014 55334 699066
rect 55386 699014 90822 699066
rect 90874 699014 90886 699066
rect 90938 699014 90950 699066
rect 91002 699014 91014 699066
rect 91066 699014 91078 699066
rect 91130 699014 91142 699066
rect 91194 699014 91206 699066
rect 91258 699014 91270 699066
rect 91322 699014 91334 699066
rect 91386 699014 126822 699066
rect 126874 699014 126886 699066
rect 126938 699014 126950 699066
rect 127002 699014 127014 699066
rect 127066 699014 127078 699066
rect 127130 699014 127142 699066
rect 127194 699014 127206 699066
rect 127258 699014 127270 699066
rect 127322 699014 127334 699066
rect 127386 699014 162822 699066
rect 162874 699014 162886 699066
rect 162938 699014 162950 699066
rect 163002 699014 163014 699066
rect 163066 699014 163078 699066
rect 163130 699014 163142 699066
rect 163194 699014 163206 699066
rect 163258 699014 163270 699066
rect 163322 699014 163334 699066
rect 163386 699014 198822 699066
rect 198874 699014 198886 699066
rect 198938 699014 198950 699066
rect 199002 699014 199014 699066
rect 199066 699014 199078 699066
rect 199130 699014 199142 699066
rect 199194 699014 199206 699066
rect 199258 699014 199270 699066
rect 199322 699014 199334 699066
rect 199386 699014 234822 699066
rect 234874 699014 234886 699066
rect 234938 699014 234950 699066
rect 235002 699014 235014 699066
rect 235066 699014 235078 699066
rect 235130 699014 235142 699066
rect 235194 699014 235206 699066
rect 235258 699014 235270 699066
rect 235322 699014 235334 699066
rect 235386 699014 270822 699066
rect 270874 699014 270886 699066
rect 270938 699014 270950 699066
rect 271002 699014 271014 699066
rect 271066 699014 271078 699066
rect 271130 699014 271142 699066
rect 271194 699014 271206 699066
rect 271258 699014 271270 699066
rect 271322 699014 271334 699066
rect 271386 699014 306822 699066
rect 306874 699014 306886 699066
rect 306938 699014 306950 699066
rect 307002 699014 307014 699066
rect 307066 699014 307078 699066
rect 307130 699014 307142 699066
rect 307194 699014 307206 699066
rect 307258 699014 307270 699066
rect 307322 699014 307334 699066
rect 307386 699014 342822 699066
rect 342874 699014 342886 699066
rect 342938 699014 342950 699066
rect 343002 699014 343014 699066
rect 343066 699014 343078 699066
rect 343130 699014 343142 699066
rect 343194 699014 343206 699066
rect 343258 699014 343270 699066
rect 343322 699014 343334 699066
rect 343386 699014 378822 699066
rect 378874 699014 378886 699066
rect 378938 699014 378950 699066
rect 379002 699014 379014 699066
rect 379066 699014 379078 699066
rect 379130 699014 379142 699066
rect 379194 699014 379206 699066
rect 379258 699014 379270 699066
rect 379322 699014 379334 699066
rect 379386 699014 414822 699066
rect 414874 699014 414886 699066
rect 414938 699014 414950 699066
rect 415002 699014 415014 699066
rect 415066 699014 415078 699066
rect 415130 699014 415142 699066
rect 415194 699014 415206 699066
rect 415258 699014 415270 699066
rect 415322 699014 415334 699066
rect 415386 699014 450822 699066
rect 450874 699014 450886 699066
rect 450938 699014 450950 699066
rect 451002 699014 451014 699066
rect 451066 699014 451078 699066
rect 451130 699014 451142 699066
rect 451194 699014 451206 699066
rect 451258 699014 451270 699066
rect 451322 699014 451334 699066
rect 451386 699014 486822 699066
rect 486874 699014 486886 699066
rect 486938 699014 486950 699066
rect 487002 699014 487014 699066
rect 487066 699014 487078 699066
rect 487130 699014 487142 699066
rect 487194 699014 487206 699066
rect 487258 699014 487270 699066
rect 487322 699014 487334 699066
rect 487386 699014 522822 699066
rect 522874 699014 522886 699066
rect 522938 699014 522950 699066
rect 523002 699014 523014 699066
rect 523066 699014 523078 699066
rect 523130 699014 523142 699066
rect 523194 699014 523206 699066
rect 523258 699014 523270 699066
rect 523322 699014 523334 699066
rect 523386 699014 558822 699066
rect 558874 699014 558886 699066
rect 558938 699014 558950 699066
rect 559002 699014 559014 699066
rect 559066 699014 559078 699066
rect 559130 699014 559142 699066
rect 559194 699014 559206 699066
rect 559258 699014 559270 699066
rect 559322 699014 559334 699066
rect 559386 699014 582820 699066
rect 1104 698992 582820 699014
rect 119154 698912 119160 698964
rect 119212 698952 119218 698964
rect 244090 698952 244096 698964
rect 119212 698924 244096 698952
rect 119212 698912 119218 698924
rect 244090 698912 244096 698924
rect 244148 698912 244154 698964
rect 244182 698912 244188 698964
rect 244240 698952 244246 698964
rect 244274 698952 244280 698964
rect 244240 698924 244280 698952
rect 244240 698912 244246 698924
rect 244274 698912 244280 698924
rect 244332 698912 244338 698964
rect 244366 698912 244372 698964
rect 244424 698952 244430 698964
rect 253750 698952 253756 698964
rect 244424 698924 253756 698952
rect 244424 698912 244430 698924
rect 253750 698912 253756 698924
rect 253808 698912 253814 698964
rect 253842 698912 253848 698964
rect 253900 698952 253906 698964
rect 282914 698952 282920 698964
rect 253900 698924 282920 698952
rect 253900 698912 253906 698924
rect 282914 698912 282920 698924
rect 282972 698912 282978 698964
rect 283009 698955 283067 698961
rect 283009 698921 283021 698955
rect 283055 698952 283067 698955
rect 303341 698955 303399 698961
rect 303341 698952 303353 698955
rect 283055 698924 303353 698952
rect 283055 698921 283067 698924
rect 283009 698915 283067 698921
rect 303341 698921 303353 698924
rect 303387 698921 303399 698955
rect 303341 698915 303399 698921
rect 303433 698955 303491 698961
rect 303433 698921 303445 698955
rect 303479 698952 303491 698955
rect 321554 698952 321560 698964
rect 303479 698924 321560 698952
rect 303479 698921 303491 698924
rect 303433 698915 303491 698921
rect 321554 698912 321560 698924
rect 321612 698912 321618 698964
rect 321646 698912 321652 698964
rect 321704 698952 321710 698964
rect 335909 698955 335967 698961
rect 335909 698952 335921 698955
rect 321704 698924 335921 698952
rect 321704 698912 321710 698924
rect 335909 698921 335921 698924
rect 335955 698921 335967 698955
rect 335909 698915 335967 698921
rect 336001 698955 336059 698961
rect 336001 698921 336013 698955
rect 336047 698952 336059 698955
rect 344833 698955 344891 698961
rect 344833 698952 344845 698955
rect 336047 698924 344845 698952
rect 336047 698921 336059 698924
rect 336001 698915 336059 698921
rect 344833 698921 344845 698924
rect 344879 698921 344891 698955
rect 344833 698915 344891 698921
rect 344922 698912 344928 698964
rect 344980 698952 344986 698964
rect 579154 698952 579160 698964
rect 344980 698924 579160 698952
rect 344980 698912 344986 698924
rect 579154 698912 579160 698924
rect 579212 698912 579218 698964
rect 57606 698844 57612 698896
rect 57664 698884 57670 698896
rect 107562 698884 107568 698896
rect 57664 698856 107568 698884
rect 57664 698844 57670 698856
rect 107562 698844 107568 698856
rect 107620 698844 107626 698896
rect 114370 698844 114376 698896
rect 114428 698884 114434 698896
rect 577774 698884 577780 698896
rect 114428 698856 577780 698884
rect 114428 698844 114434 698856
rect 577774 698844 577780 698856
rect 577832 698844 577838 698896
rect 5258 698776 5264 698828
rect 5316 698816 5322 698828
rect 474182 698816 474188 698828
rect 5316 698788 474188 698816
rect 5316 698776 5322 698788
rect 474182 698776 474188 698788
rect 474240 698776 474246 698828
rect 33962 698708 33968 698760
rect 34020 698748 34026 698760
rect 89714 698748 89720 698760
rect 34020 698720 89720 698748
rect 34020 698708 34026 698720
rect 89714 698708 89720 698720
rect 89772 698708 89778 698760
rect 104986 698708 104992 698760
rect 105044 698748 105050 698760
rect 579062 698748 579068 698760
rect 105044 698720 579068 698748
rect 105044 698708 105050 698720
rect 579062 698708 579068 698720
rect 579120 698708 579126 698760
rect 90726 698640 90732 698692
rect 90784 698680 90790 698692
rect 578970 698680 578976 698692
rect 90784 698652 578976 698680
rect 90784 698640 90790 698652
rect 578970 698640 578976 698652
rect 579028 698640 579034 698692
rect 5350 698572 5356 698624
rect 5408 698612 5414 698624
rect 502518 698612 502524 698624
rect 5408 698584 502524 698612
rect 5408 698572 5414 698584
rect 502518 698572 502524 698584
rect 502576 698572 502582 698624
rect 1104 698522 582820 698544
rect 1104 698470 36822 698522
rect 36874 698470 36886 698522
rect 36938 698470 36950 698522
rect 37002 698470 37014 698522
rect 37066 698470 37078 698522
rect 37130 698470 37142 698522
rect 37194 698470 37206 698522
rect 37258 698470 37270 698522
rect 37322 698470 37334 698522
rect 37386 698470 72822 698522
rect 72874 698470 72886 698522
rect 72938 698470 72950 698522
rect 73002 698470 73014 698522
rect 73066 698470 73078 698522
rect 73130 698470 73142 698522
rect 73194 698470 73206 698522
rect 73258 698470 73270 698522
rect 73322 698470 73334 698522
rect 73386 698470 108822 698522
rect 108874 698470 108886 698522
rect 108938 698470 108950 698522
rect 109002 698470 109014 698522
rect 109066 698470 109078 698522
rect 109130 698470 109142 698522
rect 109194 698470 109206 698522
rect 109258 698470 109270 698522
rect 109322 698470 109334 698522
rect 109386 698470 144822 698522
rect 144874 698470 144886 698522
rect 144938 698470 144950 698522
rect 145002 698470 145014 698522
rect 145066 698470 145078 698522
rect 145130 698470 145142 698522
rect 145194 698470 145206 698522
rect 145258 698470 145270 698522
rect 145322 698470 145334 698522
rect 145386 698470 180822 698522
rect 180874 698470 180886 698522
rect 180938 698470 180950 698522
rect 181002 698470 181014 698522
rect 181066 698470 181078 698522
rect 181130 698470 181142 698522
rect 181194 698470 181206 698522
rect 181258 698470 181270 698522
rect 181322 698470 181334 698522
rect 181386 698470 216822 698522
rect 216874 698470 216886 698522
rect 216938 698470 216950 698522
rect 217002 698470 217014 698522
rect 217066 698470 217078 698522
rect 217130 698470 217142 698522
rect 217194 698470 217206 698522
rect 217258 698470 217270 698522
rect 217322 698470 217334 698522
rect 217386 698470 252822 698522
rect 252874 698470 252886 698522
rect 252938 698470 252950 698522
rect 253002 698470 253014 698522
rect 253066 698470 253078 698522
rect 253130 698470 253142 698522
rect 253194 698470 253206 698522
rect 253258 698470 253270 698522
rect 253322 698470 253334 698522
rect 253386 698470 288822 698522
rect 288874 698470 288886 698522
rect 288938 698470 288950 698522
rect 289002 698470 289014 698522
rect 289066 698470 289078 698522
rect 289130 698470 289142 698522
rect 289194 698470 289206 698522
rect 289258 698470 289270 698522
rect 289322 698470 289334 698522
rect 289386 698470 324822 698522
rect 324874 698470 324886 698522
rect 324938 698470 324950 698522
rect 325002 698470 325014 698522
rect 325066 698470 325078 698522
rect 325130 698470 325142 698522
rect 325194 698470 325206 698522
rect 325258 698470 325270 698522
rect 325322 698470 325334 698522
rect 325386 698470 360822 698522
rect 360874 698470 360886 698522
rect 360938 698470 360950 698522
rect 361002 698470 361014 698522
rect 361066 698470 361078 698522
rect 361130 698470 361142 698522
rect 361194 698470 361206 698522
rect 361258 698470 361270 698522
rect 361322 698470 361334 698522
rect 361386 698470 396822 698522
rect 396874 698470 396886 698522
rect 396938 698470 396950 698522
rect 397002 698470 397014 698522
rect 397066 698470 397078 698522
rect 397130 698470 397142 698522
rect 397194 698470 397206 698522
rect 397258 698470 397270 698522
rect 397322 698470 397334 698522
rect 397386 698470 432822 698522
rect 432874 698470 432886 698522
rect 432938 698470 432950 698522
rect 433002 698470 433014 698522
rect 433066 698470 433078 698522
rect 433130 698470 433142 698522
rect 433194 698470 433206 698522
rect 433258 698470 433270 698522
rect 433322 698470 433334 698522
rect 433386 698470 468822 698522
rect 468874 698470 468886 698522
rect 468938 698470 468950 698522
rect 469002 698470 469014 698522
rect 469066 698470 469078 698522
rect 469130 698470 469142 698522
rect 469194 698470 469206 698522
rect 469258 698470 469270 698522
rect 469322 698470 469334 698522
rect 469386 698470 504822 698522
rect 504874 698470 504886 698522
rect 504938 698470 504950 698522
rect 505002 698470 505014 698522
rect 505066 698470 505078 698522
rect 505130 698470 505142 698522
rect 505194 698470 505206 698522
rect 505258 698470 505270 698522
rect 505322 698470 505334 698522
rect 505386 698470 540822 698522
rect 540874 698470 540886 698522
rect 540938 698470 540950 698522
rect 541002 698470 541014 698522
rect 541066 698470 541078 698522
rect 541130 698470 541142 698522
rect 541194 698470 541206 698522
rect 541258 698470 541270 698522
rect 541322 698470 541334 698522
rect 541386 698470 576822 698522
rect 576874 698470 576886 698522
rect 576938 698470 576950 698522
rect 577002 698470 577014 698522
rect 577066 698470 577078 698522
rect 577130 698470 577142 698522
rect 577194 698470 577206 698522
rect 577258 698470 577270 698522
rect 577322 698470 577334 698522
rect 577386 698470 582820 698522
rect 1104 698448 582820 698470
rect 76558 698368 76564 698420
rect 76616 698408 76622 698420
rect 218054 698408 218060 698420
rect 76616 698380 218060 698408
rect 76616 698368 76622 698380
rect 218054 698368 218060 698380
rect 218112 698368 218118 698420
rect 218422 698368 218428 698420
rect 218480 698408 218486 698420
rect 237469 698411 237527 698417
rect 237469 698408 237481 698411
rect 218480 698380 237481 698408
rect 218480 698368 218486 698380
rect 237469 698377 237481 698380
rect 237515 698377 237527 698411
rect 237469 698371 237527 698377
rect 237561 698411 237619 698417
rect 237561 698377 237573 698411
rect 237607 698408 237619 698411
rect 578878 698408 578884 698420
rect 237607 698380 578884 698408
rect 237607 698377 237619 698380
rect 237561 698371 237619 698377
rect 578878 698368 578884 698380
rect 578936 698368 578942 698420
rect 62298 698300 62304 698352
rect 62356 698340 62362 698352
rect 218149 698343 218207 698349
rect 218149 698340 218161 698343
rect 62356 698312 218161 698340
rect 62356 698300 62362 698312
rect 218149 698309 218161 698312
rect 218195 698309 218207 698343
rect 218149 698303 218207 698309
rect 218333 698343 218391 698349
rect 218333 698309 218345 698343
rect 218379 698340 218391 698343
rect 237377 698343 237435 698349
rect 237377 698340 237389 698343
rect 218379 698312 237389 698340
rect 218379 698309 218391 698312
rect 218333 698303 218391 698309
rect 237377 698309 237389 698312
rect 237423 698309 237435 698343
rect 237377 698303 237435 698309
rect 237653 698343 237711 698349
rect 237653 698309 237665 698343
rect 237699 698340 237711 698343
rect 577590 698340 577596 698352
rect 237699 698312 577596 698340
rect 237699 698309 237711 698312
rect 237653 698303 237711 698309
rect 577590 698300 577596 698312
rect 577648 698300 577654 698352
rect 5810 698232 5816 698284
rect 5868 698272 5874 698284
rect 218054 698272 218060 698284
rect 5868 698244 218060 698272
rect 5868 698232 5874 698244
rect 218054 698232 218060 698244
rect 218112 698232 218118 698284
rect 218422 698232 218428 698284
rect 218480 698272 218486 698284
rect 237469 698275 237527 698281
rect 237469 698272 237481 698275
rect 218480 698244 237481 698272
rect 218480 698232 218486 698244
rect 237469 698241 237481 698244
rect 237515 698241 237527 698275
rect 237469 698235 237527 698241
rect 237745 698275 237803 698281
rect 237745 698241 237757 698275
rect 237791 698272 237803 698275
rect 237791 698244 350580 698272
rect 237791 698241 237803 698244
rect 237745 698235 237803 698241
rect 5902 698164 5908 698216
rect 5960 698204 5966 698216
rect 136545 698207 136603 698213
rect 5960 698176 30328 698204
rect 5960 698164 5966 698176
rect 30300 698136 30328 698176
rect 107580 698176 129596 698204
rect 107580 698136 107608 698176
rect 30300 698108 107608 698136
rect 129568 698068 129596 698176
rect 136545 698173 136557 698207
rect 136591 698173 136603 698207
rect 153197 698207 153255 698213
rect 153197 698204 153209 698207
rect 136545 698167 136603 698173
rect 144932 698176 153209 698204
rect 136560 698136 136588 698167
rect 144932 698136 144960 698176
rect 153197 698173 153209 698176
rect 153243 698173 153255 698207
rect 153197 698167 153255 698173
rect 186317 698207 186375 698213
rect 186317 698173 186329 698207
rect 186363 698204 186375 698207
rect 215110 698204 215116 698216
rect 186363 698176 193260 698204
rect 215071 698176 215116 698204
rect 186363 698173 186375 698176
rect 186317 698167 186375 698173
rect 193232 698145 193260 698176
rect 215110 698164 215116 698176
rect 215168 698164 215174 698216
rect 215205 698207 215263 698213
rect 215205 698173 215217 698207
rect 215251 698204 215263 698207
rect 218146 698204 218152 698216
rect 215251 698176 218152 698204
rect 215251 698173 215263 698176
rect 215205 698167 215263 698173
rect 218146 698164 218152 698176
rect 218204 698164 218210 698216
rect 218330 698164 218336 698216
rect 218388 698204 218394 698216
rect 226334 698204 226340 698216
rect 218388 698176 226340 698204
rect 218388 698164 218394 698176
rect 226334 698164 226340 698176
rect 226392 698164 226398 698216
rect 235902 698164 235908 698216
rect 235960 698204 235966 698216
rect 237374 698204 237380 698216
rect 235960 698176 237380 698204
rect 235960 698164 235966 698176
rect 237374 698164 237380 698176
rect 237432 698164 237438 698216
rect 237558 698164 237564 698216
rect 237616 698204 237622 698216
rect 253842 698204 253848 698216
rect 237616 698176 253848 698204
rect 237616 698164 237622 698176
rect 253842 698164 253848 698176
rect 253900 698164 253906 698216
rect 254026 698164 254032 698216
rect 254084 698204 254090 698216
rect 350442 698204 350448 698216
rect 254084 698176 350448 698204
rect 254084 698164 254090 698176
rect 350442 698164 350448 698176
rect 350500 698164 350506 698216
rect 350552 698204 350580 698244
rect 350718 698232 350724 698284
rect 350776 698272 350782 698284
rect 365254 698272 365260 698284
rect 350776 698244 365260 698272
rect 350776 698232 350782 698244
rect 365254 698232 365260 698244
rect 365312 698232 365318 698284
rect 383657 698275 383715 698281
rect 383657 698241 383669 698275
rect 383703 698272 383715 698275
rect 393958 698272 393964 698284
rect 383703 698244 393964 698272
rect 383703 698241 383715 698244
rect 383657 698235 383715 698241
rect 393958 698232 393964 698244
rect 394016 698232 394022 698284
rect 351086 698204 351092 698216
rect 350552 698176 351092 698204
rect 351086 698164 351092 698176
rect 351144 698164 351150 698216
rect 354677 698207 354735 698213
rect 354677 698173 354689 698207
rect 354723 698204 354735 698207
rect 580534 698204 580540 698216
rect 354723 698176 580540 698204
rect 354723 698173 354735 698176
rect 354677 698167 354735 698173
rect 580534 698164 580540 698176
rect 580592 698164 580598 698216
rect 136560 698108 144960 698136
rect 157981 698139 158039 698145
rect 157981 698105 157993 698139
rect 158027 698136 158039 698139
rect 172517 698139 172575 698145
rect 172517 698136 172529 698139
rect 158027 698108 165476 698136
rect 158027 698105 158039 698108
rect 157981 698099 158039 698105
rect 136545 698071 136603 698077
rect 136545 698068 136557 698071
rect 129568 698040 136557 698068
rect 136545 698037 136557 698040
rect 136591 698037 136603 698071
rect 165448 698068 165476 698108
rect 169772 698108 172529 698136
rect 169772 698068 169800 698108
rect 172517 698105 172529 698108
rect 172563 698105 172575 698139
rect 172517 698099 172575 698105
rect 182085 698139 182143 698145
rect 182085 698105 182097 698139
rect 182131 698136 182143 698139
rect 186225 698139 186283 698145
rect 186225 698136 186237 698139
rect 182131 698108 186237 698136
rect 182131 698105 182143 698108
rect 182085 698099 182143 698105
rect 186225 698105 186237 698108
rect 186271 698105 186283 698139
rect 186225 698099 186283 698105
rect 193217 698139 193275 698145
rect 193217 698105 193229 698139
rect 193263 698105 193275 698139
rect 193217 698099 193275 698105
rect 193306 698096 193312 698148
rect 193364 698136 193370 698148
rect 193364 698108 193409 698136
rect 193364 698096 193370 698108
rect 202782 698096 202788 698148
rect 202840 698136 202846 698148
rect 208946 698136 208952 698148
rect 202840 698108 208952 698136
rect 202840 698096 202846 698108
rect 208946 698096 208952 698108
rect 209004 698096 209010 698148
rect 209038 698096 209044 698148
rect 209096 698136 209102 698148
rect 218057 698139 218115 698145
rect 218057 698136 218069 698139
rect 209096 698108 218069 698136
rect 209096 698096 209102 698108
rect 218057 698105 218069 698108
rect 218103 698105 218115 698139
rect 218057 698099 218115 698105
rect 218241 698139 218299 698145
rect 218241 698105 218253 698139
rect 218287 698136 218299 698139
rect 237469 698139 237527 698145
rect 237469 698136 237481 698139
rect 218287 698108 237481 698136
rect 218287 698105 218299 698108
rect 218241 698099 218299 698105
rect 237469 698105 237481 698108
rect 237515 698105 237527 698139
rect 237469 698099 237527 698105
rect 237745 698139 237803 698145
rect 237745 698105 237757 698139
rect 237791 698136 237803 698139
rect 576026 698136 576032 698148
rect 237791 698108 576032 698136
rect 237791 698105 237803 698108
rect 237745 698099 237803 698105
rect 576026 698096 576032 698108
rect 576084 698096 576090 698148
rect 165448 698040 169800 698068
rect 136545 698031 136603 698037
rect 213822 698028 213828 698080
rect 213880 698068 213886 698080
rect 237377 698071 237435 698077
rect 237377 698068 237389 698071
rect 213880 698040 237389 698068
rect 213880 698028 213886 698040
rect 237377 698037 237389 698040
rect 237423 698037 237435 698071
rect 237377 698031 237435 698037
rect 237653 698071 237711 698077
rect 237653 698037 237665 698071
rect 237699 698068 237711 698071
rect 579614 698068 579620 698080
rect 237699 698040 579620 698068
rect 237699 698037 237711 698040
rect 237653 698031 237711 698037
rect 579614 698028 579620 698040
rect 579672 698028 579678 698080
rect 1104 697904 6000 698000
rect 6086 697960 6092 698012
rect 6144 698000 6150 698012
rect 379514 698000 379520 698012
rect 6144 697972 379520 698000
rect 6144 697960 6150 697972
rect 379514 697960 379520 697972
rect 379572 697960 379578 698012
rect 153197 697935 153255 697941
rect 153197 697901 153209 697935
rect 153243 697932 153255 697935
rect 157981 697935 158039 697941
rect 157981 697932 157993 697935
rect 153243 697904 157993 697932
rect 153243 697901 153255 697904
rect 153197 697895 153255 697901
rect 157981 697901 157993 697904
rect 158027 697901 158039 697935
rect 157981 697895 158039 697901
rect 172517 697935 172575 697941
rect 172517 697901 172529 697935
rect 172563 697932 172575 697935
rect 182085 697935 182143 697941
rect 182085 697932 182097 697935
rect 172563 697904 182097 697932
rect 172563 697901 172575 697904
rect 172517 697895 172575 697901
rect 182085 697901 182097 697904
rect 182131 697901 182143 697935
rect 182085 697895 182143 697901
rect 194870 697892 194876 697944
rect 194928 697932 194934 697944
rect 574646 697932 574652 697944
rect 194928 697904 574652 697932
rect 194928 697892 194934 697904
rect 574646 697892 574652 697904
rect 574704 697892 574710 697944
rect 578000 697904 582820 698000
rect 6086 697824 6092 697876
rect 6144 697864 6150 697876
rect 393682 697864 393688 697876
rect 6144 697836 393688 697864
rect 6144 697824 6150 697836
rect 393682 697824 393688 697836
rect 393740 697824 393746 697876
rect 393958 697824 393964 697876
rect 394016 697864 394022 697876
rect 580626 697864 580632 697876
rect 394016 697836 580632 697864
rect 394016 697824 394022 697836
rect 580626 697824 580632 697836
rect 580684 697824 580690 697876
rect 7466 697756 7472 697808
rect 7524 697796 7530 697808
rect 398374 697796 398380 697808
rect 7524 697768 398380 697796
rect 7524 697756 7530 697768
rect 398374 697756 398380 697768
rect 398432 697756 398438 697808
rect 180702 697688 180708 697740
rect 180760 697728 180766 697740
rect 575382 697728 575388 697740
rect 180760 697700 575388 697728
rect 180760 697688 180766 697700
rect 575382 697688 575388 697700
rect 575440 697688 575446 697740
rect 6822 697620 6828 697672
rect 6880 697660 6886 697672
rect 407850 697660 407856 697672
rect 6880 697632 407856 697660
rect 6880 697620 6886 697632
rect 407850 697620 407856 697632
rect 407908 697620 407914 697672
rect 166442 697552 166448 697604
rect 166500 697592 166506 697604
rect 575290 697592 575296 697604
rect 166500 697564 575296 697592
rect 166500 697552 166506 697564
rect 575290 697552 575296 697564
rect 575348 697552 575354 697604
rect 6730 697484 6736 697536
rect 6788 697524 6794 697536
rect 422110 697524 422116 697536
rect 6788 697496 422116 697524
rect 6788 697484 6794 697496
rect 422110 697484 422116 697496
rect 422168 697484 422174 697536
rect 1104 697360 6000 697456
rect 152274 697416 152280 697468
rect 152332 697456 152338 697468
rect 575198 697456 575204 697468
rect 152332 697428 575204 697456
rect 152332 697416 152338 697428
rect 575198 697416 575204 697428
rect 575256 697416 575262 697468
rect 6546 697348 6552 697400
rect 6604 697388 6610 697400
rect 436278 697388 436284 697400
rect 6604 697360 436284 697388
rect 6604 697348 6610 697360
rect 436278 697348 436284 697360
rect 436336 697348 436342 697400
rect 578000 697360 582820 697456
rect 6362 697280 6368 697332
rect 6420 697320 6426 697332
rect 455230 697320 455236 697332
rect 6420 697292 455236 697320
rect 6420 697280 6426 697292
rect 455230 697280 455236 697292
rect 455288 697280 455294 697332
rect 6270 697212 6276 697264
rect 6328 697252 6334 697264
rect 464706 697252 464712 697264
rect 6328 697224 464712 697252
rect 6328 697212 6334 697224
rect 464706 697212 464712 697224
rect 464764 697212 464770 697264
rect 7926 697144 7932 697196
rect 7984 697184 7990 697196
rect 493042 697184 493048 697196
rect 7984 697156 493048 697184
rect 7984 697144 7990 697156
rect 493042 697144 493048 697156
rect 493100 697144 493106 697196
rect 7558 697076 7564 697128
rect 7616 697116 7622 697128
rect 535638 697116 535644 697128
rect 7616 697088 535644 697116
rect 7616 697076 7622 697088
rect 535638 697076 535644 697088
rect 535696 697076 535702 697128
rect 38654 697008 38660 697060
rect 38712 697048 38718 697060
rect 574922 697048 574928 697060
rect 38712 697020 574928 697048
rect 38712 697008 38718 697020
rect 574922 697008 574928 697020
rect 574980 697008 574986 697060
rect 24486 696940 24492 696992
rect 24544 696980 24550 696992
rect 574830 696980 574836 696992
rect 24544 696952 574836 696980
rect 24544 696940 24550 696952
rect 574830 696940 574836 696952
rect 574888 696940 574894 696992
rect 19337 696915 19395 696921
rect 1104 696816 6000 696912
rect 19337 696881 19349 696915
rect 19383 696912 19395 696915
rect 28905 696915 28963 696921
rect 28905 696912 28917 696915
rect 19383 696884 28917 696912
rect 19383 696881 19395 696884
rect 19337 696875 19395 696881
rect 28905 696881 28917 696884
rect 28951 696881 28963 696915
rect 28905 696875 28963 696881
rect 165617 696915 165675 696921
rect 165617 696881 165629 696915
rect 165663 696912 165675 696915
rect 175185 696915 175243 696921
rect 175185 696912 175197 696915
rect 165663 696884 175197 696912
rect 165663 696881 165675 696884
rect 165617 696875 165675 696881
rect 175185 696881 175197 696884
rect 175231 696881 175243 696915
rect 175185 696875 175243 696881
rect 224957 696915 225015 696921
rect 224957 696881 224969 696915
rect 225003 696912 225015 696915
rect 232958 696912 232964 696924
rect 225003 696884 232964 696912
rect 225003 696881 225015 696884
rect 224957 696875 225015 696881
rect 232958 696872 232964 696884
rect 233016 696872 233022 696924
rect 233050 696872 233056 696924
rect 233108 696912 233114 696924
rect 248322 696912 248328 696924
rect 233108 696884 248328 696912
rect 233108 696872 233114 696884
rect 248322 696872 248328 696884
rect 248380 696872 248386 696924
rect 248414 696872 248420 696924
rect 248472 696912 248478 696924
rect 253937 696915 253995 696921
rect 253937 696912 253949 696915
rect 248472 696884 253949 696912
rect 248472 696872 248478 696884
rect 253937 696881 253949 696884
rect 253983 696881 253995 696915
rect 253937 696875 253995 696881
rect 263597 696915 263655 696921
rect 263597 696881 263609 696915
rect 263643 696912 263655 696915
rect 271417 696915 271475 696921
rect 271417 696912 271429 696915
rect 263643 696884 271429 696912
rect 263643 696881 263655 696884
rect 263597 696875 263655 696881
rect 271417 696881 271429 696884
rect 271463 696881 271475 696915
rect 277581 696915 277639 696921
rect 271417 696875 271475 696881
rect 274836 696884 275048 696912
rect 6089 696847 6147 696853
rect 6089 696813 6101 696847
rect 6135 696844 6147 696847
rect 274836 696844 274864 696884
rect 6135 696816 274864 696844
rect 275020 696844 275048 696884
rect 277581 696881 277593 696915
rect 277627 696912 277639 696915
rect 284478 696912 284484 696924
rect 277627 696884 284484 696912
rect 277627 696881 277639 696884
rect 277581 696875 277639 696881
rect 284478 696872 284484 696884
rect 284536 696872 284542 696924
rect 284941 696915 284999 696921
rect 284941 696881 284953 696915
rect 284987 696912 284999 696915
rect 289817 696915 289875 696921
rect 289817 696912 289829 696915
rect 284987 696884 289829 696912
rect 284987 696881 284999 696884
rect 284941 696875 284999 696881
rect 289817 696881 289829 696884
rect 289863 696881 289875 696915
rect 289817 696875 289875 696881
rect 302237 696915 302295 696921
rect 302237 696881 302249 696915
rect 302283 696912 302295 696915
rect 311805 696915 311863 696921
rect 311805 696912 311817 696915
rect 302283 696884 311817 696912
rect 302283 696881 302295 696884
rect 302237 696875 302295 696881
rect 311805 696881 311817 696884
rect 311851 696881 311863 696915
rect 311805 696875 311863 696881
rect 321557 696915 321615 696921
rect 321557 696881 321569 696915
rect 321603 696912 321615 696915
rect 331125 696915 331183 696921
rect 331125 696912 331137 696915
rect 321603 696884 331137 696912
rect 321603 696881 321615 696884
rect 321557 696875 321615 696881
rect 331125 696881 331137 696884
rect 331171 696881 331183 696915
rect 331125 696875 331183 696881
rect 340877 696915 340935 696921
rect 340877 696881 340889 696915
rect 340923 696912 340935 696915
rect 350445 696915 350503 696921
rect 350445 696912 350457 696915
rect 340923 696884 350457 696912
rect 340923 696881 340935 696884
rect 340877 696875 340935 696881
rect 350445 696881 350457 696884
rect 350491 696881 350503 696915
rect 360194 696912 360200 696924
rect 350445 696875 350503 696881
rect 350552 696884 360200 696912
rect 289722 696844 289728 696856
rect 275020 696816 289728 696844
rect 6135 696813 6147 696816
rect 6089 696807 6147 696813
rect 289722 696804 289728 696816
rect 289780 696804 289786 696856
rect 309134 696844 309140 696856
rect 309060 696816 309140 696844
rect 309060 696788 309088 696816
rect 309134 696804 309140 696816
rect 309192 696804 309198 696856
rect 19337 696779 19395 696785
rect 19337 696776 19349 696779
rect 15856 696748 19349 696776
rect 4062 696668 4068 696720
rect 4120 696708 4126 696720
rect 6089 696711 6147 696717
rect 6089 696708 6101 696711
rect 4120 696680 6101 696708
rect 4120 696668 4126 696680
rect 6089 696677 6101 696680
rect 6135 696677 6147 696711
rect 15856 696708 15884 696748
rect 19337 696745 19349 696748
rect 19383 696745 19395 696779
rect 128357 696779 128415 696785
rect 19337 696739 19395 696745
rect 89640 696748 98500 696776
rect 6089 696671 6147 696677
rect 10336 696680 15884 696708
rect 28905 696711 28963 696717
rect 5442 696600 5448 696652
rect 5500 696640 5506 696652
rect 10336 696640 10364 696680
rect 28905 696677 28917 696711
rect 28951 696708 28963 696711
rect 89640 696708 89668 696748
rect 28951 696680 89668 696708
rect 98472 696708 98500 696748
rect 128357 696745 128369 696779
rect 128403 696776 128415 696779
rect 160094 696776 160100 696788
rect 128403 696748 160100 696776
rect 128403 696745 128415 696748
rect 128357 696739 128415 696745
rect 160094 696736 160100 696748
rect 160152 696736 160158 696788
rect 160186 696736 160192 696788
rect 160244 696776 160250 696788
rect 165617 696779 165675 696785
rect 165617 696776 165629 696779
rect 160244 696748 165629 696776
rect 160244 696736 160250 696748
rect 165617 696745 165629 696748
rect 165663 696745 165675 696779
rect 207017 696779 207075 696785
rect 207017 696776 207029 696779
rect 165617 696739 165675 696745
rect 199948 696748 207029 696776
rect 128265 696711 128323 696717
rect 128265 696708 128277 696711
rect 98472 696680 128277 696708
rect 28951 696677 28963 696680
rect 28905 696671 28963 696677
rect 128265 696677 128277 696680
rect 128311 696677 128323 696711
rect 128265 696671 128323 696677
rect 175185 696711 175243 696717
rect 175185 696677 175197 696711
rect 175231 696708 175243 696711
rect 199948 696708 199976 696748
rect 207017 696745 207029 696748
rect 207063 696745 207075 696779
rect 224957 696779 225015 696785
rect 224957 696776 224969 696779
rect 207017 696739 207075 696745
rect 218440 696748 224969 696776
rect 175231 696680 199976 696708
rect 207109 696711 207167 696717
rect 175231 696677 175243 696680
rect 175185 696671 175243 696677
rect 207109 696677 207121 696711
rect 207155 696708 207167 696711
rect 218440 696708 218468 696748
rect 224957 696745 224969 696748
rect 225003 696745 225015 696779
rect 224957 696739 225015 696745
rect 234522 696736 234528 696788
rect 234580 696776 234586 696788
rect 244274 696776 244280 696788
rect 234580 696748 244280 696776
rect 234580 696736 234586 696748
rect 244274 696736 244280 696748
rect 244332 696736 244338 696788
rect 253937 696779 253995 696785
rect 253937 696745 253949 696779
rect 253983 696776 253995 696779
rect 263597 696779 263655 696785
rect 263597 696776 263609 696779
rect 253983 696748 263609 696776
rect 253983 696745 253995 696748
rect 253937 696739 253995 696745
rect 263597 696745 263609 696748
rect 263643 696745 263655 696779
rect 263597 696739 263655 696745
rect 271417 696779 271475 696785
rect 271417 696745 271429 696779
rect 271463 696776 271475 696779
rect 284941 696779 284999 696785
rect 284941 696776 284953 696779
rect 271463 696748 284953 696776
rect 271463 696745 271475 696748
rect 271417 696739 271475 696745
rect 284941 696745 284953 696748
rect 284987 696745 284999 696779
rect 284941 696739 284999 696745
rect 289817 696779 289875 696785
rect 289817 696745 289829 696779
rect 289863 696776 289875 696779
rect 299474 696776 299480 696788
rect 289863 696748 299480 696776
rect 289863 696745 289875 696748
rect 289817 696739 289875 696745
rect 299474 696736 299480 696748
rect 299532 696736 299538 696788
rect 309042 696736 309048 696788
rect 309100 696736 309106 696788
rect 321554 696736 321560 696788
rect 321612 696776 321618 696788
rect 328454 696776 328460 696788
rect 321612 696748 328460 696776
rect 321612 696736 321618 696748
rect 328454 696736 328460 696748
rect 328512 696736 328518 696788
rect 342622 696736 342628 696788
rect 342680 696776 342686 696788
rect 350552 696776 350580 696884
rect 360194 696872 360200 696884
rect 360252 696872 360258 696924
rect 355321 696847 355379 696853
rect 355321 696813 355333 696847
rect 355367 696844 355379 696847
rect 364981 696847 365039 696853
rect 364981 696844 364993 696847
rect 355367 696816 364993 696844
rect 355367 696813 355379 696816
rect 355321 696807 355379 696813
rect 364981 696813 364993 696816
rect 365027 696813 365039 696847
rect 578000 696816 582820 696912
rect 364981 696807 365039 696813
rect 342680 696748 350580 696776
rect 371145 696779 371203 696785
rect 342680 696736 342686 696748
rect 371145 696745 371157 696779
rect 371191 696776 371203 696779
rect 388990 696776 388996 696788
rect 371191 696748 388996 696776
rect 371191 696745 371203 696748
rect 371145 696739 371203 696745
rect 388990 696736 388996 696748
rect 389048 696736 389054 696788
rect 207155 696680 218468 696708
rect 207155 696677 207167 696680
rect 207109 696671 207167 696677
rect 218514 696668 218520 696720
rect 218572 696708 218578 696720
rect 578694 696708 578700 696720
rect 218572 696680 578700 696708
rect 218572 696668 218578 696680
rect 578694 696668 578700 696680
rect 578752 696668 578758 696720
rect 5500 696612 10364 696640
rect 5500 696600 5506 696612
rect 146938 696600 146944 696652
rect 146996 696640 147002 696652
rect 208489 696643 208547 696649
rect 208489 696640 208501 696643
rect 146996 696612 208501 696640
rect 146996 696600 147002 696612
rect 208489 696609 208501 696612
rect 208535 696609 208547 696643
rect 208489 696603 208547 696609
rect 208673 696643 208731 696649
rect 208673 696609 208685 696643
rect 208719 696640 208731 696643
rect 580718 696640 580724 696652
rect 208719 696612 580724 696640
rect 208719 696609 208731 696612
rect 208673 696603 208731 696609
rect 580718 696600 580724 696612
rect 580776 696600 580782 696652
rect 113085 696575 113143 696581
rect 113085 696541 113097 696575
rect 113131 696572 113143 696575
rect 116581 696575 116639 696581
rect 116581 696572 116593 696575
rect 113131 696544 116593 696572
rect 113131 696541 113143 696544
rect 113085 696535 113143 696541
rect 116581 696541 116593 696544
rect 116627 696541 116639 696575
rect 116581 696535 116639 696541
rect 142706 696532 142712 696584
rect 142764 696572 142770 696584
rect 208397 696575 208455 696581
rect 208397 696572 208409 696575
rect 142764 696544 208409 696572
rect 142764 696532 142770 696544
rect 208397 696541 208409 696544
rect 208443 696541 208455 696575
rect 208397 696535 208455 696541
rect 208765 696575 208823 696581
rect 208765 696541 208777 696575
rect 208811 696572 208823 696575
rect 580350 696572 580356 696584
rect 208811 696544 580356 696572
rect 208811 696541 208823 696544
rect 208765 696535 208823 696541
rect 580350 696532 580356 696544
rect 580408 696532 580414 696584
rect 3142 696464 3148 696516
rect 3200 696504 3206 696516
rect 374730 696504 374736 696516
rect 3200 696476 374736 696504
rect 3200 696464 3206 696476
rect 374730 696464 374736 696476
rect 374788 696464 374794 696516
rect 403342 696464 403348 696516
rect 403400 696504 403406 696516
rect 580810 696504 580816 696516
rect 403400 696476 580816 696504
rect 403400 696464 403406 696476
rect 580810 696464 580816 696476
rect 580868 696464 580874 696516
rect 113085 696439 113143 696445
rect 113085 696436 113097 696439
rect 30300 696408 113097 696436
rect 30300 696368 30328 696408
rect 113085 696405 113097 696408
rect 113131 696405 113143 696439
rect 113085 696399 113143 696405
rect 116581 696439 116639 696445
rect 116581 696405 116593 696439
rect 116627 696436 116639 696439
rect 143721 696439 143779 696445
rect 116627 696408 131252 696436
rect 116627 696405 116639 696408
rect 116581 696399 116639 696405
rect 1104 696272 6000 696368
rect 8036 696340 30328 696368
rect 3878 696192 3884 696244
rect 3936 696232 3942 696244
rect 8036 696232 8064 696340
rect 131224 696300 131252 696408
rect 143721 696405 143733 696439
rect 143767 696436 143779 696439
rect 160097 696439 160155 696445
rect 143767 696408 149100 696436
rect 143767 696405 143779 696408
rect 143721 696399 143779 696405
rect 149072 696368 149100 696408
rect 160097 696405 160109 696439
rect 160143 696436 160155 696439
rect 165522 696436 165528 696448
rect 160143 696408 165528 696436
rect 160143 696405 160155 696408
rect 160097 696399 160155 696405
rect 165522 696396 165528 696408
rect 165580 696396 165586 696448
rect 165706 696396 165712 696448
rect 165764 696436 165770 696448
rect 165764 696408 200804 696436
rect 165764 696396 165770 696408
rect 160005 696371 160063 696377
rect 160005 696368 160017 696371
rect 149072 696340 160017 696368
rect 160005 696337 160017 696340
rect 160051 696337 160063 696371
rect 200776 696368 200804 696408
rect 204346 696396 204352 696448
rect 204404 696436 204410 696448
rect 578786 696436 578792 696448
rect 204404 696408 578792 696436
rect 204404 696396 204410 696408
rect 578786 696396 578792 696408
rect 578844 696396 578850 696448
rect 205637 696371 205695 696377
rect 205637 696368 205649 696371
rect 200776 696340 205649 696368
rect 160005 696331 160063 696337
rect 205637 696337 205649 696340
rect 205683 696337 205695 696371
rect 205637 696331 205695 696337
rect 205729 696371 205787 696377
rect 205729 696337 205741 696371
rect 205775 696368 205787 696371
rect 224954 696368 224960 696380
rect 205775 696340 224960 696368
rect 205775 696337 205787 696340
rect 205729 696331 205787 696337
rect 224954 696328 224960 696340
rect 225012 696328 225018 696380
rect 234522 696328 234528 696380
rect 234580 696368 234586 696380
rect 244274 696368 244280 696380
rect 234580 696340 244280 696368
rect 234580 696328 234586 696340
rect 244274 696328 244280 696340
rect 244332 696328 244338 696380
rect 253842 696328 253848 696380
rect 253900 696368 253906 696380
rect 263594 696368 263600 696380
rect 253900 696340 263600 696368
rect 253900 696328 253906 696340
rect 263594 696328 263600 696340
rect 263652 696328 263658 696380
rect 273162 696328 273168 696380
rect 273220 696368 273226 696380
rect 282914 696368 282920 696380
rect 273220 696340 282920 696368
rect 273220 696328 273226 696340
rect 282914 696328 282920 696340
rect 282972 696328 282978 696380
rect 292482 696328 292488 696380
rect 292540 696368 292546 696380
rect 302237 696371 302295 696377
rect 302237 696368 302249 696371
rect 292540 696340 302249 696368
rect 292540 696328 292546 696340
rect 302237 696337 302249 696340
rect 302283 696337 302295 696371
rect 302237 696331 302295 696337
rect 311805 696371 311863 696377
rect 311805 696337 311817 696371
rect 311851 696368 311863 696371
rect 321557 696371 321615 696377
rect 321557 696368 321569 696371
rect 311851 696340 321569 696368
rect 311851 696337 311863 696340
rect 311805 696331 311863 696337
rect 321557 696337 321569 696340
rect 321603 696337 321615 696371
rect 321557 696331 321615 696337
rect 331125 696371 331183 696377
rect 331125 696337 331137 696371
rect 331171 696368 331183 696371
rect 340877 696371 340935 696377
rect 340877 696368 340889 696371
rect 331171 696340 340889 696368
rect 331171 696337 331183 696340
rect 331125 696331 331183 696337
rect 340877 696337 340889 696340
rect 340923 696337 340935 696371
rect 340877 696331 340935 696337
rect 350445 696371 350503 696377
rect 350445 696337 350457 696371
rect 350491 696368 350503 696371
rect 355321 696371 355379 696377
rect 355321 696368 355333 696371
rect 350491 696340 355333 696368
rect 350491 696337 350503 696340
rect 350445 696331 350503 696337
rect 355321 696337 355333 696340
rect 355367 696337 355379 696371
rect 355321 696331 355379 696337
rect 364981 696371 365039 696377
rect 364981 696337 364993 696371
rect 365027 696368 365039 696371
rect 371145 696371 371203 696377
rect 371145 696368 371157 696371
rect 365027 696340 371157 696368
rect 365027 696337 365039 696340
rect 364981 696331 365039 696337
rect 371145 696337 371157 696340
rect 371191 696337 371203 696371
rect 371145 696331 371203 696337
rect 143721 696303 143779 696309
rect 143721 696300 143733 696303
rect 131224 696272 143733 696300
rect 143721 696269 143733 696272
rect 143767 696269 143779 696303
rect 143721 696263 143779 696269
rect 190178 696260 190184 696312
rect 190236 696300 190242 696312
rect 563425 696303 563483 696309
rect 563425 696300 563437 696303
rect 190236 696272 563437 696300
rect 190236 696260 190242 696272
rect 563425 696269 563437 696272
rect 563471 696269 563483 696303
rect 578000 696272 582820 696368
rect 563425 696263 563483 696269
rect 81250 696232 81256 696244
rect 3936 696204 8064 696232
rect 81211 696204 81256 696232
rect 3936 696192 3942 696204
rect 81250 696192 81256 696204
rect 81308 696192 81314 696244
rect 107562 696192 107568 696244
rect 107620 696232 107626 696244
rect 580442 696232 580448 696244
rect 107620 696204 580448 696232
rect 107620 696192 107626 696204
rect 580442 696192 580448 696204
rect 580500 696192 580506 696244
rect 3326 696124 3332 696176
rect 3384 696164 3390 696176
rect 403158 696164 403164 696176
rect 3384 696136 403164 696164
rect 3384 696124 3390 696136
rect 403158 696124 403164 696136
rect 403216 696124 403222 696176
rect 563425 696167 563483 696173
rect 563425 696133 563437 696167
rect 563471 696164 563483 696167
rect 579522 696164 579528 696176
rect 563471 696136 579528 696164
rect 563471 696133 563483 696136
rect 563425 696127 563483 696133
rect 579522 696124 579528 696136
rect 579580 696124 579586 696176
rect 8202 696056 8208 696108
rect 8260 696096 8266 696108
rect 412634 696096 412640 696108
rect 8260 696068 412640 696096
rect 8260 696056 8266 696068
rect 412634 696056 412640 696068
rect 412692 696056 412698 696108
rect 425146 696056 425152 696108
rect 425204 696096 425210 696108
rect 426894 696096 426900 696108
rect 425204 696068 426900 696096
rect 425204 696056 425210 696068
rect 426894 696056 426900 696068
rect 426952 696056 426958 696108
rect 5166 695988 5172 696040
rect 5224 696028 5230 696040
rect 431310 696028 431316 696040
rect 5224 696000 431316 696028
rect 5224 695988 5230 696000
rect 431310 695988 431316 696000
rect 431368 695988 431374 696040
rect 6454 695920 6460 695972
rect 6512 695960 6518 695972
rect 450078 695960 450084 695972
rect 6512 695932 450084 695960
rect 6512 695920 6518 695932
rect 450078 695920 450084 695932
rect 450136 695920 450142 695972
rect 3786 695852 3792 695904
rect 3844 695892 3850 695904
rect 469214 695892 469220 695904
rect 3844 695864 469220 695892
rect 3844 695852 3850 695864
rect 469214 695852 469220 695864
rect 469272 695852 469278 695904
rect 1104 695728 6000 695824
rect 8018 695784 8024 695836
rect 8076 695824 8082 695836
rect 478782 695824 478788 695836
rect 8076 695796 478788 695824
rect 8076 695784 8082 695796
rect 478782 695784 478788 695796
rect 478840 695784 478846 695836
rect 485774 695784 485780 695836
rect 485832 695824 485838 695836
rect 492582 695824 492588 695836
rect 485832 695796 492588 695824
rect 485832 695784 485838 695796
rect 492582 695784 492588 695796
rect 492640 695784 492646 695836
rect 487982 695756 487988 695768
rect 6104 695728 487988 695756
rect 4890 695648 4896 695700
rect 4948 695688 4954 695700
rect 6104 695688 6132 695728
rect 487982 695716 487988 695728
rect 488040 695716 488046 695768
rect 562318 695716 562324 695768
rect 562376 695756 562382 695768
rect 567102 695756 567108 695768
rect 562376 695728 567108 695756
rect 562376 695716 562382 695728
rect 567102 695716 567108 695728
rect 567160 695716 567166 695768
rect 578000 695728 582820 695824
rect 4948 695660 6132 695688
rect 4948 695648 4954 695660
rect 7742 695648 7748 695700
rect 7800 695688 7806 695700
rect 506934 695688 506940 695700
rect 7800 695660 506940 695688
rect 7800 695648 7806 695660
rect 506934 695648 506940 695660
rect 506992 695648 506998 695700
rect 540974 695648 540980 695700
rect 541032 695688 541038 695700
rect 543826 695688 543832 695700
rect 541032 695660 543832 695688
rect 541032 695648 541038 695660
rect 543826 695648 543832 695660
rect 543884 695648 543890 695700
rect 53282 695580 53288 695632
rect 53340 695620 53346 695632
rect 575014 695620 575020 695632
rect 53340 695592 575020 695620
rect 53340 695580 53346 695592
rect 575014 695580 575020 695592
rect 575072 695580 575078 695632
rect 3510 695512 3516 695564
rect 3568 695552 3574 695564
rect 530670 695552 530676 695564
rect 3568 695524 530676 695552
rect 3568 695512 3574 695524
rect 530670 695512 530676 695524
rect 530728 695512 530734 695564
rect 7282 695444 7288 695496
rect 7340 695484 7346 695496
rect 355502 695484 355508 695496
rect 7340 695456 355508 695484
rect 7340 695444 7346 695456
rect 355502 695444 355508 695456
rect 355560 695444 355566 695496
rect 355597 695487 355655 695493
rect 355597 695453 355609 695487
rect 355643 695484 355655 695487
rect 364981 695487 365039 695493
rect 364981 695484 364993 695487
rect 355643 695456 364993 695484
rect 355643 695453 355655 695456
rect 355597 695447 355655 695453
rect 364981 695453 364993 695456
rect 365027 695453 365039 695487
rect 364981 695447 365039 695453
rect 375374 695444 375380 695496
rect 375432 695484 375438 695496
rect 384942 695484 384948 695496
rect 375432 695456 384948 695484
rect 375432 695444 375438 695456
rect 384942 695444 384948 695456
rect 385000 695444 385006 695496
rect 7374 695376 7380 695428
rect 7432 695416 7438 695428
rect 369946 695416 369952 695428
rect 7432 695388 369952 695416
rect 7432 695376 7438 695388
rect 369946 695376 369952 695388
rect 370004 695376 370010 695428
rect 374641 695419 374699 695425
rect 374641 695385 374653 695419
rect 374687 695416 374699 695419
rect 384301 695419 384359 695425
rect 384301 695416 384313 695419
rect 374687 695388 384313 695416
rect 374687 695385 374699 695388
rect 374641 695379 374699 695385
rect 384301 695385 384313 695388
rect 384347 695385 384359 695419
rect 384301 695379 384359 695385
rect 432601 695419 432659 695425
rect 432601 695385 432613 695419
rect 432647 695416 432659 695419
rect 442261 695419 442319 695425
rect 442261 695416 442273 695419
rect 432647 695388 442273 695416
rect 432647 695385 432659 695388
rect 432601 695379 432659 695385
rect 442261 695385 442273 695388
rect 442307 695385 442319 695419
rect 442261 695379 442319 695385
rect 3234 695308 3240 695360
rect 3292 695348 3298 695360
rect 383838 695348 383844 695360
rect 3292 695320 383844 695348
rect 3292 695308 3298 695320
rect 383838 695308 383844 695320
rect 383896 695308 383902 695360
rect 393961 695351 394019 695357
rect 393961 695317 393973 695351
rect 394007 695348 394019 695351
rect 403621 695351 403679 695357
rect 403621 695348 403633 695351
rect 394007 695320 403633 695348
rect 394007 695317 394019 695320
rect 393961 695311 394019 695317
rect 403621 695317 403633 695320
rect 403667 695317 403679 695351
rect 403621 695311 403679 695317
rect 413281 695351 413339 695357
rect 413281 695317 413293 695351
rect 413327 695348 413339 695351
rect 422941 695351 422999 695357
rect 422941 695348 422953 695351
rect 413327 695320 422953 695348
rect 413327 695317 413339 695320
rect 413281 695311 413339 695317
rect 422941 695317 422953 695320
rect 422987 695317 422999 695351
rect 440694 695348 440700 695360
rect 440655 695320 440700 695348
rect 422941 695311 422999 695317
rect 440694 695308 440700 695320
rect 440752 695308 440758 695360
rect 483382 695348 483388 695360
rect 483343 695320 483388 695348
rect 483382 695308 483388 695320
rect 483440 695308 483446 695360
rect 497550 695348 497556 695360
rect 497511 695320 497556 695348
rect 497550 695308 497556 695320
rect 497608 695308 497614 695360
rect 511902 695348 511908 695360
rect 511863 695320 511908 695348
rect 511902 695308 511908 695320
rect 511960 695308 511966 695360
rect 578142 695348 578148 695360
rect 577516 695320 578148 695348
rect 29546 695280 29552 695292
rect 1104 695184 6000 695280
rect 29507 695252 29552 695280
rect 29546 695240 29552 695252
rect 29604 695240 29610 695292
rect 43714 695280 43720 695292
rect 43675 695252 43720 695280
rect 43714 695240 43720 695252
rect 43772 695240 43778 695292
rect 67450 695280 67456 695292
rect 67411 695252 67456 695280
rect 67450 695240 67456 695252
rect 67508 695240 67514 695292
rect 86402 695280 86408 695292
rect 86363 695252 86408 695280
rect 86402 695240 86408 695252
rect 86460 695240 86466 695292
rect 95786 695280 95792 695292
rect 95747 695252 95792 695280
rect 95786 695240 95792 695252
rect 95844 695240 95850 695292
rect 109954 695280 109960 695292
rect 109915 695252 109960 695280
rect 109954 695240 109960 695252
rect 110012 695240 110018 695292
rect 124122 695280 124128 695292
rect 124083 695252 124128 695280
rect 124122 695240 124128 695252
rect 124180 695240 124186 695292
rect 128906 695280 128912 695292
rect 128867 695252 128912 695280
rect 128906 695240 128912 695252
rect 128964 695240 128970 695292
rect 138474 695280 138480 695292
rect 138435 695252 138480 695280
rect 138474 695240 138480 695252
rect 138532 695240 138538 695292
rect 140593 695283 140651 695289
rect 140593 695249 140605 695283
rect 140639 695280 140651 695283
rect 152461 695283 152519 695289
rect 152461 695280 152473 695283
rect 140639 695252 152473 695280
rect 140639 695249 140651 695252
rect 140593 695243 140651 695249
rect 152461 695249 152473 695252
rect 152507 695249 152519 695283
rect 152461 695243 152519 695249
rect 171594 695240 171600 695292
rect 171652 695240 171658 695292
rect 185762 695240 185768 695292
rect 185820 695240 185826 695292
rect 199930 695240 199936 695292
rect 199988 695280 199994 695292
rect 577406 695280 577412 695292
rect 199988 695252 577412 695280
rect 199988 695240 199994 695252
rect 577406 695240 577412 695252
rect 577464 695240 577470 695292
rect 14001 695215 14059 695221
rect 14001 695181 14013 695215
rect 14047 695212 14059 695215
rect 103425 695215 103483 695221
rect 103425 695212 103437 695215
rect 14047 695184 103437 695212
rect 14047 695181 14059 695184
rect 14001 695175 14059 695181
rect 103425 695181 103437 695184
rect 103471 695181 103483 695215
rect 144917 695215 144975 695221
rect 144917 695212 144929 695215
rect 103425 695175 103483 695181
rect 120092 695184 144929 695212
rect 103517 695147 103575 695153
rect 103517 695113 103529 695147
rect 103563 695144 103575 695147
rect 120092 695144 120120 695184
rect 144917 695181 144929 695184
rect 144963 695181 144975 695215
rect 144917 695175 144975 695181
rect 145009 695215 145067 695221
rect 145009 695181 145021 695215
rect 145055 695212 145067 695215
rect 164329 695215 164387 695221
rect 145055 695184 164280 695212
rect 145055 695181 145067 695184
rect 145009 695175 145067 695181
rect 164252 695153 164280 695184
rect 164329 695181 164341 695215
rect 164375 695212 164387 695215
rect 171505 695215 171563 695221
rect 171505 695212 171517 695215
rect 164375 695184 171517 695212
rect 164375 695181 164387 695184
rect 164329 695175 164387 695181
rect 171505 695181 171517 695184
rect 171551 695181 171563 695215
rect 171505 695175 171563 695181
rect 103563 695116 120120 695144
rect 164237 695147 164295 695153
rect 103563 695113 103575 695116
rect 103517 695107 103575 695113
rect 164237 695113 164249 695147
rect 164283 695113 164295 695147
rect 171612 695144 171640 695240
rect 185780 695212 185808 695240
rect 577516 695212 577544 695320
rect 578142 695308 578148 695320
rect 578200 695308 578206 695360
rect 185780 695184 577544 695212
rect 578000 695184 582820 695280
rect 578050 695144 578056 695156
rect 171612 695116 578056 695144
rect 164237 695107 164295 695113
rect 578050 695104 578056 695116
rect 578108 695104 578114 695156
rect 3970 695036 3976 695088
rect 4028 695076 4034 695088
rect 8021 695079 8079 695085
rect 8021 695076 8033 695079
rect 4028 695048 8033 695076
rect 4028 695036 4034 695048
rect 8021 695045 8033 695048
rect 8067 695045 8079 695079
rect 8021 695039 8079 695045
rect 8110 695036 8116 695088
rect 8168 695076 8174 695088
rect 15013 695079 15071 695085
rect 15013 695076 15025 695079
rect 8168 695048 15025 695076
rect 8168 695036 8174 695048
rect 15013 695045 15025 695048
rect 15059 695045 15071 695079
rect 15013 695039 15071 695045
rect 15197 695079 15255 695085
rect 15197 695045 15209 695079
rect 15243 695076 15255 695079
rect 440697 695079 440755 695085
rect 440697 695076 440709 695079
rect 15243 695048 440709 695076
rect 15243 695045 15255 695048
rect 15197 695039 15255 695045
rect 440697 695045 440709 695048
rect 440743 695045 440755 695079
rect 440697 695039 440755 695045
rect 450265 695079 450323 695085
rect 450265 695045 450277 695079
rect 450311 695076 450323 695079
rect 459925 695079 459983 695085
rect 459925 695076 459937 695079
rect 450311 695048 459937 695076
rect 450311 695045 450323 695048
rect 450265 695039 450323 695045
rect 459925 695045 459937 695048
rect 459971 695045 459983 695079
rect 459925 695039 459983 695045
rect 469585 695079 469643 695085
rect 469585 695045 469597 695079
rect 469631 695076 469643 695079
rect 483385 695079 483443 695085
rect 483385 695076 483397 695079
rect 469631 695048 483397 695076
rect 469631 695045 469643 695048
rect 469585 695039 469643 695045
rect 483385 695045 483397 695048
rect 483431 695045 483443 695079
rect 483385 695039 483443 695045
rect 138477 695011 138535 695017
rect 138477 694977 138489 695011
rect 138523 695008 138535 695011
rect 576762 695008 576768 695020
rect 138523 694980 576768 695008
rect 138523 694977 138535 694980
rect 138477 694971 138535 694977
rect 576762 694968 576768 694980
rect 576820 694968 576826 695020
rect 8021 694943 8079 694949
rect 8021 694909 8033 694943
rect 8067 694940 8079 694943
rect 14001 694943 14059 694949
rect 14001 694940 14013 694943
rect 8067 694912 14013 694940
rect 8067 694909 8079 694912
rect 8021 694903 8079 694909
rect 14001 694909 14013 694912
rect 14047 694909 14059 694943
rect 125597 694943 125655 694949
rect 125597 694940 125609 694943
rect 14001 694903 14059 694909
rect 123496 694912 125609 694940
rect 123496 694872 123524 694912
rect 125597 694909 125609 694912
rect 125643 694909 125655 694943
rect 125597 694903 125655 694909
rect 128909 694943 128967 694949
rect 128909 694909 128921 694943
rect 128955 694940 128967 694943
rect 577866 694940 577872 694952
rect 128955 694912 577872 694940
rect 128955 694909 128967 694912
rect 128909 694903 128967 694909
rect 577866 694900 577872 694912
rect 577924 694900 577930 694952
rect 108316 694844 123524 694872
rect 124125 694875 124183 694881
rect 108316 694804 108344 694844
rect 124125 694841 124137 694875
rect 124171 694872 124183 694875
rect 576670 694872 576676 694884
rect 124171 694844 576676 694872
rect 124171 694841 124183 694844
rect 124125 694835 124183 694841
rect 576670 694832 576676 694844
rect 576728 694832 576734 694884
rect 22112 694776 108344 694804
rect 109957 694807 110015 694813
rect 22112 694736 22140 694776
rect 109957 694773 109969 694807
rect 110003 694804 110015 694807
rect 576578 694804 576584 694816
rect 110003 694776 576584 694804
rect 110003 694773 110015 694776
rect 109957 694767 110015 694773
rect 576578 694764 576584 694776
rect 576636 694764 576642 694816
rect 1104 694640 6000 694736
rect 7852 694708 22140 694736
rect 125597 694739 125655 694745
rect 7852 694668 7880 694708
rect 125597 694705 125609 694739
rect 125643 694736 125655 694739
rect 140593 694739 140651 694745
rect 140593 694736 140605 694739
rect 125643 694708 140605 694736
rect 125643 694705 125655 694708
rect 125597 694699 125655 694705
rect 140593 694705 140605 694708
rect 140639 694705 140651 694739
rect 140593 694699 140651 694705
rect 152461 694739 152519 694745
rect 152461 694705 152473 694739
rect 152507 694736 152519 694739
rect 355597 694739 355655 694745
rect 355597 694736 355609 694739
rect 152507 694708 355609 694736
rect 152507 694705 152519 694708
rect 152461 694699 152519 694705
rect 355597 694705 355609 694708
rect 355643 694705 355655 694739
rect 355597 694699 355655 694705
rect 364981 694739 365039 694745
rect 364981 694705 364993 694739
rect 365027 694736 365039 694739
rect 374641 694739 374699 694745
rect 374641 694736 374653 694739
rect 365027 694708 374653 694736
rect 365027 694705 365039 694708
rect 364981 694699 365039 694705
rect 374641 694705 374653 694708
rect 374687 694705 374699 694739
rect 374641 694699 374699 694705
rect 384301 694739 384359 694745
rect 384301 694705 384313 694739
rect 384347 694736 384359 694739
rect 393961 694739 394019 694745
rect 393961 694736 393973 694739
rect 384347 694708 393973 694736
rect 384347 694705 384359 694708
rect 384301 694699 384359 694705
rect 393961 694705 393973 694708
rect 394007 694705 394019 694739
rect 393961 694699 394019 694705
rect 403621 694739 403679 694745
rect 403621 694705 403633 694739
rect 403667 694736 403679 694739
rect 413281 694739 413339 694745
rect 413281 694736 413293 694739
rect 403667 694708 413293 694736
rect 403667 694705 403679 694708
rect 403621 694699 403679 694705
rect 413281 694705 413293 694708
rect 413327 694705 413339 694739
rect 413281 694699 413339 694705
rect 422941 694739 422999 694745
rect 422941 694705 422953 694739
rect 422987 694736 422999 694739
rect 432601 694739 432659 694745
rect 432601 694736 432613 694739
rect 422987 694708 432613 694736
rect 422987 694705 422999 694708
rect 422941 694699 422999 694705
rect 432601 694705 432613 694708
rect 432647 694705 432659 694739
rect 432601 694699 432659 694705
rect 442261 694739 442319 694745
rect 442261 694705 442273 694739
rect 442307 694736 442319 694739
rect 450265 694739 450323 694745
rect 450265 694736 450277 694739
rect 442307 694708 450277 694736
rect 442307 694705 442319 694708
rect 442261 694699 442319 694705
rect 450265 694705 450277 694708
rect 450311 694705 450323 694739
rect 450265 694699 450323 694705
rect 459925 694739 459983 694745
rect 459925 694705 459937 694739
rect 459971 694736 459983 694739
rect 469585 694739 469643 694745
rect 469585 694736 469597 694739
rect 459971 694708 469597 694736
rect 459971 694705 459983 694708
rect 459925 694699 459983 694705
rect 469585 694705 469597 694708
rect 469631 694705 469643 694739
rect 469585 694699 469643 694705
rect 569310 694696 569316 694748
rect 569368 694736 569374 694748
rect 577498 694736 577504 694748
rect 569368 694708 577504 694736
rect 569368 694696 569374 694708
rect 577498 694696 577504 694708
rect 577556 694696 577562 694748
rect 7760 694640 7880 694668
rect 95789 694671 95847 694677
rect 3694 694560 3700 694612
rect 3752 694600 3758 694612
rect 7760 694600 7788 694640
rect 95789 694637 95801 694671
rect 95835 694668 95847 694671
rect 576486 694668 576492 694680
rect 95835 694640 576492 694668
rect 95835 694637 95847 694640
rect 95789 694631 95847 694637
rect 576486 694628 576492 694640
rect 576544 694628 576550 694680
rect 578000 694640 582820 694736
rect 3752 694572 7788 694600
rect 3752 694560 3758 694572
rect 7834 694560 7840 694612
rect 7892 694600 7898 694612
rect 497553 694603 497611 694609
rect 497553 694600 497565 694603
rect 7892 694572 497565 694600
rect 7892 694560 7898 694572
rect 497553 694569 497565 694572
rect 497599 694569 497611 694603
rect 497553 694563 497611 694569
rect 86405 694535 86463 694541
rect 86405 694501 86417 694535
rect 86451 694532 86463 694535
rect 577682 694532 577688 694544
rect 86451 694504 577688 694532
rect 86451 694501 86463 694504
rect 86405 694495 86463 694501
rect 577682 694492 577688 694504
rect 577740 694492 577746 694544
rect 81253 694467 81311 694473
rect 81253 694433 81265 694467
rect 81299 694464 81311 694467
rect 576394 694464 576400 694476
rect 81299 694436 576400 694464
rect 81299 694433 81311 694436
rect 81253 694427 81311 694433
rect 576394 694424 576400 694436
rect 576452 694424 576458 694476
rect 67453 694399 67511 694405
rect 67453 694365 67465 694399
rect 67499 694396 67511 694399
rect 575106 694396 575112 694408
rect 67499 694368 575112 694396
rect 67499 694365 67511 694368
rect 67453 694359 67511 694365
rect 575106 694356 575112 694368
rect 575164 694356 575170 694408
rect 3602 694288 3608 694340
rect 3660 694328 3666 694340
rect 511905 694331 511963 694337
rect 511905 694328 511917 694331
rect 3660 694300 511917 694328
rect 3660 694288 3666 694300
rect 511905 694297 511917 694300
rect 511951 694297 511963 694331
rect 511905 694291 511963 694297
rect 43717 694263 43775 694269
rect 43717 694229 43729 694263
rect 43763 694260 43775 694263
rect 576302 694260 576308 694272
rect 43763 694232 576308 694260
rect 43763 694229 43775 694232
rect 43717 694223 43775 694229
rect 576302 694220 576308 694232
rect 576360 694220 576366 694272
rect 29549 694195 29607 694201
rect 1104 694096 6000 694192
rect 29549 694161 29561 694195
rect 29595 694192 29607 694195
rect 576210 694192 576216 694204
rect 29595 694164 576216 694192
rect 29595 694161 29607 694164
rect 29549 694155 29607 694161
rect 576210 694152 576216 694164
rect 576268 694152 576274 694204
rect 578000 694096 582820 694192
rect 1104 693552 6000 693648
rect 578000 693552 582820 693648
rect 1104 693008 6000 693104
rect 578000 693008 582820 693104
rect 1104 692464 6000 692560
rect 578000 692464 582820 692560
rect 1104 691920 6000 692016
rect 578000 691920 582820 692016
rect 1104 691376 6000 691472
rect 578000 691376 582820 691472
rect 1104 690832 6000 690928
rect 578000 690832 582820 690928
rect 1104 690288 6000 690384
rect 578000 690288 582820 690384
rect 1104 689744 6000 689840
rect 578000 689744 582820 689840
rect 1104 689200 6000 689296
rect 578000 689200 582820 689296
rect 1104 688656 6000 688752
rect 578000 688656 582820 688752
rect 1104 688112 6000 688208
rect 578000 688112 582820 688208
rect 1104 687568 6000 687664
rect 578000 687568 582820 687664
rect 578694 687148 578700 687200
rect 578752 687188 578758 687200
rect 580902 687188 580908 687200
rect 578752 687160 580908 687188
rect 578752 687148 578758 687160
rect 580902 687148 580908 687160
rect 580960 687148 580966 687200
rect 1104 687024 6000 687120
rect 578000 687024 582820 687120
rect 1104 686480 6000 686576
rect 578000 686480 582820 686576
rect 1104 685936 6000 686032
rect 578000 685936 582820 686032
rect 1104 685392 6000 685488
rect 578000 685392 582820 685488
rect 1104 684848 6000 684944
rect 578000 684848 582820 684944
rect 1104 684304 6000 684400
rect 578000 684304 582820 684400
rect 1104 683760 6000 683856
rect 578000 683760 582820 683856
rect 1104 683216 6000 683312
rect 578000 683216 582820 683312
rect 1104 682672 6000 682768
rect 578000 682672 582820 682768
rect 2958 682524 2964 682576
rect 3016 682564 3022 682576
rect 5810 682564 5816 682576
rect 3016 682536 5816 682564
rect 3016 682524 3022 682536
rect 5810 682524 5816 682536
rect 5868 682524 5874 682576
rect 1104 682128 6000 682224
rect 578000 682128 582820 682224
rect 1104 681584 6000 681680
rect 578000 681584 582820 681680
rect 1104 681040 6000 681136
rect 578000 681040 582820 681136
rect 1104 680496 6000 680592
rect 578000 680496 582820 680592
rect 1104 679952 6000 680048
rect 578000 679952 582820 680048
rect 1104 679408 6000 679504
rect 578000 679408 582820 679504
rect 1104 678864 6000 678960
rect 578000 678864 582820 678960
rect 1104 678320 6000 678416
rect 578000 678320 582820 678416
rect 1104 677776 6000 677872
rect 578000 677776 582820 677872
rect 1104 677232 6000 677328
rect 578000 677232 582820 677328
rect 1104 676688 6000 676784
rect 578000 676688 582820 676784
rect 1104 676144 6000 676240
rect 578000 676144 582820 676240
rect 1104 675600 6000 675696
rect 578000 675600 582820 675696
rect 1104 675056 6000 675152
rect 578000 675056 582820 675152
rect 576026 674772 576032 674824
rect 576084 674812 576090 674824
rect 579798 674812 579804 674824
rect 576084 674784 579804 674812
rect 576084 674772 576090 674784
rect 579798 674772 579804 674784
rect 579856 674772 579862 674824
rect 1104 674512 6000 674608
rect 578000 674512 582820 674608
rect 1104 673968 6000 674064
rect 578000 673968 582820 674064
rect 1104 673424 6000 673520
rect 578000 673424 582820 673520
rect 1104 672880 6000 672976
rect 578000 672880 582820 672976
rect 1104 672336 6000 672432
rect 578000 672336 582820 672432
rect 1104 671792 6000 671888
rect 578000 671792 582820 671888
rect 1104 671248 6000 671344
rect 578000 671248 582820 671344
rect 1104 670704 6000 670800
rect 578000 670704 582820 670800
rect 1104 670160 6000 670256
rect 578000 670160 582820 670256
rect 1104 669616 6000 669712
rect 578000 669616 582820 669712
rect 1104 669072 6000 669168
rect 578000 669072 582820 669168
rect 1104 668528 6000 668624
rect 578000 668528 582820 668624
rect 2774 668176 2780 668228
rect 2832 668216 2838 668228
rect 5442 668216 5448 668228
rect 2832 668188 5448 668216
rect 2832 668176 2838 668188
rect 5442 668176 5448 668188
rect 5500 668176 5506 668228
rect 1104 667984 6000 668080
rect 578000 667984 582820 668080
rect 1104 667440 6000 667536
rect 578000 667440 582820 667536
rect 1104 666896 6000 666992
rect 578000 666896 582820 666992
rect 1104 666352 6000 666448
rect 578000 666352 582820 666448
rect 1104 665808 6000 665904
rect 578000 665808 582820 665904
rect 1104 665264 6000 665360
rect 578000 665264 582820 665360
rect 1104 664720 6000 664816
rect 578000 664720 582820 664816
rect 1104 664176 6000 664272
rect 578000 664176 582820 664272
rect 1104 663632 6000 663728
rect 578000 663632 582820 663728
rect 1104 663088 6000 663184
rect 578000 663088 582820 663184
rect 1104 662544 6000 662640
rect 578000 662544 582820 662640
rect 1104 662000 6000 662096
rect 578000 662000 582820 662096
rect 1104 661456 6000 661552
rect 578000 661456 582820 661552
rect 1104 660912 6000 661008
rect 578000 660912 582820 661008
rect 1104 660368 6000 660464
rect 578000 660368 582820 660464
rect 1104 659824 6000 659920
rect 578000 659824 582820 659920
rect 1104 659280 6000 659376
rect 578000 659280 582820 659376
rect 1104 658736 6000 658832
rect 578000 658736 582820 658832
rect 1104 658192 6000 658288
rect 578000 658192 582820 658288
rect 1104 657648 6000 657744
rect 578000 657648 582820 657744
rect 1104 657104 6000 657200
rect 578000 657104 582820 657200
rect 1104 656560 6000 656656
rect 578000 656560 582820 656656
rect 1104 656016 6000 656112
rect 578000 656016 582820 656112
rect 1104 655472 6000 655568
rect 578000 655472 582820 655568
rect 1104 654928 6000 655024
rect 578000 654928 582820 655024
rect 1104 654384 6000 654480
rect 578000 654384 582820 654480
rect 3050 653964 3056 654016
rect 3108 654004 3114 654016
rect 7282 654004 7288 654016
rect 3108 653976 7288 654004
rect 3108 653964 3114 653976
rect 7282 653964 7288 653976
rect 7340 653964 7346 654016
rect 1104 653840 6000 653936
rect 578000 653840 582820 653936
rect 1104 653296 6000 653392
rect 578000 653296 582820 653392
rect 1104 652752 6000 652848
rect 578000 652752 582820 652848
rect 1104 652208 6000 652304
rect 578000 652208 582820 652304
rect 1104 651664 6000 651760
rect 578000 651664 582820 651760
rect 577406 651312 577412 651364
rect 577464 651352 577470 651364
rect 579614 651352 579620 651364
rect 577464 651324 579620 651352
rect 577464 651312 577470 651324
rect 579614 651312 579620 651324
rect 579672 651312 579678 651364
rect 1104 651120 6000 651216
rect 578000 651120 582820 651216
rect 1104 650576 6000 650672
rect 578000 650576 582820 650672
rect 1104 650032 6000 650128
rect 578000 650032 582820 650128
rect 1104 649488 6000 649584
rect 578000 649488 582820 649584
rect 1104 648944 6000 649040
rect 578000 648944 582820 649040
rect 1104 648400 6000 648496
rect 578000 648400 582820 648496
rect 1104 647856 6000 647952
rect 578000 647856 582820 647952
rect 1104 647312 6000 647408
rect 578000 647312 582820 647408
rect 1104 646768 6000 646864
rect 578000 646768 582820 646864
rect 1104 646224 6000 646320
rect 578000 646224 582820 646320
rect 1104 645680 6000 645776
rect 578000 645680 582820 645776
rect 1104 645136 6000 645232
rect 578000 645136 582820 645232
rect 1104 644592 6000 644688
rect 578000 644592 582820 644688
rect 1104 644048 6000 644144
rect 578000 644048 582820 644144
rect 1104 643504 6000 643600
rect 578000 643504 582820 643600
rect 1104 642960 6000 643056
rect 578000 642960 582820 643056
rect 1104 642416 6000 642512
rect 578000 642416 582820 642512
rect 1104 641872 6000 641968
rect 578000 641872 582820 641968
rect 1104 641328 6000 641424
rect 578000 641328 582820 641424
rect 1104 640784 6000 640880
rect 578000 640784 582820 640880
rect 1104 640240 6000 640336
rect 578000 640240 582820 640336
rect 578786 640160 578792 640212
rect 578844 640200 578850 640212
rect 580902 640200 580908 640212
rect 578844 640172 580908 640200
rect 578844 640160 578850 640172
rect 580902 640160 580908 640172
rect 580960 640160 580966 640212
rect 1104 639696 6000 639792
rect 578000 639696 582820 639792
rect 1104 639152 6000 639248
rect 578000 639152 582820 639248
rect 1104 638608 6000 638704
rect 578000 638608 582820 638704
rect 1104 638064 6000 638160
rect 578000 638064 582820 638160
rect 1104 637520 6000 637616
rect 578000 637520 582820 637616
rect 1104 636976 6000 637072
rect 578000 636976 582820 637072
rect 1104 636432 6000 636528
rect 578000 636432 582820 636528
rect 1104 635888 6000 635984
rect 578000 635888 582820 635984
rect 1104 635344 6000 635440
rect 578000 635344 582820 635440
rect 1104 634800 6000 634896
rect 578000 634800 582820 634896
rect 1104 634256 6000 634352
rect 578000 634256 582820 634352
rect 1104 633712 6000 633808
rect 578000 633712 582820 633808
rect 1104 633168 6000 633264
rect 578000 633168 582820 633264
rect 1104 632624 6000 632720
rect 578000 632624 582820 632720
rect 1104 632080 6000 632176
rect 578000 632080 582820 632176
rect 1104 631536 6000 631632
rect 578000 631536 582820 631632
rect 1104 630992 6000 631088
rect 578000 630992 582820 631088
rect 1104 630448 6000 630544
rect 578000 630448 582820 630544
rect 1104 629904 6000 630000
rect 578000 629904 582820 630000
rect 1104 629360 6000 629456
rect 578000 629360 582820 629456
rect 1104 628816 6000 628912
rect 578000 628816 582820 628912
rect 1104 628272 6000 628368
rect 578000 628272 582820 628368
rect 575474 627852 575480 627904
rect 575532 627892 575538 627904
rect 579798 627892 579804 627904
rect 575532 627864 579804 627892
rect 575532 627852 575538 627864
rect 579798 627852 579804 627864
rect 579856 627852 579862 627904
rect 1104 627728 6000 627824
rect 578000 627728 582820 627824
rect 1104 627184 6000 627280
rect 578000 627184 582820 627280
rect 1104 626640 6000 626736
rect 578000 626640 582820 626736
rect 1104 626096 6000 626192
rect 578000 626096 582820 626192
rect 1104 625552 6000 625648
rect 578000 625552 582820 625648
rect 1104 625008 6000 625104
rect 578000 625008 582820 625104
rect 2958 624860 2964 624912
rect 3016 624900 3022 624912
rect 5902 624900 5908 624912
rect 3016 624872 5908 624900
rect 3016 624860 3022 624872
rect 5902 624860 5908 624872
rect 5960 624860 5966 624912
rect 1104 624464 6000 624560
rect 578000 624464 582820 624560
rect 1104 623920 6000 624016
rect 578000 623920 582820 624016
rect 1104 623376 6000 623472
rect 578000 623376 582820 623472
rect 1104 622832 6000 622928
rect 578000 622832 582820 622928
rect 1104 622288 6000 622384
rect 578000 622288 582820 622384
rect 1104 621744 6000 621840
rect 578000 621744 582820 621840
rect 1104 621200 6000 621296
rect 578000 621200 582820 621296
rect 1104 620656 6000 620752
rect 578000 620656 582820 620752
rect 1104 620112 6000 620208
rect 578000 620112 582820 620208
rect 1104 619568 6000 619664
rect 578000 619568 582820 619664
rect 1104 619024 6000 619120
rect 578000 619024 582820 619120
rect 1104 618480 6000 618576
rect 578000 618480 582820 618576
rect 1104 617936 6000 618032
rect 578000 617936 582820 618032
rect 1104 617392 6000 617488
rect 578000 617392 582820 617488
rect 1104 616848 6000 616944
rect 578000 616848 582820 616944
rect 1104 616304 6000 616400
rect 578000 616304 582820 616400
rect 1104 615760 6000 615856
rect 578000 615760 582820 615856
rect 1104 615216 6000 615312
rect 578000 615216 582820 615312
rect 1104 614672 6000 614768
rect 578000 614672 582820 614768
rect 1104 614128 6000 614224
rect 578000 614128 582820 614224
rect 1104 613584 6000 613680
rect 578000 613584 582820 613680
rect 1104 613040 6000 613136
rect 578000 613040 582820 613136
rect 1104 612496 6000 612592
rect 578000 612496 582820 612592
rect 1104 611952 6000 612048
rect 578000 611952 582820 612048
rect 1104 611408 6000 611504
rect 578000 611408 582820 611504
rect 1104 610864 6000 610960
rect 578000 610864 582820 610960
rect 1104 610320 6000 610416
rect 578000 610320 582820 610416
rect 1104 609776 6000 609872
rect 578000 609776 582820 609872
rect 1104 609232 6000 609328
rect 578000 609232 582820 609328
rect 1104 608688 6000 608784
rect 578000 608688 582820 608784
rect 1104 608144 6000 608240
rect 578000 608144 582820 608240
rect 1104 607600 6000 607696
rect 578000 607600 582820 607696
rect 1104 607056 6000 607152
rect 578000 607056 582820 607152
rect 1104 606512 6000 606608
rect 578000 606512 582820 606608
rect 1104 605968 6000 606064
rect 578000 605968 582820 606064
rect 1104 605424 6000 605520
rect 578000 605424 582820 605520
rect 1104 604880 6000 604976
rect 578000 604880 582820 604976
rect 1104 604336 6000 604432
rect 578000 604336 582820 604432
rect 578142 604256 578148 604308
rect 578200 604296 578206 604308
rect 579614 604296 579620 604308
rect 578200 604268 579620 604296
rect 578200 604256 578206 604268
rect 579614 604256 579620 604268
rect 579672 604256 579678 604308
rect 1104 603792 6000 603888
rect 578000 603792 582820 603888
rect 1104 603248 6000 603344
rect 578000 603248 582820 603344
rect 1104 602704 6000 602800
rect 578000 602704 582820 602800
rect 1104 602160 6000 602256
rect 578000 602160 582820 602256
rect 1104 601616 6000 601712
rect 578000 601616 582820 601712
rect 1104 601072 6000 601168
rect 578000 601072 582820 601168
rect 1104 600528 6000 600624
rect 578000 600528 582820 600624
rect 1104 599984 6000 600080
rect 578000 599984 582820 600080
rect 1104 599440 6000 599536
rect 578000 599440 582820 599536
rect 1104 598896 6000 598992
rect 578000 598896 582820 598992
rect 1104 598352 6000 598448
rect 578000 598352 582820 598448
rect 1104 597808 6000 597904
rect 578000 597808 582820 597904
rect 1104 597264 6000 597360
rect 578000 597264 582820 597360
rect 1104 596720 6000 596816
rect 578000 596720 582820 596816
rect 1104 596176 6000 596272
rect 578000 596176 582820 596272
rect 3142 596028 3148 596080
rect 3200 596068 3206 596080
rect 7374 596068 7380 596080
rect 3200 596040 7380 596068
rect 3200 596028 3206 596040
rect 7374 596028 7380 596040
rect 7432 596028 7438 596080
rect 1104 595632 6000 595728
rect 578000 595632 582820 595728
rect 1104 595088 6000 595184
rect 578000 595088 582820 595184
rect 1104 594544 6000 594640
rect 578000 594544 582820 594640
rect 1104 594000 6000 594096
rect 578000 594000 582820 594096
rect 1104 593456 6000 593552
rect 578000 593456 582820 593552
rect 1104 592912 6000 593008
rect 578000 592912 582820 593008
rect 1104 592368 6000 592464
rect 578000 592368 582820 592464
rect 1104 591824 6000 591920
rect 578000 591824 582820 591920
rect 1104 591280 6000 591376
rect 578000 591280 582820 591376
rect 1104 590736 6000 590832
rect 578000 590736 582820 590832
rect 1104 590192 6000 590288
rect 578000 590192 582820 590288
rect 1104 589648 6000 589744
rect 578000 589648 582820 589744
rect 1104 589104 6000 589200
rect 578000 589104 582820 589200
rect 1104 588560 6000 588656
rect 578000 588560 582820 588656
rect 1104 588016 6000 588112
rect 578000 588016 582820 588112
rect 1104 587472 6000 587568
rect 578000 587472 582820 587568
rect 1104 586928 6000 587024
rect 578000 586928 582820 587024
rect 1104 586384 6000 586480
rect 578000 586384 582820 586480
rect 1104 585840 6000 585936
rect 578000 585840 582820 585936
rect 1104 585296 6000 585392
rect 578000 585296 582820 585392
rect 1104 584752 6000 584848
rect 578000 584752 582820 584848
rect 1104 584208 6000 584304
rect 578000 584208 582820 584304
rect 1104 583664 6000 583760
rect 578000 583664 582820 583760
rect 1104 583120 6000 583216
rect 578000 583120 582820 583216
rect 1104 582576 6000 582672
rect 578000 582576 582820 582672
rect 1104 582032 6000 582128
rect 578000 582032 582820 582128
rect 1104 581488 6000 581584
rect 578000 581488 582820 581584
rect 1104 580944 6000 581040
rect 578000 580944 582820 581040
rect 575382 580864 575388 580916
rect 575440 580904 575446 580916
rect 580166 580904 580172 580916
rect 575440 580876 580172 580904
rect 575440 580864 575446 580876
rect 580166 580864 580172 580876
rect 580224 580864 580230 580916
rect 1104 580400 6000 580496
rect 578000 580400 582820 580496
rect 1104 579856 6000 579952
rect 578000 579856 582820 579952
rect 1104 579312 6000 579408
rect 578000 579312 582820 579408
rect 1104 578768 6000 578864
rect 578000 578768 582820 578864
rect 1104 578224 6000 578320
rect 578000 578224 582820 578320
rect 1104 577680 6000 577776
rect 578000 577680 582820 577776
rect 1104 577136 6000 577232
rect 578000 577136 582820 577232
rect 1104 576592 6000 576688
rect 578000 576592 582820 576688
rect 1104 576048 6000 576144
rect 578000 576048 582820 576144
rect 1104 575504 6000 575600
rect 578000 575504 582820 575600
rect 1104 574960 6000 575056
rect 578000 574960 582820 575056
rect 1104 574416 6000 574512
rect 578000 574416 582820 574512
rect 1104 573872 6000 573968
rect 578000 573872 582820 573968
rect 1104 573328 6000 573424
rect 578000 573328 582820 573424
rect 1104 572784 6000 572880
rect 578000 572784 582820 572880
rect 1104 572240 6000 572336
rect 578000 572240 582820 572336
rect 1104 571696 6000 571792
rect 578000 571696 582820 571792
rect 1104 571152 6000 571248
rect 578000 571152 582820 571248
rect 1104 570608 6000 570704
rect 578000 570608 582820 570704
rect 1104 570064 6000 570160
rect 578000 570064 582820 570160
rect 1104 569520 6000 569616
rect 578000 569520 582820 569616
rect 1104 568976 6000 569072
rect 578000 568976 582820 569072
rect 1104 568432 6000 568528
rect 578000 568432 582820 568528
rect 1104 567888 6000 567984
rect 578000 567888 582820 567984
rect 3050 567604 3056 567656
rect 3108 567644 3114 567656
rect 5994 567644 6000 567656
rect 3108 567616 6000 567644
rect 3108 567604 3114 567616
rect 5994 567604 6000 567616
rect 6052 567604 6058 567656
rect 1104 567344 6000 567440
rect 578000 567344 582820 567440
rect 1104 566800 6000 566896
rect 578000 566800 582820 566896
rect 1104 566256 6000 566352
rect 578000 566256 582820 566352
rect 1104 565712 6000 565808
rect 578000 565712 582820 565808
rect 1104 565168 6000 565264
rect 578000 565168 582820 565264
rect 1104 564624 6000 564720
rect 578000 564624 582820 564720
rect 1104 564080 6000 564176
rect 578000 564080 582820 564176
rect 1104 563536 6000 563632
rect 578000 563536 582820 563632
rect 1104 562992 6000 563088
rect 578000 562992 582820 563088
rect 1104 562448 6000 562544
rect 578000 562448 582820 562544
rect 1104 561904 6000 562000
rect 578000 561904 582820 562000
rect 1104 561360 6000 561456
rect 578000 561360 582820 561456
rect 1104 560816 6000 560912
rect 578000 560816 582820 560912
rect 1104 560272 6000 560368
rect 578000 560272 582820 560368
rect 1104 559728 6000 559824
rect 578000 559728 582820 559824
rect 1104 559184 6000 559280
rect 578000 559184 582820 559280
rect 1104 558640 6000 558736
rect 578000 558640 582820 558736
rect 1104 558096 6000 558192
rect 578000 558096 582820 558192
rect 1104 557552 6000 557648
rect 578000 557552 582820 557648
rect 578050 557336 578056 557388
rect 578108 557376 578114 557388
rect 579614 557376 579620 557388
rect 578108 557348 579620 557376
rect 578108 557336 578114 557348
rect 579614 557336 579620 557348
rect 579672 557336 579678 557388
rect 1104 557008 6000 557104
rect 578000 557008 582820 557104
rect 1104 556464 6000 556560
rect 578000 556464 582820 556560
rect 1104 555920 6000 556016
rect 578000 555920 582820 556016
rect 1104 555376 6000 555472
rect 578000 555376 582820 555472
rect 1104 554832 6000 554928
rect 578000 554832 582820 554928
rect 1104 554288 6000 554384
rect 578000 554288 582820 554384
rect 1104 553744 6000 553840
rect 578000 553744 582820 553840
rect 1104 553200 6000 553296
rect 578000 553200 582820 553296
rect 1104 552656 6000 552752
rect 578000 552656 582820 552752
rect 1104 552112 6000 552208
rect 578000 552112 582820 552208
rect 1104 551568 6000 551664
rect 578000 551568 582820 551664
rect 1104 551024 6000 551120
rect 578000 551024 582820 551120
rect 1104 550480 6000 550576
rect 578000 550480 582820 550576
rect 1104 549936 6000 550032
rect 578000 549936 582820 550032
rect 1104 549392 6000 549488
rect 578000 549392 582820 549488
rect 1104 548848 6000 548944
rect 578000 548848 582820 548944
rect 1104 548304 6000 548400
rect 578000 548304 582820 548400
rect 1104 547760 6000 547856
rect 578000 547760 582820 547856
rect 1104 547216 6000 547312
rect 578000 547216 582820 547312
rect 1104 546672 6000 546768
rect 578000 546672 582820 546768
rect 1104 546128 6000 546224
rect 578000 546128 582820 546224
rect 1104 545584 6000 545680
rect 578000 545584 582820 545680
rect 1104 545040 6000 545136
rect 578000 545040 582820 545136
rect 1104 544496 6000 544592
rect 578000 544496 582820 544592
rect 1104 543952 6000 544048
rect 578000 543952 582820 544048
rect 1104 543408 6000 543504
rect 578000 543408 582820 543504
rect 1104 542864 6000 542960
rect 578000 542864 582820 542960
rect 1104 542320 6000 542416
rect 578000 542320 582820 542416
rect 1104 541776 6000 541872
rect 578000 541776 582820 541872
rect 1104 541232 6000 541328
rect 578000 541232 582820 541328
rect 1104 540688 6000 540784
rect 578000 540688 582820 540784
rect 1104 540144 6000 540240
rect 578000 540144 582820 540240
rect 1104 539600 6000 539696
rect 578000 539600 582820 539696
rect 3878 539384 3884 539436
rect 3936 539424 3942 539436
rect 5350 539424 5356 539436
rect 3936 539396 5356 539424
rect 3936 539384 3942 539396
rect 5350 539384 5356 539396
rect 5408 539384 5414 539436
rect 1104 539056 6000 539152
rect 578000 539056 582820 539152
rect 1104 538512 6000 538608
rect 578000 538512 582820 538608
rect 1104 537968 6000 538064
rect 578000 537968 582820 538064
rect 1104 537424 6000 537520
rect 578000 537424 582820 537520
rect 1104 536880 6000 536976
rect 578000 536880 582820 536976
rect 1104 536336 6000 536432
rect 578000 536336 582820 536432
rect 1104 535792 6000 535888
rect 578000 535792 582820 535888
rect 1104 535248 6000 535344
rect 578000 535248 582820 535344
rect 1104 534704 6000 534800
rect 578000 534704 582820 534800
rect 1104 534160 6000 534256
rect 578000 534160 582820 534256
rect 575290 534012 575296 534064
rect 575348 534052 575354 534064
rect 579798 534052 579804 534064
rect 575348 534024 579804 534052
rect 575348 534012 575354 534024
rect 579798 534012 579804 534024
rect 579856 534012 579862 534064
rect 1104 533616 6000 533712
rect 578000 533616 582820 533712
rect 1104 533072 6000 533168
rect 578000 533072 582820 533168
rect 1104 532528 6000 532624
rect 578000 532528 582820 532624
rect 1104 531984 6000 532080
rect 578000 531984 582820 532080
rect 1104 531440 6000 531536
rect 578000 531440 582820 531536
rect 1104 530896 6000 530992
rect 578000 530896 582820 530992
rect 1104 530352 6000 530448
rect 578000 530352 582820 530448
rect 1104 529808 6000 529904
rect 578000 529808 582820 529904
rect 1104 529264 6000 529360
rect 578000 529264 582820 529360
rect 1104 528720 6000 528816
rect 578000 528720 582820 528816
rect 1104 528176 6000 528272
rect 578000 528176 582820 528272
rect 1104 527632 6000 527728
rect 578000 527632 582820 527728
rect 1104 527088 6000 527184
rect 578000 527088 582820 527184
rect 1104 526544 6000 526640
rect 578000 526544 582820 526640
rect 1104 526000 6000 526096
rect 578000 526000 582820 526096
rect 1104 525456 6000 525552
rect 578000 525456 582820 525552
rect 1104 524912 6000 525008
rect 578000 524912 582820 525008
rect 1104 524368 6000 524464
rect 578000 524368 582820 524464
rect 1104 523824 6000 523920
rect 578000 523824 582820 523920
rect 1104 523280 6000 523376
rect 578000 523280 582820 523376
rect 1104 522736 6000 522832
rect 578000 522736 582820 522832
rect 1104 522192 6000 522288
rect 578000 522192 582820 522288
rect 1104 521648 6000 521744
rect 578000 521648 582820 521744
rect 1104 521104 6000 521200
rect 578000 521104 582820 521200
rect 1104 520560 6000 520656
rect 578000 520560 582820 520656
rect 1104 520016 6000 520112
rect 578000 520016 582820 520112
rect 1104 519472 6000 519568
rect 578000 519472 582820 519568
rect 1104 518928 6000 519024
rect 578000 518928 582820 519024
rect 1104 518384 6000 518480
rect 578000 518384 582820 518480
rect 1104 517840 6000 517936
rect 578000 517840 582820 517936
rect 1104 517296 6000 517392
rect 578000 517296 582820 517392
rect 1104 516752 6000 516848
rect 578000 516752 582820 516848
rect 1104 516208 6000 516304
rect 578000 516208 582820 516304
rect 1104 515664 6000 515760
rect 578000 515664 582820 515760
rect 1104 515120 6000 515216
rect 578000 515120 582820 515216
rect 1104 514576 6000 514672
rect 578000 514576 582820 514672
rect 1104 514032 6000 514128
rect 578000 514032 582820 514128
rect 1104 513488 6000 513584
rect 578000 513488 582820 513584
rect 1104 512944 6000 513040
rect 578000 512944 582820 513040
rect 1104 512400 6000 512496
rect 578000 512400 582820 512496
rect 1104 511856 6000 511952
rect 578000 511856 582820 511952
rect 1104 511312 6000 511408
rect 578000 511312 582820 511408
rect 1104 510768 6000 510864
rect 578000 510768 582820 510864
rect 577958 510552 577964 510604
rect 578016 510592 578022 510604
rect 580074 510592 580080 510604
rect 578016 510564 580080 510592
rect 578016 510552 578022 510564
rect 580074 510552 580080 510564
rect 580132 510552 580138 510604
rect 3050 510348 3056 510400
rect 3108 510388 3114 510400
rect 6086 510388 6092 510400
rect 3108 510360 6092 510388
rect 3108 510348 3114 510360
rect 6086 510348 6092 510360
rect 6144 510348 6150 510400
rect 1104 510224 6000 510320
rect 578000 510224 582820 510320
rect 1104 509680 6000 509776
rect 578000 509680 582820 509776
rect 1104 509136 6000 509232
rect 578000 509136 582820 509232
rect 1104 508592 6000 508688
rect 578000 508592 582820 508688
rect 1104 508048 6000 508144
rect 578000 508048 582820 508144
rect 1104 507504 6000 507600
rect 578000 507504 582820 507600
rect 1104 506960 6000 507056
rect 578000 506960 582820 507056
rect 1104 506416 6000 506512
rect 578000 506416 582820 506512
rect 1104 505872 6000 505968
rect 578000 505872 582820 505968
rect 1104 505328 6000 505424
rect 578000 505328 582820 505424
rect 1104 504784 6000 504880
rect 578000 504784 582820 504880
rect 1104 504240 6000 504336
rect 578000 504240 582820 504336
rect 1104 503696 6000 503792
rect 578000 503696 582820 503792
rect 1104 503152 6000 503248
rect 578000 503152 582820 503248
rect 1104 502608 6000 502704
rect 578000 502608 582820 502704
rect 1104 502064 6000 502160
rect 578000 502064 582820 502160
rect 1104 501520 6000 501616
rect 578000 501520 582820 501616
rect 1104 500976 6000 501072
rect 578000 500976 582820 501072
rect 1104 500432 6000 500528
rect 578000 500432 582820 500528
rect 1104 499888 6000 499984
rect 578000 499888 582820 499984
rect 1104 499344 6000 499440
rect 578000 499344 582820 499440
rect 1104 498800 6000 498896
rect 578000 498800 582820 498896
rect 1104 498256 6000 498352
rect 578000 498256 582820 498352
rect 1104 497712 6000 497808
rect 578000 497712 582820 497808
rect 1104 497168 6000 497264
rect 578000 497168 582820 497264
rect 1104 496624 6000 496720
rect 578000 496624 582820 496720
rect 1104 496080 6000 496176
rect 578000 496080 582820 496176
rect 1104 495536 6000 495632
rect 578000 495536 582820 495632
rect 1104 494992 6000 495088
rect 578000 494992 582820 495088
rect 1104 494448 6000 494544
rect 578000 494448 582820 494544
rect 1104 493904 6000 494000
rect 578000 493904 582820 494000
rect 1104 493360 6000 493456
rect 578000 493360 582820 493456
rect 1104 492816 6000 492912
rect 578000 492816 582820 492912
rect 1104 492272 6000 492368
rect 578000 492272 582820 492368
rect 1104 491728 6000 491824
rect 578000 491728 582820 491824
rect 1104 491184 6000 491280
rect 578000 491184 582820 491280
rect 1104 490640 6000 490736
rect 578000 490640 582820 490736
rect 1104 490096 6000 490192
rect 578000 490096 582820 490192
rect 1104 489552 6000 489648
rect 578000 489552 582820 489648
rect 1104 489008 6000 489104
rect 578000 489008 582820 489104
rect 1104 488464 6000 488560
rect 578000 488464 582820 488560
rect 1104 487920 6000 488016
rect 578000 487920 582820 488016
rect 1104 487376 6000 487472
rect 578000 487376 582820 487472
rect 575198 487092 575204 487144
rect 575256 487132 575262 487144
rect 580166 487132 580172 487144
rect 575256 487104 580172 487132
rect 575256 487092 575262 487104
rect 580166 487092 580172 487104
rect 580224 487092 580230 487144
rect 1104 486832 6000 486928
rect 578000 486832 582820 486928
rect 1104 486288 6000 486384
rect 578000 486288 582820 486384
rect 1104 485744 6000 485840
rect 578000 485744 582820 485840
rect 1104 485200 6000 485296
rect 578000 485200 582820 485296
rect 1104 484656 6000 484752
rect 578000 484656 582820 484752
rect 1104 484112 6000 484208
rect 578000 484112 582820 484208
rect 1104 483568 6000 483664
rect 578000 483568 582820 483664
rect 1104 483024 6000 483120
rect 578000 483024 582820 483120
rect 1104 482480 6000 482576
rect 578000 482480 582820 482576
rect 1104 481936 6000 482032
rect 578000 481936 582820 482032
rect 1104 481392 6000 481488
rect 578000 481392 582820 481488
rect 3326 481108 3332 481160
rect 3384 481148 3390 481160
rect 7466 481148 7472 481160
rect 3384 481120 7472 481148
rect 3384 481108 3390 481120
rect 7466 481108 7472 481120
rect 7524 481108 7530 481160
rect 1104 480848 6000 480944
rect 578000 480848 582820 480944
rect 1104 480304 6000 480400
rect 578000 480304 582820 480400
rect 1104 479760 6000 479856
rect 578000 479760 582820 479856
rect 1104 479216 6000 479312
rect 578000 479216 582820 479312
rect 1104 478672 6000 478768
rect 578000 478672 582820 478768
rect 1104 478128 6000 478224
rect 578000 478128 582820 478224
rect 1104 477584 6000 477680
rect 578000 477584 582820 477680
rect 1104 477040 6000 477136
rect 578000 477040 582820 477136
rect 1104 476496 6000 476592
rect 578000 476496 582820 476592
rect 1104 475952 6000 476048
rect 578000 475952 582820 476048
rect 1104 475408 6000 475504
rect 578000 475408 582820 475504
rect 1104 474864 6000 474960
rect 578000 474864 582820 474960
rect 1104 474320 6000 474416
rect 578000 474320 582820 474416
rect 1104 473776 6000 473872
rect 578000 473776 582820 473872
rect 1104 473232 6000 473328
rect 578000 473232 582820 473328
rect 1104 472688 6000 472784
rect 578000 472688 582820 472784
rect 1104 472144 6000 472240
rect 578000 472144 582820 472240
rect 1104 471600 6000 471696
rect 578000 471600 582820 471696
rect 1104 471056 6000 471152
rect 578000 471056 582820 471152
rect 1104 470512 6000 470608
rect 578000 470512 582820 470608
rect 1104 469968 6000 470064
rect 578000 469968 582820 470064
rect 1104 469424 6000 469520
rect 578000 469424 582820 469520
rect 1104 468880 6000 468976
rect 578000 468880 582820 468976
rect 1104 468336 6000 468432
rect 578000 468336 582820 468432
rect 1104 467792 6000 467888
rect 578000 467792 582820 467888
rect 1104 467248 6000 467344
rect 578000 467248 582820 467344
rect 1104 466704 6000 466800
rect 578000 466704 582820 466800
rect 1104 466160 6000 466256
rect 578000 466160 582820 466256
rect 1104 465616 6000 465712
rect 578000 465616 582820 465712
rect 1104 465072 6000 465168
rect 578000 465072 582820 465168
rect 1104 464528 6000 464624
rect 578000 464528 582820 464624
rect 1104 463984 6000 464080
rect 578000 463984 582820 464080
rect 1104 463440 6000 463536
rect 578000 463440 582820 463536
rect 1104 462896 6000 462992
rect 578000 462896 582820 462992
rect 1104 462352 6000 462448
rect 578000 462352 582820 462448
rect 1104 461808 6000 461904
rect 578000 461808 582820 461904
rect 1104 461264 6000 461360
rect 578000 461264 582820 461360
rect 1104 460720 6000 460816
rect 578000 460720 582820 460816
rect 1104 460176 6000 460272
rect 578000 460176 582820 460272
rect 1104 459632 6000 459728
rect 578000 459632 582820 459728
rect 1104 459088 6000 459184
rect 578000 459088 582820 459184
rect 1104 458544 6000 458640
rect 578000 458544 582820 458640
rect 1104 458000 6000 458096
rect 578000 458000 582820 458096
rect 1104 457456 6000 457552
rect 578000 457456 582820 457552
rect 1104 456912 6000 457008
rect 578000 456912 582820 457008
rect 1104 456368 6000 456464
rect 578000 456368 582820 456464
rect 1104 455824 6000 455920
rect 578000 455824 582820 455920
rect 1104 455280 6000 455376
rect 578000 455280 582820 455376
rect 1104 454736 6000 454832
rect 578000 454736 582820 454832
rect 1104 454192 6000 454288
rect 578000 454192 582820 454288
rect 1104 453648 6000 453744
rect 578000 453648 582820 453744
rect 1104 453104 6000 453200
rect 578000 453104 582820 453200
rect 1104 452560 6000 452656
rect 578000 452560 582820 452656
rect 3326 452412 3332 452464
rect 3384 452452 3390 452464
rect 6822 452452 6828 452464
rect 3384 452424 6828 452452
rect 3384 452412 3390 452424
rect 6822 452412 6828 452424
rect 6880 452412 6886 452464
rect 1104 452016 6000 452112
rect 578000 452016 582820 452112
rect 1104 451472 6000 451568
rect 578000 451472 582820 451568
rect 1104 450928 6000 451024
rect 578000 450928 582820 451024
rect 1104 450384 6000 450480
rect 578000 450384 582820 450480
rect 1104 449840 6000 449936
rect 578000 449840 582820 449936
rect 1104 449296 6000 449392
rect 578000 449296 582820 449392
rect 1104 448752 6000 448848
rect 578000 448752 582820 448848
rect 1104 448208 6000 448304
rect 578000 448208 582820 448304
rect 1104 447664 6000 447760
rect 578000 447664 582820 447760
rect 1104 447120 6000 447216
rect 578000 447120 582820 447216
rect 1104 446576 6000 446672
rect 578000 446576 582820 446672
rect 1104 446032 6000 446128
rect 578000 446032 582820 446128
rect 1104 445488 6000 445584
rect 578000 445488 582820 445584
rect 1104 444944 6000 445040
rect 578000 444944 582820 445040
rect 1104 444400 6000 444496
rect 578000 444400 582820 444496
rect 1104 443856 6000 443952
rect 578000 443856 582820 443952
rect 1104 443312 6000 443408
rect 578000 443312 582820 443408
rect 1104 442768 6000 442864
rect 578000 442768 582820 442864
rect 1104 442224 6000 442320
rect 578000 442224 582820 442320
rect 1104 441680 6000 441776
rect 578000 441680 582820 441776
rect 1104 441136 6000 441232
rect 578000 441136 582820 441232
rect 1104 440592 6000 440688
rect 578000 440592 582820 440688
rect 576762 440172 576768 440224
rect 576820 440212 576826 440224
rect 579982 440212 579988 440224
rect 576820 440184 579988 440212
rect 576820 440172 576826 440184
rect 579982 440172 579988 440184
rect 580040 440172 580046 440224
rect 1104 440048 6000 440144
rect 578000 440048 582820 440144
rect 1104 439504 6000 439600
rect 578000 439504 582820 439600
rect 1104 438960 6000 439056
rect 578000 438960 582820 439056
rect 3326 438880 3332 438932
rect 3384 438920 3390 438932
rect 5258 438920 5264 438932
rect 3384 438892 5264 438920
rect 3384 438880 3390 438892
rect 5258 438880 5264 438892
rect 5316 438880 5322 438932
rect 1104 438416 6000 438512
rect 578000 438416 582820 438512
rect 1104 437872 6000 437968
rect 578000 437872 582820 437968
rect 1104 437328 6000 437424
rect 578000 437328 582820 437424
rect 1104 436784 6000 436880
rect 578000 436784 582820 436880
rect 1104 436240 6000 436336
rect 578000 436240 582820 436336
rect 1104 435696 6000 435792
rect 578000 435696 582820 435792
rect 1104 435152 6000 435248
rect 578000 435152 582820 435248
rect 1104 434608 6000 434704
rect 578000 434608 582820 434704
rect 1104 434064 6000 434160
rect 578000 434064 582820 434160
rect 1104 433520 6000 433616
rect 578000 433520 582820 433616
rect 1104 432976 6000 433072
rect 578000 432976 582820 433072
rect 1104 432432 6000 432528
rect 578000 432432 582820 432528
rect 1104 431888 6000 431984
rect 578000 431888 582820 431984
rect 1104 431344 6000 431440
rect 578000 431344 582820 431440
rect 1104 430800 6000 430896
rect 578000 430800 582820 430896
rect 1104 430256 6000 430352
rect 578000 430256 582820 430352
rect 1104 429712 6000 429808
rect 578000 429712 582820 429808
rect 1104 429168 6000 429264
rect 578000 429168 582820 429264
rect 1104 428624 6000 428720
rect 578000 428624 582820 428720
rect 1104 428080 6000 428176
rect 578000 428080 582820 428176
rect 1104 427536 6000 427632
rect 578000 427536 582820 427632
rect 1104 426992 6000 427088
rect 578000 426992 582820 427088
rect 1104 426448 6000 426544
rect 578000 426448 582820 426544
rect 1104 425904 6000 426000
rect 578000 425904 582820 426000
rect 1104 425360 6000 425456
rect 578000 425360 582820 425456
rect 1104 424816 6000 424912
rect 578000 424816 582820 424912
rect 1104 424272 6000 424368
rect 578000 424272 582820 424368
rect 2866 423852 2872 423904
rect 2924 423892 2930 423904
rect 8202 423892 8208 423904
rect 2924 423864 8208 423892
rect 2924 423852 2930 423864
rect 8202 423852 8208 423864
rect 8260 423852 8266 423904
rect 1104 423728 6000 423824
rect 578000 423728 582820 423824
rect 1104 423184 6000 423280
rect 578000 423184 582820 423280
rect 1104 422640 6000 422736
rect 578000 422640 582820 422736
rect 1104 422096 6000 422192
rect 578000 422096 582820 422192
rect 1104 421552 6000 421648
rect 578000 421552 582820 421648
rect 1104 421008 6000 421104
rect 578000 421008 582820 421104
rect 1104 420464 6000 420560
rect 578000 420464 582820 420560
rect 1104 419920 6000 420016
rect 578000 419920 582820 420016
rect 1104 419376 6000 419472
rect 578000 419376 582820 419472
rect 1104 418832 6000 418928
rect 578000 418832 582820 418928
rect 1104 418288 6000 418384
rect 578000 418288 582820 418384
rect 1104 417744 6000 417840
rect 578000 417744 582820 417840
rect 1104 417200 6000 417296
rect 578000 417200 582820 417296
rect 1104 416656 6000 416752
rect 578000 416656 582820 416752
rect 577866 416576 577872 416628
rect 577924 416616 577930 416628
rect 579614 416616 579620 416628
rect 577924 416588 579620 416616
rect 577924 416576 577930 416588
rect 579614 416576 579620 416588
rect 579672 416576 579678 416628
rect 1104 416112 6000 416208
rect 578000 416112 582820 416208
rect 1104 415568 6000 415664
rect 578000 415568 582820 415664
rect 1104 415024 6000 415120
rect 578000 415024 582820 415120
rect 1104 414480 6000 414576
rect 578000 414480 582820 414576
rect 1104 413936 6000 414032
rect 578000 413936 582820 414032
rect 1104 413392 6000 413488
rect 578000 413392 582820 413488
rect 1104 412848 6000 412944
rect 578000 412848 582820 412944
rect 1104 412304 6000 412400
rect 578000 412304 582820 412400
rect 1104 411760 6000 411856
rect 578000 411760 582820 411856
rect 1104 411216 6000 411312
rect 578000 411216 582820 411312
rect 1104 410672 6000 410768
rect 578000 410672 582820 410768
rect 1104 410128 6000 410224
rect 578000 410128 582820 410224
rect 1104 409584 6000 409680
rect 578000 409584 582820 409680
rect 1104 409040 6000 409136
rect 578000 409040 582820 409136
rect 1104 408496 6000 408592
rect 578000 408496 582820 408592
rect 1104 407952 6000 408048
rect 578000 407952 582820 408048
rect 1104 407408 6000 407504
rect 578000 407408 582820 407504
rect 1104 406864 6000 406960
rect 578000 406864 582820 406960
rect 1104 406320 6000 406416
rect 578000 406320 582820 406416
rect 1104 405776 6000 405872
rect 578000 405776 582820 405872
rect 1104 405232 6000 405328
rect 578000 405232 582820 405328
rect 1104 404688 6000 404784
rect 578000 404688 582820 404784
rect 1104 404144 6000 404240
rect 578000 404144 582820 404240
rect 1104 403600 6000 403696
rect 578000 403600 582820 403696
rect 1104 403056 6000 403152
rect 578000 403056 582820 403152
rect 1104 402512 6000 402608
rect 578000 402512 582820 402608
rect 1104 401968 6000 402064
rect 578000 401968 582820 402064
rect 1104 401424 6000 401520
rect 578000 401424 582820 401520
rect 1104 400880 6000 400976
rect 578000 400880 582820 400976
rect 1104 400336 6000 400432
rect 578000 400336 582820 400432
rect 1104 399792 6000 399888
rect 578000 399792 582820 399888
rect 1104 399248 6000 399344
rect 578000 399248 582820 399344
rect 1104 398704 6000 398800
rect 578000 398704 582820 398800
rect 1104 398160 6000 398256
rect 578000 398160 582820 398256
rect 1104 397616 6000 397712
rect 578000 397616 582820 397712
rect 1104 397072 6000 397168
rect 578000 397072 582820 397168
rect 1104 396528 6000 396624
rect 578000 396528 582820 396624
rect 1104 395984 6000 396080
rect 578000 395984 582820 396080
rect 3234 395700 3240 395752
rect 3292 395740 3298 395752
rect 6730 395740 6736 395752
rect 3292 395712 6736 395740
rect 3292 395700 3298 395712
rect 6730 395700 6736 395712
rect 6788 395700 6794 395752
rect 1104 395440 6000 395536
rect 578000 395440 582820 395536
rect 1104 394896 6000 394992
rect 578000 394896 582820 394992
rect 1104 394352 6000 394448
rect 578000 394352 582820 394448
rect 1104 393808 6000 393904
rect 578000 393808 582820 393904
rect 1104 393264 6000 393360
rect 578000 393264 582820 393360
rect 576670 393184 576676 393236
rect 576728 393224 576734 393236
rect 579614 393224 579620 393236
rect 576728 393196 579620 393224
rect 576728 393184 576734 393196
rect 579614 393184 579620 393196
rect 579672 393184 579678 393236
rect 1104 392720 6000 392816
rect 578000 392720 582820 392816
rect 1104 392176 6000 392272
rect 578000 392176 582820 392272
rect 1104 391632 6000 391728
rect 578000 391632 582820 391728
rect 1104 391088 6000 391184
rect 578000 391088 582820 391184
rect 1104 390544 6000 390640
rect 578000 390544 582820 390640
rect 1104 390000 6000 390096
rect 578000 390000 582820 390096
rect 1104 389456 6000 389552
rect 578000 389456 582820 389552
rect 1104 388912 6000 389008
rect 578000 388912 582820 389008
rect 1104 388368 6000 388464
rect 578000 388368 582820 388464
rect 1104 387824 6000 387920
rect 578000 387824 582820 387920
rect 1104 387280 6000 387376
rect 578000 387280 582820 387376
rect 1104 386736 6000 386832
rect 578000 386736 582820 386832
rect 1104 386192 6000 386288
rect 578000 386192 582820 386288
rect 1104 385648 6000 385744
rect 578000 385648 582820 385744
rect 1104 385104 6000 385200
rect 578000 385104 582820 385200
rect 1104 384560 6000 384656
rect 578000 384560 582820 384656
rect 1104 384016 6000 384112
rect 578000 384016 582820 384112
rect 1104 383472 6000 383568
rect 578000 383472 582820 383568
rect 1104 382928 6000 383024
rect 578000 382928 582820 383024
rect 1104 382384 6000 382480
rect 578000 382384 582820 382480
rect 1104 381840 6000 381936
rect 578000 381840 582820 381936
rect 1104 381296 6000 381392
rect 578000 381296 582820 381392
rect 1104 380752 6000 380848
rect 578000 380752 582820 380848
rect 2774 380604 2780 380656
rect 2832 380644 2838 380656
rect 5166 380644 5172 380656
rect 2832 380616 5172 380644
rect 2832 380604 2838 380616
rect 5166 380604 5172 380616
rect 5224 380604 5230 380656
rect 1104 380208 6000 380304
rect 578000 380208 582820 380304
rect 1104 379664 6000 379760
rect 578000 379664 582820 379760
rect 1104 379120 6000 379216
rect 578000 379120 582820 379216
rect 1104 378576 6000 378672
rect 578000 378576 582820 378672
rect 1104 378032 6000 378128
rect 578000 378032 582820 378128
rect 1104 377488 6000 377584
rect 578000 377488 582820 377584
rect 1104 376944 6000 377040
rect 578000 376944 582820 377040
rect 1104 376400 6000 376496
rect 578000 376400 582820 376496
rect 1104 375856 6000 375952
rect 578000 375856 582820 375952
rect 1104 375312 6000 375408
rect 578000 375312 582820 375408
rect 1104 374768 6000 374864
rect 578000 374768 582820 374864
rect 1104 374224 6000 374320
rect 578000 374224 582820 374320
rect 1104 373680 6000 373776
rect 578000 373680 582820 373776
rect 1104 373136 6000 373232
rect 578000 373136 582820 373232
rect 1104 372592 6000 372688
rect 578000 372592 582820 372688
rect 1104 372048 6000 372144
rect 578000 372048 582820 372144
rect 1104 371504 6000 371600
rect 578000 371504 582820 371600
rect 1104 370960 6000 371056
rect 578000 370960 582820 371056
rect 1104 370416 6000 370512
rect 578000 370416 582820 370512
rect 1104 369872 6000 369968
rect 578000 369872 582820 369968
rect 577774 369792 577780 369844
rect 577832 369832 577838 369844
rect 580718 369832 580724 369844
rect 577832 369804 580724 369832
rect 577832 369792 577838 369804
rect 580718 369792 580724 369804
rect 580776 369792 580782 369844
rect 1104 369328 6000 369424
rect 578000 369328 582820 369424
rect 1104 368784 6000 368880
rect 578000 368784 582820 368880
rect 1104 368240 6000 368336
rect 578000 368240 582820 368336
rect 1104 367696 6000 367792
rect 578000 367696 582820 367792
rect 1104 367152 6000 367248
rect 578000 367152 582820 367248
rect 3234 367004 3240 367056
rect 3292 367044 3298 367056
rect 6638 367044 6644 367056
rect 3292 367016 6644 367044
rect 3292 367004 3298 367016
rect 6638 367004 6644 367016
rect 6696 367004 6702 367056
rect 1104 366608 6000 366704
rect 578000 366608 582820 366704
rect 1104 366064 6000 366160
rect 578000 366064 582820 366160
rect 1104 365520 6000 365616
rect 578000 365520 582820 365616
rect 1104 364976 6000 365072
rect 578000 364976 582820 365072
rect 1104 364432 6000 364528
rect 578000 364432 582820 364528
rect 1104 363888 6000 363984
rect 578000 363888 582820 363984
rect 1104 363344 6000 363440
rect 578000 363344 582820 363440
rect 1104 362800 6000 362896
rect 578000 362800 582820 362896
rect 1104 362256 6000 362352
rect 578000 362256 582820 362352
rect 1104 361712 6000 361808
rect 578000 361712 582820 361808
rect 1104 361168 6000 361264
rect 578000 361168 582820 361264
rect 1104 360624 6000 360720
rect 578000 360624 582820 360720
rect 1104 360080 6000 360176
rect 578000 360080 582820 360176
rect 1104 359536 6000 359632
rect 578000 359536 582820 359632
rect 1104 358992 6000 359088
rect 578000 358992 582820 359088
rect 1104 358448 6000 358544
rect 578000 358448 582820 358544
rect 1104 357904 6000 358000
rect 578000 357904 582820 358000
rect 1104 357360 6000 357456
rect 578000 357360 582820 357456
rect 1104 356816 6000 356912
rect 578000 356816 582820 356912
rect 1104 356272 6000 356368
rect 578000 356272 582820 356368
rect 1104 355728 6000 355824
rect 578000 355728 582820 355824
rect 1104 355184 6000 355280
rect 578000 355184 582820 355280
rect 1104 354640 6000 354736
rect 578000 354640 582820 354736
rect 1104 354096 6000 354192
rect 578000 354096 582820 354192
rect 1104 353552 6000 353648
rect 578000 353552 582820 353648
rect 1104 353008 6000 353104
rect 578000 353008 582820 353104
rect 1104 352464 6000 352560
rect 578000 352464 582820 352560
rect 1104 351920 6000 352016
rect 578000 351920 582820 352016
rect 1104 351376 6000 351472
rect 578000 351376 582820 351472
rect 1104 350832 6000 350928
rect 578000 350832 582820 350928
rect 1104 350288 6000 350384
rect 578000 350288 582820 350384
rect 1104 349744 6000 349840
rect 578000 349744 582820 349840
rect 1104 349200 6000 349296
rect 578000 349200 582820 349296
rect 1104 348656 6000 348752
rect 578000 348656 582820 348752
rect 1104 348112 6000 348208
rect 578000 348112 582820 348208
rect 1104 347568 6000 347664
rect 578000 347568 582820 347664
rect 1104 347024 6000 347120
rect 578000 347024 582820 347120
rect 1104 346480 6000 346576
rect 578000 346480 582820 346576
rect 576578 346332 576584 346384
rect 576636 346372 576642 346384
rect 580166 346372 580172 346384
rect 576636 346344 580172 346372
rect 576636 346332 576642 346344
rect 580166 346332 580172 346344
rect 580224 346332 580230 346384
rect 1104 345936 6000 346032
rect 578000 345936 582820 346032
rect 1104 345392 6000 345488
rect 578000 345392 582820 345488
rect 1104 344848 6000 344944
rect 578000 344848 582820 344944
rect 1104 344304 6000 344400
rect 578000 344304 582820 344400
rect 1104 343760 6000 343856
rect 578000 343760 582820 343856
rect 1104 343216 6000 343312
rect 578000 343216 582820 343312
rect 1104 342672 6000 342768
rect 578000 342672 582820 342768
rect 1104 342128 6000 342224
rect 578000 342128 582820 342224
rect 1104 341584 6000 341680
rect 578000 341584 582820 341680
rect 1104 341040 6000 341136
rect 578000 341040 582820 341136
rect 1104 340496 6000 340592
rect 578000 340496 582820 340592
rect 1104 339952 6000 340048
rect 578000 339952 582820 340048
rect 1104 339408 6000 339504
rect 578000 339408 582820 339504
rect 1104 338864 6000 338960
rect 578000 338864 582820 338960
rect 1104 338320 6000 338416
rect 578000 338320 582820 338416
rect 1104 337776 6000 337872
rect 578000 337776 582820 337872
rect 3234 337628 3240 337680
rect 3292 337668 3298 337680
rect 6546 337668 6552 337680
rect 3292 337640 6552 337668
rect 3292 337628 3298 337640
rect 6546 337628 6552 337640
rect 6604 337628 6610 337680
rect 1104 337232 6000 337328
rect 578000 337232 582820 337328
rect 1104 336688 6000 336784
rect 578000 336688 582820 336784
rect 1104 336144 6000 336240
rect 578000 336144 582820 336240
rect 1104 335600 6000 335696
rect 578000 335600 582820 335696
rect 1104 335056 6000 335152
rect 578000 335056 582820 335152
rect 1104 334512 6000 334608
rect 578000 334512 582820 334608
rect 1104 333968 6000 334064
rect 578000 333968 582820 334064
rect 1104 333424 6000 333520
rect 578000 333424 582820 333520
rect 1104 332880 6000 332976
rect 578000 332880 582820 332976
rect 1104 332336 6000 332432
rect 578000 332336 582820 332432
rect 1104 331792 6000 331888
rect 578000 331792 582820 331888
rect 1104 331248 6000 331344
rect 578000 331248 582820 331344
rect 1104 330704 6000 330800
rect 578000 330704 582820 330800
rect 1104 330160 6000 330256
rect 578000 330160 582820 330256
rect 1104 329616 6000 329712
rect 578000 329616 582820 329712
rect 1104 329072 6000 329168
rect 578000 329072 582820 329168
rect 1104 328528 6000 328624
rect 578000 328528 582820 328624
rect 1104 327984 6000 328080
rect 578000 327984 582820 328080
rect 1104 327440 6000 327536
rect 578000 327440 582820 327536
rect 1104 326896 6000 326992
rect 578000 326896 582820 326992
rect 1104 326352 6000 326448
rect 578000 326352 582820 326448
rect 1104 325808 6000 325904
rect 578000 325808 582820 325904
rect 1104 325264 6000 325360
rect 578000 325264 582820 325360
rect 1104 324720 6000 324816
rect 578000 324720 582820 324816
rect 1104 324176 6000 324272
rect 578000 324176 582820 324272
rect 1104 323632 6000 323728
rect 578000 323632 582820 323728
rect 1104 323088 6000 323184
rect 578000 323088 582820 323184
rect 1104 322544 6000 322640
rect 578000 322544 582820 322640
rect 1104 322000 6000 322096
rect 578000 322000 582820 322096
rect 1104 321456 6000 321552
rect 578000 321456 582820 321552
rect 1104 320912 6000 321008
rect 578000 320912 582820 321008
rect 1104 320368 6000 320464
rect 578000 320368 582820 320464
rect 1104 319824 6000 319920
rect 578000 319824 582820 319920
rect 1104 319280 6000 319376
rect 578000 319280 582820 319376
rect 1104 318736 6000 318832
rect 578000 318736 582820 318832
rect 1104 318192 6000 318288
rect 578000 318192 582820 318288
rect 1104 317648 6000 317744
rect 578000 317648 582820 317744
rect 1104 317104 6000 317200
rect 578000 317104 582820 317200
rect 1104 316560 6000 316656
rect 578000 316560 582820 316656
rect 1104 316016 6000 316112
rect 578000 316016 582820 316112
rect 1104 315472 6000 315568
rect 578000 315472 582820 315568
rect 1104 314928 6000 315024
rect 578000 314928 582820 315024
rect 1104 314384 6000 314480
rect 578000 314384 582820 314480
rect 1104 313840 6000 313936
rect 578000 313840 582820 313936
rect 1104 313296 6000 313392
rect 578000 313296 582820 313392
rect 1104 312752 6000 312848
rect 578000 312752 582820 312848
rect 1104 312208 6000 312304
rect 578000 312208 582820 312304
rect 1104 311664 6000 311760
rect 578000 311664 582820 311760
rect 1104 311120 6000 311216
rect 578000 311120 582820 311216
rect 1104 310576 6000 310672
rect 578000 310576 582820 310672
rect 1104 310032 6000 310128
rect 578000 310032 582820 310128
rect 1104 309488 6000 309584
rect 578000 309488 582820 309584
rect 1104 308944 6000 309040
rect 578000 308944 582820 309040
rect 3234 308864 3240 308916
rect 3292 308904 3298 308916
rect 8110 308904 8116 308916
rect 3292 308876 8116 308904
rect 3292 308864 3298 308876
rect 8110 308864 8116 308876
rect 8168 308864 8174 308916
rect 1104 308400 6000 308496
rect 578000 308400 582820 308496
rect 1104 307856 6000 307952
rect 578000 307856 582820 307952
rect 1104 307312 6000 307408
rect 578000 307312 582820 307408
rect 1104 306768 6000 306864
rect 578000 306768 582820 306864
rect 1104 306224 6000 306320
rect 578000 306224 582820 306320
rect 1104 305680 6000 305776
rect 578000 305680 582820 305776
rect 1104 305136 6000 305232
rect 578000 305136 582820 305232
rect 1104 304592 6000 304688
rect 578000 304592 582820 304688
rect 1104 304048 6000 304144
rect 578000 304048 582820 304144
rect 1104 303504 6000 303600
rect 578000 303504 582820 303600
rect 1104 302960 6000 303056
rect 578000 302960 582820 303056
rect 1104 302416 6000 302512
rect 578000 302416 582820 302512
rect 1104 301872 6000 301968
rect 578000 301872 582820 301968
rect 1104 301328 6000 301424
rect 578000 301328 582820 301424
rect 1104 300784 6000 300880
rect 578000 300784 582820 300880
rect 1104 300240 6000 300336
rect 578000 300240 582820 300336
rect 1104 299696 6000 299792
rect 578000 299696 582820 299792
rect 576486 299412 576492 299464
rect 576544 299452 576550 299464
rect 580166 299452 580172 299464
rect 576544 299424 580172 299452
rect 576544 299412 576550 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 1104 299152 6000 299248
rect 578000 299152 582820 299248
rect 1104 298608 6000 298704
rect 578000 298608 582820 298704
rect 1104 298064 6000 298160
rect 578000 298064 582820 298160
rect 1104 297520 6000 297616
rect 578000 297520 582820 297616
rect 1104 296976 6000 297072
rect 578000 296976 582820 297072
rect 1104 296432 6000 296528
rect 578000 296432 582820 296528
rect 1104 295888 6000 295984
rect 578000 295888 582820 295984
rect 1104 295344 6000 295440
rect 578000 295344 582820 295440
rect 1104 294800 6000 294896
rect 578000 294800 582820 294896
rect 3234 294720 3240 294772
rect 3292 294760 3298 294772
rect 6454 294760 6460 294772
rect 3292 294732 6460 294760
rect 3292 294720 3298 294732
rect 6454 294720 6460 294732
rect 6512 294720 6518 294772
rect 1104 294256 6000 294352
rect 578000 294256 582820 294352
rect 1104 293712 6000 293808
rect 578000 293712 582820 293808
rect 1104 293168 6000 293264
rect 578000 293168 582820 293264
rect 1104 292624 6000 292720
rect 578000 292624 582820 292720
rect 1104 292080 6000 292176
rect 578000 292080 582820 292176
rect 1104 291536 6000 291632
rect 578000 291536 582820 291632
rect 1104 290992 6000 291088
rect 578000 290992 582820 291088
rect 1104 290448 6000 290544
rect 578000 290448 582820 290544
rect 1104 289904 6000 290000
rect 578000 289904 582820 290000
rect 1104 289360 6000 289456
rect 578000 289360 582820 289456
rect 1104 288816 6000 288912
rect 578000 288816 582820 288912
rect 1104 288272 6000 288368
rect 578000 288272 582820 288368
rect 1104 287728 6000 287824
rect 578000 287728 582820 287824
rect 1104 287184 6000 287280
rect 578000 287184 582820 287280
rect 1104 286640 6000 286736
rect 578000 286640 582820 286736
rect 1104 286096 6000 286192
rect 578000 286096 582820 286192
rect 1104 285552 6000 285648
rect 578000 285552 582820 285648
rect 1104 285008 6000 285104
rect 578000 285008 582820 285104
rect 1104 284464 6000 284560
rect 578000 284464 582820 284560
rect 1104 283920 6000 284016
rect 578000 283920 582820 284016
rect 1104 283376 6000 283472
rect 578000 283376 582820 283472
rect 1104 282832 6000 282928
rect 578000 282832 582820 282928
rect 1104 282288 6000 282384
rect 578000 282288 582820 282384
rect 1104 281744 6000 281840
rect 578000 281744 582820 281840
rect 1104 281200 6000 281296
rect 578000 281200 582820 281296
rect 1104 280656 6000 280752
rect 578000 280656 582820 280752
rect 1104 280112 6000 280208
rect 578000 280112 582820 280208
rect 2774 280032 2780 280084
rect 2832 280072 2838 280084
rect 5074 280072 5080 280084
rect 2832 280044 5080 280072
rect 2832 280032 2838 280044
rect 5074 280032 5080 280044
rect 5132 280032 5138 280084
rect 1104 279568 6000 279664
rect 578000 279568 582820 279664
rect 1104 279024 6000 279120
rect 578000 279024 582820 279120
rect 1104 278480 6000 278576
rect 578000 278480 582820 278576
rect 1104 277936 6000 278032
rect 578000 277936 582820 278032
rect 1104 277392 6000 277488
rect 578000 277392 582820 277488
rect 1104 276848 6000 276944
rect 578000 276848 582820 276944
rect 1104 276304 6000 276400
rect 578000 276304 582820 276400
rect 577682 275952 577688 276004
rect 577740 275992 577746 276004
rect 579614 275992 579620 276004
rect 577740 275964 579620 275992
rect 577740 275952 577746 275964
rect 579614 275952 579620 275964
rect 579672 275952 579678 276004
rect 1104 275760 6000 275856
rect 578000 275760 582820 275856
rect 1104 275216 6000 275312
rect 578000 275216 582820 275312
rect 1104 274672 6000 274768
rect 578000 274672 582820 274768
rect 1104 274128 6000 274224
rect 578000 274128 582820 274224
rect 1104 273584 6000 273680
rect 578000 273584 582820 273680
rect 1104 273040 6000 273136
rect 578000 273040 582820 273136
rect 1104 272496 6000 272592
rect 578000 272496 582820 272592
rect 1104 271952 6000 272048
rect 578000 271952 582820 272048
rect 1104 271408 6000 271504
rect 578000 271408 582820 271504
rect 1104 270864 6000 270960
rect 578000 270864 582820 270960
rect 1104 270320 6000 270416
rect 578000 270320 582820 270416
rect 1104 269776 6000 269872
rect 578000 269776 582820 269872
rect 1104 269232 6000 269328
rect 578000 269232 582820 269328
rect 1104 268688 6000 268784
rect 578000 268688 582820 268784
rect 1104 268144 6000 268240
rect 578000 268144 582820 268240
rect 1104 267600 6000 267696
rect 578000 267600 582820 267696
rect 1104 267056 6000 267152
rect 578000 267056 582820 267152
rect 1104 266512 6000 266608
rect 578000 266512 582820 266608
rect 2958 266296 2964 266348
rect 3016 266336 3022 266348
rect 6362 266336 6368 266348
rect 3016 266308 6368 266336
rect 3016 266296 3022 266308
rect 6362 266296 6368 266308
rect 6420 266296 6426 266348
rect 1104 265968 6000 266064
rect 578000 265968 582820 266064
rect 1104 265424 6000 265520
rect 578000 265424 582820 265520
rect 1104 264880 6000 264976
rect 578000 264880 582820 264976
rect 1104 264336 6000 264432
rect 578000 264336 582820 264432
rect 1104 263792 6000 263888
rect 578000 263792 582820 263888
rect 1104 263248 6000 263344
rect 578000 263248 582820 263344
rect 1104 262704 6000 262800
rect 578000 262704 582820 262800
rect 1104 262160 6000 262256
rect 578000 262160 582820 262256
rect 1104 261616 6000 261712
rect 578000 261616 582820 261712
rect 1104 261072 6000 261168
rect 578000 261072 582820 261168
rect 1104 260528 6000 260624
rect 578000 260528 582820 260624
rect 1104 259984 6000 260080
rect 578000 259984 582820 260080
rect 1104 259440 6000 259536
rect 578000 259440 582820 259536
rect 1104 258896 6000 258992
rect 578000 258896 582820 258992
rect 1104 258352 6000 258448
rect 578000 258352 582820 258448
rect 1104 257808 6000 257904
rect 578000 257808 582820 257904
rect 1104 257264 6000 257360
rect 578000 257264 582820 257360
rect 1104 256720 6000 256816
rect 578000 256720 582820 256816
rect 1104 256176 6000 256272
rect 578000 256176 582820 256272
rect 1104 255632 6000 255728
rect 578000 255632 582820 255728
rect 1104 255088 6000 255184
rect 578000 255088 582820 255184
rect 1104 254544 6000 254640
rect 578000 254544 582820 254640
rect 1104 254000 6000 254096
rect 578000 254000 582820 254096
rect 1104 253456 6000 253552
rect 578000 253456 582820 253552
rect 1104 252912 6000 253008
rect 578000 252912 582820 253008
rect 3234 252492 3240 252544
rect 3292 252532 3298 252544
rect 6270 252532 6276 252544
rect 3292 252504 6276 252532
rect 3292 252492 3298 252504
rect 6270 252492 6276 252504
rect 6328 252492 6334 252544
rect 576394 252492 576400 252544
rect 576452 252532 576458 252544
rect 580166 252532 580172 252544
rect 576452 252504 580172 252532
rect 576452 252492 576458 252504
rect 580166 252492 580172 252504
rect 580224 252492 580230 252544
rect 1104 252368 6000 252464
rect 578000 252368 582820 252464
rect 1104 251824 6000 251920
rect 578000 251824 582820 251920
rect 1104 251280 6000 251376
rect 578000 251280 582820 251376
rect 1104 250736 6000 250832
rect 578000 250736 582820 250832
rect 1104 250192 6000 250288
rect 578000 250192 582820 250288
rect 1104 249648 6000 249744
rect 578000 249648 582820 249744
rect 1104 249104 6000 249200
rect 578000 249104 582820 249200
rect 1104 248560 6000 248656
rect 578000 248560 582820 248656
rect 1104 248016 6000 248112
rect 578000 248016 582820 248112
rect 1104 247472 6000 247568
rect 578000 247472 582820 247568
rect 1104 246928 6000 247024
rect 578000 246928 582820 247024
rect 1104 246384 6000 246480
rect 578000 246384 582820 246480
rect 1104 245840 6000 245936
rect 578000 245840 582820 245936
rect 1104 245296 6000 245392
rect 578000 245296 582820 245392
rect 1104 244752 6000 244848
rect 578000 244752 582820 244848
rect 1104 244208 6000 244304
rect 578000 244208 582820 244304
rect 1104 243664 6000 243760
rect 578000 243664 582820 243760
rect 1104 243120 6000 243216
rect 578000 243120 582820 243216
rect 1104 242576 6000 242672
rect 578000 242576 582820 242672
rect 1104 242032 6000 242128
rect 578000 242032 582820 242128
rect 1104 241488 6000 241584
rect 578000 241488 582820 241584
rect 1104 240944 6000 241040
rect 578000 240944 582820 241040
rect 1104 240400 6000 240496
rect 578000 240400 582820 240496
rect 1104 239856 6000 239952
rect 578000 239856 582820 239952
rect 1104 239312 6000 239408
rect 578000 239312 582820 239408
rect 1104 238768 6000 238864
rect 578000 238768 582820 238864
rect 1104 238224 6000 238320
rect 578000 238224 582820 238320
rect 1104 237680 6000 237776
rect 578000 237680 582820 237776
rect 1104 237136 6000 237232
rect 578000 237136 582820 237232
rect 1104 236592 6000 236688
rect 578000 236592 582820 236688
rect 1104 236048 6000 236144
rect 578000 236048 582820 236144
rect 1104 235504 6000 235600
rect 578000 235504 582820 235600
rect 1104 234960 6000 235056
rect 578000 234960 582820 235056
rect 1104 234416 6000 234512
rect 578000 234416 582820 234512
rect 1104 233872 6000 233968
rect 578000 233872 582820 233968
rect 1104 233328 6000 233424
rect 578000 233328 582820 233424
rect 1104 232784 6000 232880
rect 578000 232784 582820 232880
rect 1104 232240 6000 232336
rect 578000 232240 582820 232336
rect 1104 231696 6000 231792
rect 578000 231696 582820 231792
rect 1104 231152 6000 231248
rect 578000 231152 582820 231248
rect 1104 230608 6000 230704
rect 578000 230608 582820 230704
rect 1104 230064 6000 230160
rect 578000 230064 582820 230160
rect 1104 229520 6000 229616
rect 578000 229520 582820 229616
rect 1104 228976 6000 229072
rect 578000 228976 582820 229072
rect 1104 228432 6000 228528
rect 578000 228432 582820 228528
rect 1104 227888 6000 227984
rect 578000 227888 582820 227984
rect 1104 227344 6000 227440
rect 578000 227344 582820 227440
rect 1104 226800 6000 226896
rect 578000 226800 582820 226896
rect 1104 226256 6000 226352
rect 578000 226256 582820 226352
rect 1104 225712 6000 225808
rect 578000 225712 582820 225808
rect 1104 225168 6000 225264
rect 578000 225168 582820 225264
rect 1104 224624 6000 224720
rect 578000 224624 582820 224720
rect 1104 224080 6000 224176
rect 578000 224080 582820 224176
rect 1104 223536 6000 223632
rect 578000 223536 582820 223632
rect 1104 222992 6000 223088
rect 578000 222992 582820 223088
rect 1104 222448 6000 222544
rect 578000 222448 582820 222544
rect 1104 221904 6000 222000
rect 578000 221904 582820 222000
rect 1104 221360 6000 221456
rect 578000 221360 582820 221456
rect 1104 220816 6000 220912
rect 578000 220816 582820 220912
rect 1104 220272 6000 220368
rect 578000 220272 582820 220368
rect 1104 219728 6000 219824
rect 578000 219728 582820 219824
rect 1104 219184 6000 219280
rect 578000 219184 582820 219280
rect 1104 218640 6000 218736
rect 578000 218640 582820 218736
rect 1104 218096 6000 218192
rect 578000 218096 582820 218192
rect 1104 217552 6000 217648
rect 578000 217552 582820 217648
rect 1104 217008 6000 217104
rect 578000 217008 582820 217104
rect 1104 216464 6000 216560
rect 578000 216464 582820 216560
rect 1104 215920 6000 216016
rect 578000 215920 582820 216016
rect 1104 215376 6000 215472
rect 578000 215376 582820 215472
rect 1104 214832 6000 214928
rect 578000 214832 582820 214928
rect 1104 214288 6000 214384
rect 578000 214288 582820 214384
rect 1104 213744 6000 213840
rect 578000 213744 582820 213840
rect 1104 213200 6000 213296
rect 578000 213200 582820 213296
rect 1104 212656 6000 212752
rect 578000 212656 582820 212752
rect 1104 212112 6000 212208
rect 578000 212112 582820 212208
rect 1104 211568 6000 211664
rect 578000 211568 582820 211664
rect 1104 211024 6000 211120
rect 578000 211024 582820 211120
rect 1104 210480 6000 210576
rect 578000 210480 582820 210576
rect 1104 209936 6000 210032
rect 578000 209936 582820 210032
rect 1104 209392 6000 209488
rect 578000 209392 582820 209488
rect 1104 208848 6000 208944
rect 578000 208848 582820 208944
rect 1104 208304 6000 208400
rect 578000 208304 582820 208400
rect 3326 208156 3332 208208
rect 3384 208196 3390 208208
rect 8018 208196 8024 208208
rect 3384 208168 8024 208196
rect 3384 208156 3390 208168
rect 8018 208156 8024 208168
rect 8076 208156 8082 208208
rect 1104 207760 6000 207856
rect 578000 207760 582820 207856
rect 1104 207216 6000 207312
rect 578000 207216 582820 207312
rect 1104 206672 6000 206768
rect 578000 206672 582820 206768
rect 1104 206128 6000 206224
rect 578000 206128 582820 206224
rect 1104 205584 6000 205680
rect 578000 205584 582820 205680
rect 575106 205504 575112 205556
rect 575164 205544 575170 205556
rect 580166 205544 580172 205556
rect 575164 205516 580172 205544
rect 575164 205504 575170 205516
rect 580166 205504 580172 205516
rect 580224 205504 580230 205556
rect 1104 205040 6000 205136
rect 578000 205040 582820 205136
rect 1104 204496 6000 204592
rect 578000 204496 582820 204592
rect 1104 203952 6000 204048
rect 578000 203952 582820 204048
rect 1104 203408 6000 203504
rect 578000 203408 582820 203504
rect 1104 202864 6000 202960
rect 578000 202864 582820 202960
rect 1104 202320 6000 202416
rect 578000 202320 582820 202416
rect 1104 201776 6000 201872
rect 578000 201776 582820 201872
rect 1104 201232 6000 201328
rect 578000 201232 582820 201328
rect 1104 200688 6000 200784
rect 578000 200688 582820 200784
rect 1104 200144 6000 200240
rect 578000 200144 582820 200240
rect 1104 199600 6000 199696
rect 578000 199600 582820 199696
rect 1104 199056 6000 199152
rect 578000 199056 582820 199152
rect 1104 198512 6000 198608
rect 578000 198512 582820 198608
rect 1104 197968 6000 198064
rect 578000 197968 582820 198064
rect 1104 197424 6000 197520
rect 578000 197424 582820 197520
rect 1104 196880 6000 196976
rect 578000 196880 582820 196976
rect 1104 196336 6000 196432
rect 578000 196336 582820 196432
rect 1104 195792 6000 195888
rect 578000 195792 582820 195888
rect 1104 195248 6000 195344
rect 578000 195248 582820 195344
rect 1104 194704 6000 194800
rect 578000 194704 582820 194800
rect 2774 194420 2780 194472
rect 2832 194460 2838 194472
rect 4890 194460 4896 194472
rect 2832 194432 4896 194460
rect 2832 194420 2838 194432
rect 4890 194420 4896 194432
rect 4948 194420 4954 194472
rect 1104 194160 6000 194256
rect 578000 194160 582820 194256
rect 1104 193616 6000 193712
rect 578000 193616 582820 193712
rect 1104 193072 6000 193168
rect 578000 193072 582820 193168
rect 1104 192528 6000 192624
rect 578000 192528 582820 192624
rect 1104 191984 6000 192080
rect 578000 191984 582820 192080
rect 1104 191440 6000 191536
rect 578000 191440 582820 191536
rect 1104 190896 6000 190992
rect 578000 190896 582820 190992
rect 1104 190352 6000 190448
rect 578000 190352 582820 190448
rect 1104 189808 6000 189904
rect 578000 189808 582820 189904
rect 1104 189264 6000 189360
rect 578000 189264 582820 189360
rect 1104 188720 6000 188816
rect 578000 188720 582820 188816
rect 1104 188176 6000 188272
rect 578000 188176 582820 188272
rect 1104 187632 6000 187728
rect 578000 187632 582820 187728
rect 1104 187088 6000 187184
rect 578000 187088 582820 187184
rect 1104 186544 6000 186640
rect 578000 186544 582820 186640
rect 1104 186000 6000 186096
rect 578000 186000 582820 186096
rect 1104 185456 6000 185552
rect 578000 185456 582820 185552
rect 1104 184912 6000 185008
rect 578000 184912 582820 185008
rect 1104 184368 6000 184464
rect 578000 184368 582820 184464
rect 1104 183824 6000 183920
rect 578000 183824 582820 183920
rect 1104 183280 6000 183376
rect 578000 183280 582820 183376
rect 1104 182736 6000 182832
rect 578000 182736 582820 182832
rect 1104 182192 6000 182288
rect 578000 182192 582820 182288
rect 1104 181648 6000 181744
rect 578000 181648 582820 181744
rect 1104 181104 6000 181200
rect 578000 181104 582820 181200
rect 1104 180560 6000 180656
rect 578000 180560 582820 180656
rect 1104 180016 6000 180112
rect 578000 180016 582820 180112
rect 1104 179472 6000 179568
rect 578000 179472 582820 179568
rect 1104 178928 6000 179024
rect 578000 178928 582820 179024
rect 1104 178384 6000 178480
rect 578000 178384 582820 178480
rect 1104 177840 6000 177936
rect 578000 177840 582820 177936
rect 1104 177296 6000 177392
rect 578000 177296 582820 177392
rect 1104 176752 6000 176848
rect 578000 176752 582820 176848
rect 1104 176208 6000 176304
rect 578000 176208 582820 176304
rect 1104 175664 6000 175760
rect 578000 175664 582820 175760
rect 1104 175120 6000 175216
rect 578000 175120 582820 175216
rect 1104 174576 6000 174672
rect 578000 174576 582820 174672
rect 1104 174032 6000 174128
rect 578000 174032 582820 174128
rect 1104 173488 6000 173584
rect 578000 173488 582820 173584
rect 1104 172944 6000 173040
rect 578000 172944 582820 173040
rect 1104 172400 6000 172496
rect 578000 172400 582820 172496
rect 1104 171856 6000 171952
rect 578000 171856 582820 171952
rect 1104 171312 6000 171408
rect 578000 171312 582820 171408
rect 1104 170768 6000 170864
rect 578000 170768 582820 170864
rect 577590 170620 577596 170672
rect 577648 170660 577654 170672
rect 580626 170660 580632 170672
rect 577648 170632 580632 170660
rect 577648 170620 577654 170632
rect 580626 170620 580632 170632
rect 580684 170620 580690 170672
rect 1104 170224 6000 170320
rect 578000 170224 582820 170320
rect 1104 169680 6000 169776
rect 578000 169680 582820 169776
rect 1104 169136 6000 169232
rect 578000 169136 582820 169232
rect 1104 168592 6000 168688
rect 578000 168592 582820 168688
rect 1104 168048 6000 168144
rect 578000 168048 582820 168144
rect 1104 167504 6000 167600
rect 578000 167504 582820 167600
rect 1104 166960 6000 167056
rect 578000 166960 582820 167056
rect 1104 166416 6000 166512
rect 578000 166416 582820 166512
rect 1104 165872 6000 165968
rect 578000 165872 582820 165968
rect 1104 165328 6000 165424
rect 578000 165328 582820 165424
rect 3326 165044 3332 165096
rect 3384 165084 3390 165096
rect 7926 165084 7932 165096
rect 3384 165056 7932 165084
rect 3384 165044 3390 165056
rect 7926 165044 7932 165056
rect 7984 165044 7990 165096
rect 1104 164784 6000 164880
rect 578000 164784 582820 164880
rect 1104 164240 6000 164336
rect 578000 164240 582820 164336
rect 1104 163696 6000 163792
rect 578000 163696 582820 163792
rect 1104 163152 6000 163248
rect 578000 163152 582820 163248
rect 1104 162608 6000 162704
rect 578000 162608 582820 162704
rect 1104 162064 6000 162160
rect 578000 162064 582820 162160
rect 1104 161520 6000 161616
rect 578000 161520 582820 161616
rect 1104 160976 6000 161072
rect 578000 160976 582820 161072
rect 1104 160432 6000 160528
rect 578000 160432 582820 160528
rect 1104 159888 6000 159984
rect 578000 159888 582820 159984
rect 1104 159344 6000 159440
rect 578000 159344 582820 159440
rect 1104 158800 6000 158896
rect 578000 158800 582820 158896
rect 575014 158652 575020 158704
rect 575072 158692 575078 158704
rect 579614 158692 579620 158704
rect 575072 158664 579620 158692
rect 575072 158652 575078 158664
rect 579614 158652 579620 158664
rect 579672 158652 579678 158704
rect 1104 158256 6000 158352
rect 578000 158256 582820 158352
rect 1104 157712 6000 157808
rect 578000 157712 582820 157808
rect 1104 157168 6000 157264
rect 578000 157168 582820 157264
rect 1104 156624 6000 156720
rect 578000 156624 582820 156720
rect 1104 156080 6000 156176
rect 578000 156080 582820 156176
rect 1104 155536 6000 155632
rect 578000 155536 582820 155632
rect 1104 154992 6000 155088
rect 578000 154992 582820 155088
rect 1104 154448 6000 154544
rect 578000 154448 582820 154544
rect 1104 153904 6000 154000
rect 578000 153904 582820 154000
rect 1104 153360 6000 153456
rect 578000 153360 582820 153456
rect 1104 152816 6000 152912
rect 578000 152816 582820 152912
rect 1104 152272 6000 152368
rect 578000 152272 582820 152368
rect 1104 151728 6000 151824
rect 578000 151728 582820 151824
rect 1104 151184 6000 151280
rect 578000 151184 582820 151280
rect 1104 150640 6000 150736
rect 578000 150640 582820 150736
rect 1104 150096 6000 150192
rect 578000 150096 582820 150192
rect 1104 149552 6000 149648
rect 578000 149552 582820 149648
rect 1104 149008 6000 149104
rect 578000 149008 582820 149104
rect 1104 148464 6000 148560
rect 578000 148464 582820 148560
rect 1104 147920 6000 148016
rect 578000 147920 582820 148016
rect 1104 147376 6000 147472
rect 578000 147376 582820 147472
rect 1104 146832 6000 146928
rect 578000 146832 582820 146928
rect 1104 146288 6000 146384
rect 578000 146288 582820 146384
rect 1104 145744 6000 145840
rect 578000 145744 582820 145840
rect 1104 145200 6000 145296
rect 578000 145200 582820 145296
rect 1104 144656 6000 144752
rect 578000 144656 582820 144752
rect 1104 144112 6000 144208
rect 578000 144112 582820 144208
rect 1104 143568 6000 143664
rect 578000 143568 582820 143664
rect 1104 143024 6000 143120
rect 578000 143024 582820 143120
rect 1104 142480 6000 142576
rect 578000 142480 582820 142576
rect 1104 141936 6000 142032
rect 578000 141936 582820 142032
rect 1104 141392 6000 141488
rect 578000 141392 582820 141488
rect 1104 140848 6000 140944
rect 578000 140848 582820 140944
rect 1104 140304 6000 140400
rect 578000 140304 582820 140400
rect 1104 139760 6000 139856
rect 578000 139760 582820 139856
rect 1104 139216 6000 139312
rect 578000 139216 582820 139312
rect 1104 138672 6000 138768
rect 578000 138672 582820 138768
rect 1104 138128 6000 138224
rect 578000 138128 582820 138224
rect 1104 137584 6000 137680
rect 578000 137584 582820 137680
rect 1104 137040 6000 137136
rect 578000 137040 582820 137136
rect 1104 136496 6000 136592
rect 578000 136496 582820 136592
rect 3326 136348 3332 136400
rect 3384 136388 3390 136400
rect 7834 136388 7840 136400
rect 3384 136360 7840 136388
rect 3384 136348 3390 136360
rect 7834 136348 7840 136360
rect 7892 136348 7898 136400
rect 1104 135952 6000 136048
rect 578000 135952 582820 136048
rect 1104 135408 6000 135504
rect 578000 135408 582820 135504
rect 576302 135192 576308 135244
rect 576360 135232 576366 135244
rect 580166 135232 580172 135244
rect 576360 135204 580172 135232
rect 576360 135192 576366 135204
rect 580166 135192 580172 135204
rect 580224 135192 580230 135244
rect 1104 134864 6000 134960
rect 578000 134864 582820 134960
rect 1104 134320 6000 134416
rect 578000 134320 582820 134416
rect 1104 133776 6000 133872
rect 578000 133776 582820 133872
rect 1104 133232 6000 133328
rect 578000 133232 582820 133328
rect 1104 132688 6000 132784
rect 578000 132688 582820 132784
rect 1104 132144 6000 132240
rect 578000 132144 582820 132240
rect 1104 131600 6000 131696
rect 578000 131600 582820 131696
rect 1104 131056 6000 131152
rect 578000 131056 582820 131152
rect 1104 130512 6000 130608
rect 578000 130512 582820 130608
rect 1104 129968 6000 130064
rect 578000 129968 582820 130064
rect 1104 129424 6000 129520
rect 578000 129424 582820 129520
rect 1104 128880 6000 128976
rect 578000 128880 582820 128976
rect 1104 128336 6000 128432
rect 578000 128336 582820 128432
rect 1104 127792 6000 127888
rect 578000 127792 582820 127888
rect 1104 127248 6000 127344
rect 578000 127248 582820 127344
rect 1104 126704 6000 126800
rect 578000 126704 582820 126800
rect 1104 126160 6000 126256
rect 578000 126160 582820 126256
rect 1104 125616 6000 125712
rect 578000 125616 582820 125712
rect 1104 125072 6000 125168
rect 578000 125072 582820 125168
rect 1104 124528 6000 124624
rect 578000 124528 582820 124624
rect 1104 123984 6000 124080
rect 578000 123984 582820 124080
rect 1104 123440 6000 123536
rect 578000 123440 582820 123536
rect 1104 122896 6000 122992
rect 578000 122896 582820 122992
rect 1104 122352 6000 122448
rect 578000 122352 582820 122448
rect 3326 122136 3332 122188
rect 3384 122176 3390 122188
rect 7742 122176 7748 122188
rect 3384 122148 7748 122176
rect 3384 122136 3390 122148
rect 7742 122136 7748 122148
rect 7800 122136 7806 122188
rect 1104 121808 6000 121904
rect 578000 121808 582820 121904
rect 1104 121264 6000 121360
rect 578000 121264 582820 121360
rect 1104 120720 6000 120816
rect 578000 120720 582820 120816
rect 1104 120176 6000 120272
rect 578000 120176 582820 120272
rect 1104 119632 6000 119728
rect 578000 119632 582820 119728
rect 1104 119088 6000 119184
rect 578000 119088 582820 119184
rect 1104 118544 6000 118640
rect 578000 118544 582820 118640
rect 1104 118000 6000 118096
rect 578000 118000 582820 118096
rect 1104 117456 6000 117552
rect 578000 117456 582820 117552
rect 1104 116912 6000 117008
rect 578000 116912 582820 117008
rect 1104 116368 6000 116464
rect 578000 116368 582820 116464
rect 1104 115824 6000 115920
rect 578000 115824 582820 115920
rect 1104 115280 6000 115376
rect 578000 115280 582820 115376
rect 1104 114736 6000 114832
rect 578000 114736 582820 114832
rect 1104 114192 6000 114288
rect 578000 114192 582820 114288
rect 1104 113648 6000 113744
rect 578000 113648 582820 113744
rect 1104 113104 6000 113200
rect 578000 113104 582820 113200
rect 1104 112560 6000 112656
rect 578000 112560 582820 112656
rect 1104 112016 6000 112112
rect 578000 112016 582820 112112
rect 574922 111732 574928 111784
rect 574980 111772 574986 111784
rect 580166 111772 580172 111784
rect 574980 111744 580172 111772
rect 574980 111732 574986 111744
rect 580166 111732 580172 111744
rect 580224 111732 580230 111784
rect 1104 111472 6000 111568
rect 578000 111472 582820 111568
rect 1104 110928 6000 111024
rect 578000 110928 582820 111024
rect 1104 110384 6000 110480
rect 578000 110384 582820 110480
rect 1104 109840 6000 109936
rect 578000 109840 582820 109936
rect 1104 109296 6000 109392
rect 578000 109296 582820 109392
rect 1104 108752 6000 108848
rect 578000 108752 582820 108848
rect 1104 108208 6000 108304
rect 578000 108208 582820 108304
rect 2774 107992 2780 108044
rect 2832 108032 2838 108044
rect 4982 108032 4988 108044
rect 2832 108004 4988 108032
rect 2832 107992 2838 108004
rect 4982 107992 4988 108004
rect 5040 107992 5046 108044
rect 1104 107664 6000 107760
rect 578000 107664 582820 107760
rect 1104 107120 6000 107216
rect 578000 107120 582820 107216
rect 1104 106576 6000 106672
rect 578000 106576 582820 106672
rect 1104 106032 6000 106128
rect 578000 106032 582820 106128
rect 1104 105488 6000 105584
rect 578000 105488 582820 105584
rect 1104 104944 6000 105040
rect 578000 104944 582820 105040
rect 1104 104400 6000 104496
rect 578000 104400 582820 104496
rect 1104 103856 6000 103952
rect 578000 103856 582820 103952
rect 1104 103312 6000 103408
rect 578000 103312 582820 103408
rect 1104 102768 6000 102864
rect 578000 102768 582820 102864
rect 1104 102224 6000 102320
rect 578000 102224 582820 102320
rect 1104 101680 6000 101776
rect 578000 101680 582820 101776
rect 1104 101136 6000 101232
rect 578000 101136 582820 101232
rect 1104 100592 6000 100688
rect 578000 100592 582820 100688
rect 1104 100048 6000 100144
rect 578000 100048 582820 100144
rect 1104 99504 6000 99600
rect 578000 99504 582820 99600
rect 1104 98960 6000 99056
rect 578000 98960 582820 99056
rect 1104 98416 6000 98512
rect 578000 98416 582820 98512
rect 1104 97872 6000 97968
rect 578000 97872 582820 97968
rect 1104 97328 6000 97424
rect 578000 97328 582820 97424
rect 1104 96784 6000 96880
rect 578000 96784 582820 96880
rect 1104 96240 6000 96336
rect 578000 96240 582820 96336
rect 1104 95696 6000 95792
rect 578000 95696 582820 95792
rect 1104 95152 6000 95248
rect 578000 95152 582820 95248
rect 1104 94608 6000 94704
rect 578000 94608 582820 94704
rect 1104 94064 6000 94160
rect 578000 94064 582820 94160
rect 1104 93520 6000 93616
rect 578000 93520 582820 93616
rect 1104 92976 6000 93072
rect 578000 92976 582820 93072
rect 1104 92432 6000 92528
rect 578000 92432 582820 92528
rect 1104 91888 6000 91984
rect 578000 91888 582820 91984
rect 1104 91344 6000 91440
rect 578000 91344 582820 91440
rect 1104 90800 6000 90896
rect 578000 90800 582820 90896
rect 1104 90256 6000 90352
rect 578000 90256 582820 90352
rect 1104 89712 6000 89808
rect 578000 89712 582820 89808
rect 1104 89168 6000 89264
rect 578000 89168 582820 89264
rect 1104 88624 6000 88720
rect 578000 88624 582820 88720
rect 576210 88272 576216 88324
rect 576268 88312 576274 88324
rect 579890 88312 579896 88324
rect 576268 88284 579896 88312
rect 576268 88272 576274 88284
rect 579890 88272 579896 88284
rect 579948 88272 579954 88324
rect 1104 88080 6000 88176
rect 578000 88080 582820 88176
rect 1104 87536 6000 87632
rect 578000 87536 582820 87632
rect 1104 86992 6000 87088
rect 578000 86992 582820 87088
rect 1104 86448 6000 86544
rect 578000 86448 582820 86544
rect 1104 85904 6000 86000
rect 578000 85904 582820 86000
rect 1104 85360 6000 85456
rect 578000 85360 582820 85456
rect 1104 84816 6000 84912
rect 578000 84816 582820 84912
rect 1104 84272 6000 84368
rect 578000 84272 582820 84368
rect 1104 83728 6000 83824
rect 578000 83728 582820 83824
rect 1104 83184 6000 83280
rect 578000 83184 582820 83280
rect 1104 82640 6000 82736
rect 578000 82640 582820 82736
rect 1104 82096 6000 82192
rect 578000 82096 582820 82192
rect 1104 81552 6000 81648
rect 578000 81552 582820 81648
rect 1104 81008 6000 81104
rect 578000 81008 582820 81104
rect 1104 80464 6000 80560
rect 578000 80464 582820 80560
rect 1104 79920 6000 80016
rect 578000 79920 582820 80016
rect 3050 79840 3056 79892
rect 3108 79880 3114 79892
rect 7650 79880 7656 79892
rect 3108 79852 7656 79880
rect 3108 79840 3114 79852
rect 7650 79840 7656 79852
rect 7708 79840 7714 79892
rect 1104 79376 6000 79472
rect 578000 79376 582820 79472
rect 1104 78832 6000 78928
rect 578000 78832 582820 78928
rect 1104 78288 6000 78384
rect 578000 78288 582820 78384
rect 1104 77744 6000 77840
rect 578000 77744 582820 77840
rect 1104 77200 6000 77296
rect 578000 77200 582820 77296
rect 1104 76656 6000 76752
rect 578000 76656 582820 76752
rect 1104 76112 6000 76208
rect 578000 76112 582820 76208
rect 1104 75568 6000 75664
rect 578000 75568 582820 75664
rect 1104 75024 6000 75120
rect 578000 75024 582820 75120
rect 1104 74480 6000 74576
rect 578000 74480 582820 74576
rect 1104 73936 6000 74032
rect 578000 73936 582820 74032
rect 1104 73392 6000 73488
rect 578000 73392 582820 73488
rect 1104 72848 6000 72944
rect 578000 72848 582820 72944
rect 1104 72304 6000 72400
rect 578000 72304 582820 72400
rect 1104 71760 6000 71856
rect 578000 71760 582820 71856
rect 1104 71216 6000 71312
rect 578000 71216 582820 71312
rect 1104 70672 6000 70768
rect 578000 70672 582820 70768
rect 1104 70128 6000 70224
rect 578000 70128 582820 70224
rect 1104 69584 6000 69680
rect 578000 69584 582820 69680
rect 1104 69040 6000 69136
rect 578000 69040 582820 69136
rect 1104 68496 6000 68592
rect 578000 68496 582820 68592
rect 1104 67952 6000 68048
rect 578000 67952 582820 68048
rect 1104 67408 6000 67504
rect 578000 67408 582820 67504
rect 1104 66864 6000 66960
rect 578000 66864 582820 66960
rect 1104 66320 6000 66416
rect 578000 66320 582820 66416
rect 1104 65776 6000 65872
rect 578000 65776 582820 65872
rect 1104 65232 6000 65328
rect 578000 65232 582820 65328
rect 574922 64812 574928 64864
rect 574980 64852 574986 64864
rect 579798 64852 579804 64864
rect 574980 64824 579804 64852
rect 574980 64812 574986 64824
rect 579798 64812 579804 64824
rect 579856 64812 579862 64864
rect 1104 64688 6000 64784
rect 578000 64688 582820 64784
rect 1104 64144 6000 64240
rect 578000 64144 582820 64240
rect 1104 63600 6000 63696
rect 578000 63600 582820 63696
rect 1104 63056 6000 63152
rect 578000 63056 582820 63152
rect 1104 62512 6000 62608
rect 578000 62512 582820 62608
rect 1104 61968 6000 62064
rect 578000 61968 582820 62064
rect 1104 61424 6000 61520
rect 578000 61424 582820 61520
rect 1104 60880 6000 60976
rect 578000 60880 582820 60976
rect 1104 60336 6000 60432
rect 578000 60336 582820 60432
rect 1104 59792 6000 59888
rect 578000 59792 582820 59888
rect 1104 59248 6000 59344
rect 578000 59248 582820 59344
rect 1104 58704 6000 58800
rect 578000 58704 582820 58800
rect 1104 58160 6000 58256
rect 578000 58160 582820 58256
rect 1104 57616 6000 57712
rect 578000 57616 582820 57712
rect 1104 57072 6000 57168
rect 578000 57072 582820 57168
rect 1104 56528 6000 56624
rect 578000 56528 582820 56624
rect 1104 55984 6000 56080
rect 578000 55984 582820 56080
rect 1104 55440 6000 55536
rect 578000 55440 582820 55536
rect 1104 54896 6000 54992
rect 578000 54896 582820 54992
rect 1104 54352 6000 54448
rect 578000 54352 582820 54448
rect 1104 53808 6000 53904
rect 578000 53808 582820 53904
rect 1104 53264 6000 53360
rect 578000 53264 582820 53360
rect 1104 52720 6000 52816
rect 578000 52720 582820 52816
rect 1104 52176 6000 52272
rect 578000 52176 582820 52272
rect 1104 51632 6000 51728
rect 578000 51632 582820 51728
rect 1104 51088 6000 51184
rect 578000 51088 582820 51184
rect 1104 50544 6000 50640
rect 578000 50544 582820 50640
rect 1104 50000 6000 50096
rect 578000 50000 582820 50096
rect 1104 49456 6000 49552
rect 578000 49456 582820 49552
rect 1104 48912 6000 49008
rect 578000 48912 582820 49008
rect 1104 48368 6000 48464
rect 578000 48368 582820 48464
rect 1104 47824 6000 47920
rect 578000 47824 582820 47920
rect 1104 47280 6000 47376
rect 578000 47280 582820 47376
rect 1104 46736 6000 46832
rect 578000 46736 582820 46832
rect 1104 46192 6000 46288
rect 578000 46192 582820 46288
rect 1104 45648 6000 45744
rect 578000 45648 582820 45744
rect 1104 45104 6000 45200
rect 578000 45104 582820 45200
rect 1104 44560 6000 44656
rect 578000 44560 582820 44656
rect 1104 44016 6000 44112
rect 578000 44016 582820 44112
rect 1104 43472 6000 43568
rect 578000 43472 582820 43568
rect 1104 42928 6000 43024
rect 578000 42928 582820 43024
rect 1104 42384 6000 42480
rect 578000 42384 582820 42480
rect 1104 41840 6000 41936
rect 578000 41840 582820 41936
rect 1104 41296 6000 41392
rect 578000 41296 582820 41392
rect 576118 41216 576124 41268
rect 576176 41256 576182 41268
rect 580166 41256 580172 41268
rect 576176 41228 580172 41256
rect 576176 41216 576182 41228
rect 580166 41216 580172 41228
rect 580224 41216 580230 41268
rect 1104 40752 6000 40848
rect 578000 40752 582820 40848
rect 1104 40208 6000 40304
rect 578000 40208 582820 40304
rect 1104 39664 6000 39760
rect 578000 39664 582820 39760
rect 1104 39120 6000 39216
rect 578000 39120 582820 39216
rect 1104 38576 6000 38672
rect 578000 38576 582820 38672
rect 1104 38032 6000 38128
rect 578000 38032 582820 38128
rect 1104 37488 6000 37584
rect 578000 37488 582820 37584
rect 1104 36944 6000 37040
rect 578000 36944 582820 37040
rect 1104 36400 6000 36496
rect 578000 36400 582820 36496
rect 1104 35856 6000 35952
rect 578000 35856 582820 35952
rect 3418 35776 3424 35828
rect 3476 35816 3482 35828
rect 7558 35816 7564 35828
rect 3476 35788 7564 35816
rect 3476 35776 3482 35788
rect 7558 35776 7564 35788
rect 7616 35776 7622 35828
rect 1104 35312 6000 35408
rect 578000 35312 582820 35408
rect 1104 34768 6000 34864
rect 578000 34768 582820 34864
rect 1104 34224 6000 34320
rect 578000 34224 582820 34320
rect 1104 33680 6000 33776
rect 578000 33680 582820 33776
rect 1104 33136 6000 33232
rect 578000 33136 582820 33232
rect 1104 32592 6000 32688
rect 578000 32592 582820 32688
rect 1104 32048 6000 32144
rect 578000 32048 582820 32144
rect 1104 31504 6000 31600
rect 578000 31504 582820 31600
rect 1104 30960 6000 31056
rect 578000 30960 582820 31056
rect 1104 30416 6000 30512
rect 578000 30416 582820 30512
rect 577498 30268 577504 30320
rect 577556 30308 577562 30320
rect 579614 30308 579620 30320
rect 577556 30280 579620 30308
rect 577556 30268 577562 30280
rect 579614 30268 579620 30280
rect 579672 30268 579678 30320
rect 1104 29872 6000 29968
rect 578000 29872 582820 29968
rect 1104 29328 6000 29424
rect 578000 29328 582820 29424
rect 1104 28784 6000 28880
rect 578000 28784 582820 28880
rect 1104 28240 6000 28336
rect 578000 28240 582820 28336
rect 1104 27696 6000 27792
rect 578000 27696 582820 27792
rect 1104 27152 6000 27248
rect 578000 27152 582820 27248
rect 1104 26608 6000 26704
rect 578000 26608 582820 26704
rect 1104 26064 6000 26160
rect 578000 26064 582820 26160
rect 1104 25520 6000 25616
rect 578000 25520 582820 25616
rect 1104 24976 6000 25072
rect 578000 24976 582820 25072
rect 1104 24432 6000 24528
rect 578000 24432 582820 24528
rect 1104 23888 6000 23984
rect 578000 23888 582820 23984
rect 1104 23344 6000 23440
rect 578000 23344 582820 23440
rect 1104 22800 6000 22896
rect 578000 22800 582820 22896
rect 1104 22256 6000 22352
rect 578000 22256 582820 22352
rect 2774 21836 2780 21888
rect 2832 21876 2838 21888
rect 4798 21876 4804 21888
rect 2832 21848 4804 21876
rect 2832 21836 2838 21848
rect 4798 21836 4804 21848
rect 4856 21836 4862 21888
rect 1104 21712 6000 21808
rect 578000 21712 582820 21808
rect 1104 21168 6000 21264
rect 578000 21168 582820 21264
rect 1104 20624 6000 20720
rect 578000 20624 582820 20720
rect 1104 20080 6000 20176
rect 578000 20080 582820 20176
rect 1104 19536 6000 19632
rect 578000 19536 582820 19632
rect 1104 18992 6000 19088
rect 578000 18992 582820 19088
rect 1104 18448 6000 18544
rect 578000 18448 582820 18544
rect 1104 17904 6000 18000
rect 578000 17904 582820 18000
rect 575014 17824 575020 17876
rect 575072 17864 575078 17876
rect 580166 17864 580172 17876
rect 575072 17836 580172 17864
rect 575072 17824 575078 17836
rect 580166 17824 580172 17836
rect 580224 17824 580230 17876
rect 1104 17360 6000 17456
rect 578000 17360 582820 17456
rect 1104 16816 6000 16912
rect 578000 16816 582820 16912
rect 1104 16272 6000 16368
rect 578000 16272 582820 16368
rect 1104 15728 6000 15824
rect 578000 15728 582820 15824
rect 1104 15184 6000 15280
rect 578000 15184 582820 15280
rect 1104 14640 6000 14736
rect 578000 14640 582820 14736
rect 1104 14096 6000 14192
rect 578000 14096 582820 14192
rect 1104 13552 6000 13648
rect 578000 13552 582820 13648
rect 1104 13008 6000 13104
rect 578000 13008 582820 13104
rect 1104 12464 6000 12560
rect 578000 12464 582820 12560
rect 1104 11920 6000 12016
rect 578000 11920 582820 12016
rect 1104 11376 6000 11472
rect 578000 11376 582820 11472
rect 1104 10832 6000 10928
rect 578000 10832 582820 10928
rect 1104 10288 6000 10384
rect 578000 10288 582820 10384
rect 1104 9744 6000 9840
rect 578000 9744 582820 9840
rect 1104 9200 6000 9296
rect 578000 9200 582820 9296
rect 1104 8656 6000 8752
rect 578000 8656 582820 8752
rect 1104 8112 6000 8208
rect 578000 8112 582820 8208
rect 1104 7568 6000 7664
rect 578000 7568 582820 7664
rect 3142 7148 3148 7200
rect 3200 7188 3206 7200
rect 6178 7188 6184 7200
rect 3200 7160 6184 7188
rect 3200 7148 3206 7160
rect 6178 7148 6184 7160
rect 6236 7148 6242 7200
rect 1104 7024 6000 7120
rect 578000 7024 582820 7120
rect 378134 6808 378140 6860
rect 378192 6848 378198 6860
rect 388254 6848 388260 6860
rect 378192 6820 388260 6848
rect 378192 6808 378198 6820
rect 388254 6808 388260 6820
rect 388312 6808 388318 6860
rect 399662 6808 399668 6860
rect 399720 6848 399726 6860
rect 408494 6848 408500 6860
rect 399720 6820 408500 6848
rect 399720 6808 399726 6820
rect 408494 6808 408500 6820
rect 408552 6808 408558 6860
rect 423490 6808 423496 6860
rect 423548 6848 423554 6860
rect 433886 6848 433892 6860
rect 423548 6820 433892 6848
rect 423548 6808 423554 6820
rect 433886 6808 433892 6820
rect 433944 6808 433950 6860
rect 451826 6808 451832 6860
rect 451884 6848 451890 6860
rect 463326 6848 463332 6860
rect 451884 6820 463332 6848
rect 451884 6808 451890 6820
rect 463326 6808 463332 6820
rect 463384 6808 463390 6860
rect 473354 6808 473360 6860
rect 473412 6848 473418 6860
rect 484394 6848 484400 6860
rect 473412 6820 484400 6848
rect 473412 6808 473418 6820
rect 484394 6808 484400 6820
rect 484452 6808 484458 6860
rect 485866 6808 485872 6860
rect 485924 6848 485930 6860
rect 496814 6848 496820 6860
rect 485924 6820 496820 6848
rect 485924 6808 485930 6820
rect 496814 6808 496820 6820
rect 496872 6808 496878 6860
rect 499482 6808 499488 6860
rect 499540 6848 499546 6860
rect 510430 6848 510436 6860
rect 499540 6820 510436 6848
rect 499540 6808 499546 6820
rect 510430 6808 510436 6820
rect 510488 6808 510494 6860
rect 514202 6808 514208 6860
rect 514260 6848 514266 6860
rect 524506 6848 524512 6860
rect 514260 6820 524512 6848
rect 514260 6808 514266 6820
rect 524506 6808 524512 6820
rect 524564 6808 524570 6860
rect 373626 6740 373632 6792
rect 373684 6780 373690 6792
rect 383562 6780 383568 6792
rect 373684 6752 383568 6780
rect 373684 6740 373690 6752
rect 383562 6740 383568 6752
rect 383620 6740 383626 6792
rect 383838 6740 383844 6792
rect 383896 6780 383902 6792
rect 394234 6780 394240 6792
rect 383896 6752 394240 6780
rect 383896 6740 383902 6752
rect 394234 6740 394240 6752
rect 394292 6740 394298 6792
rect 400766 6740 400772 6792
rect 400824 6780 400830 6792
rect 412082 6780 412088 6792
rect 400824 6752 412088 6780
rect 400824 6740 400830 6752
rect 412082 6740 412088 6752
rect 412140 6740 412146 6792
rect 415578 6740 415584 6792
rect 415636 6780 415642 6792
rect 426526 6780 426532 6792
rect 415636 6752 426532 6780
rect 415636 6740 415642 6752
rect 426526 6740 426532 6752
rect 426584 6740 426590 6792
rect 426894 6740 426900 6792
rect 426952 6780 426958 6792
rect 437474 6780 437480 6792
rect 426952 6752 437480 6780
rect 426952 6740 426958 6752
rect 437474 6740 437480 6752
rect 437532 6740 437538 6792
rect 441614 6740 441620 6792
rect 441672 6780 441678 6792
rect 453114 6780 453120 6792
rect 441672 6752 453120 6780
rect 441672 6740 441678 6752
rect 453114 6740 453120 6752
rect 453172 6740 453178 6792
rect 462038 6740 462044 6792
rect 462096 6780 462102 6792
rect 472894 6780 472900 6792
rect 462096 6752 472900 6780
rect 462096 6740 462102 6752
rect 472894 6740 472900 6752
rect 472952 6740 472958 6792
rect 479058 6740 479064 6792
rect 479116 6780 479122 6792
rect 491110 6780 491116 6792
rect 479116 6752 491116 6780
rect 479116 6740 479122 6752
rect 491110 6740 491116 6752
rect 491168 6740 491174 6792
rect 498286 6740 498292 6792
rect 498344 6780 498350 6792
rect 510522 6780 510528 6792
rect 498344 6752 510528 6780
rect 498344 6740 498350 6752
rect 510522 6740 510528 6752
rect 510580 6740 510586 6792
rect 515306 6740 515312 6792
rect 515364 6780 515370 6792
rect 525794 6780 525800 6792
rect 515364 6752 525800 6780
rect 515364 6740 515370 6752
rect 525794 6740 525800 6752
rect 525852 6740 525858 6792
rect 371326 6672 371332 6724
rect 371384 6712 371390 6724
rect 381170 6712 381176 6724
rect 371384 6684 381176 6712
rect 371384 6672 371390 6684
rect 381170 6672 381176 6684
rect 381228 6672 381234 6724
rect 384942 6672 384948 6724
rect 385000 6712 385006 6724
rect 385000 6684 387196 6712
rect 385000 6672 385006 6684
rect 331674 6604 331680 6656
rect 331732 6644 331738 6656
rect 333974 6644 333980 6656
rect 331732 6616 333980 6644
rect 331732 6604 331738 6616
rect 333974 6604 333980 6616
rect 334032 6604 334038 6656
rect 377030 6604 377036 6656
rect 377088 6644 377094 6656
rect 387058 6644 387064 6656
rect 377088 6616 387064 6644
rect 377088 6604 377094 6616
rect 387058 6604 387064 6616
rect 387116 6604 387122 6656
rect 387168 6644 387196 6684
rect 390554 6672 390560 6724
rect 390612 6712 390618 6724
rect 401318 6712 401324 6724
rect 390612 6684 401324 6712
rect 390612 6672 390618 6684
rect 401318 6672 401324 6684
rect 401376 6672 401382 6724
rect 403066 6672 403072 6724
rect 403124 6712 403130 6724
rect 414474 6712 414480 6724
rect 403124 6684 414480 6712
rect 403124 6672 403130 6684
rect 414474 6672 414480 6684
rect 414532 6672 414538 6724
rect 419166 6712 419172 6724
rect 415872 6684 419172 6712
rect 394050 6644 394056 6656
rect 387168 6616 394056 6644
rect 394050 6604 394056 6616
rect 394108 6604 394114 6656
rect 396258 6604 396264 6656
rect 396316 6644 396322 6656
rect 407298 6644 407304 6656
rect 396316 6616 407304 6644
rect 396316 6604 396322 6616
rect 407298 6604 407304 6616
rect 407356 6604 407362 6656
rect 412545 6647 412603 6653
rect 412545 6613 412557 6647
rect 412591 6644 412603 6647
rect 415872 6644 415900 6684
rect 419166 6672 419172 6684
rect 419224 6672 419230 6724
rect 434806 6672 434812 6724
rect 434864 6712 434870 6724
rect 445846 6712 445852 6724
rect 434864 6684 445852 6712
rect 434864 6672 434870 6684
rect 445846 6672 445852 6684
rect 445904 6672 445910 6724
rect 449526 6672 449532 6724
rect 449584 6712 449590 6724
rect 459554 6712 459560 6724
rect 449584 6684 459560 6712
rect 449584 6672 449590 6684
rect 459554 6672 459560 6684
rect 459612 6672 459618 6724
rect 460934 6672 460940 6724
rect 460992 6712 460998 6724
rect 472526 6712 472532 6724
rect 460992 6684 472532 6712
rect 460992 6672 460998 6684
rect 472526 6672 472532 6684
rect 472584 6672 472590 6724
rect 476758 6672 476764 6724
rect 476816 6712 476822 6724
rect 487430 6712 487436 6724
rect 476816 6684 487436 6712
rect 476816 6672 476822 6684
rect 487430 6672 487436 6684
rect 487488 6672 487494 6724
rect 493778 6672 493784 6724
rect 493836 6712 493842 6724
rect 503898 6712 503904 6724
rect 493836 6684 503904 6712
rect 493836 6672 493842 6684
rect 503898 6672 503904 6684
rect 503956 6672 503962 6724
rect 505094 6672 505100 6724
rect 505152 6712 505158 6724
rect 521470 6712 521476 6724
rect 505152 6684 521476 6712
rect 505152 6672 505158 6684
rect 521470 6672 521476 6684
rect 521528 6672 521534 6724
rect 523218 6672 523224 6724
rect 523276 6712 523282 6724
rect 540514 6712 540520 6724
rect 523276 6684 540520 6712
rect 523276 6672 523282 6684
rect 540514 6672 540520 6684
rect 540572 6672 540578 6724
rect 412591 6616 415900 6644
rect 412591 6613 412603 6616
rect 412545 6607 412603 6613
rect 418982 6604 418988 6656
rect 419040 6644 419046 6656
rect 429194 6644 429200 6656
rect 419040 6616 429200 6644
rect 419040 6604 419046 6616
rect 429194 6604 429200 6616
rect 429252 6604 429258 6656
rect 431402 6604 431408 6656
rect 431460 6644 431466 6656
rect 442350 6644 442356 6656
rect 431460 6616 442356 6644
rect 431460 6604 431466 6616
rect 442350 6604 442356 6616
rect 442408 6604 442414 6656
rect 446122 6604 446128 6656
rect 446180 6644 446186 6656
rect 456794 6644 456800 6656
rect 446180 6616 456800 6644
rect 446180 6604 446186 6616
rect 456794 6604 456800 6616
rect 456852 6604 456858 6656
rect 464246 6604 464252 6656
rect 464304 6644 464310 6656
rect 474734 6644 474740 6656
rect 464304 6616 474740 6644
rect 464304 6604 464310 6616
rect 474734 6604 474740 6616
rect 474792 6604 474798 6656
rect 477862 6604 477868 6656
rect 477920 6644 477926 6656
rect 488534 6644 488540 6656
rect 477920 6616 488540 6644
rect 477920 6604 477926 6616
rect 488534 6604 488540 6616
rect 488592 6604 488598 6656
rect 506198 6604 506204 6656
rect 506256 6644 506262 6656
rect 520826 6644 520832 6656
rect 506256 6616 520832 6644
rect 506256 6604 506262 6616
rect 520826 6604 520832 6616
rect 520884 6604 520890 6656
rect 524414 6604 524420 6656
rect 524472 6644 524478 6656
rect 536742 6644 536748 6656
rect 524472 6616 536748 6644
rect 524472 6604 524478 6616
rect 536742 6604 536748 6616
rect 536800 6604 536806 6656
rect 1104 6480 6000 6576
rect 360010 6536 360016 6588
rect 360068 6576 360074 6588
rect 369210 6576 369216 6588
rect 360068 6548 369216 6576
rect 360068 6536 360074 6548
rect 369210 6536 369216 6548
rect 369268 6536 369274 6588
rect 370222 6536 370228 6588
rect 370280 6576 370286 6588
rect 379974 6576 379980 6588
rect 370280 6548 379980 6576
rect 370280 6536 370286 6548
rect 379974 6536 379980 6548
rect 380032 6536 380038 6588
rect 401962 6536 401968 6588
rect 402020 6576 402026 6588
rect 413278 6576 413284 6588
rect 402020 6548 413284 6576
rect 402020 6536 402026 6548
rect 413278 6536 413284 6548
rect 413336 6536 413342 6588
rect 416682 6536 416688 6588
rect 416740 6576 416746 6588
rect 426434 6576 426440 6588
rect 416740 6548 426440 6576
rect 416740 6536 416746 6548
rect 426434 6536 426440 6548
rect 426492 6536 426498 6588
rect 426526 6536 426532 6588
rect 426584 6576 426590 6588
rect 427538 6576 427544 6588
rect 426584 6548 427544 6576
rect 426584 6536 426590 6548
rect 427538 6536 427544 6548
rect 427596 6536 427602 6588
rect 430298 6536 430304 6588
rect 430356 6576 430362 6588
rect 439038 6576 439044 6588
rect 430356 6548 439044 6576
rect 430356 6536 430362 6548
rect 439038 6536 439044 6548
rect 439096 6536 439102 6588
rect 442718 6536 442724 6588
rect 442776 6576 442782 6588
rect 453666 6576 453672 6588
rect 442776 6548 453672 6576
rect 442776 6536 442782 6548
rect 453666 6536 453672 6548
rect 453724 6536 453730 6588
rect 454126 6536 454132 6588
rect 454184 6576 454190 6588
rect 464430 6576 464436 6588
rect 454184 6548 464436 6576
rect 454184 6536 454190 6548
rect 464430 6536 464436 6548
rect 464488 6536 464494 6588
rect 467650 6536 467656 6588
rect 467708 6576 467714 6588
rect 477586 6576 477592 6588
rect 467708 6548 477592 6576
rect 467708 6536 467714 6548
rect 477586 6536 477592 6548
rect 477644 6536 477650 6588
rect 482462 6536 482468 6588
rect 482520 6576 482526 6588
rect 497734 6576 497740 6588
rect 482520 6548 497740 6576
rect 482520 6536 482526 6548
rect 497734 6536 497740 6548
rect 497792 6536 497798 6588
rect 502794 6536 502800 6588
rect 502852 6576 502858 6588
rect 519078 6576 519084 6588
rect 502852 6548 519084 6576
rect 502852 6536 502858 6548
rect 519078 6536 519084 6548
rect 519136 6536 519142 6588
rect 521010 6536 521016 6588
rect 521068 6576 521074 6588
rect 535914 6576 535920 6588
rect 521068 6548 535920 6576
rect 521068 6536 521074 6548
rect 535914 6536 535920 6548
rect 535972 6536 535978 6588
rect 70670 6468 70676 6520
rect 70728 6508 70734 6520
rect 75454 6508 75460 6520
rect 70728 6480 75460 6508
rect 70728 6468 70734 6480
rect 75454 6468 75460 6480
rect 75512 6468 75518 6520
rect 356606 6468 356612 6520
rect 356664 6508 356670 6520
rect 365714 6508 365720 6520
rect 356664 6480 365720 6508
rect 356664 6468 356670 6480
rect 365714 6468 365720 6480
rect 365772 6468 365778 6520
rect 369026 6468 369032 6520
rect 369084 6508 369090 6520
rect 378686 6508 378692 6520
rect 369084 6480 378692 6508
rect 369084 6468 369090 6480
rect 378686 6468 378692 6480
rect 378744 6468 378750 6520
rect 382642 6468 382648 6520
rect 382700 6508 382706 6520
rect 392762 6508 392768 6520
rect 382700 6480 392768 6508
rect 382700 6468 382706 6480
rect 392762 6468 392768 6480
rect 392820 6468 392826 6520
rect 392854 6468 392860 6520
rect 392912 6508 392918 6520
rect 403710 6508 403716 6520
rect 392912 6480 403716 6508
rect 392912 6468 392918 6480
rect 403710 6468 403716 6480
rect 403768 6468 403774 6520
rect 407574 6468 407580 6520
rect 407632 6508 407638 6520
rect 407632 6480 409828 6508
rect 407632 6468 407638 6480
rect 362218 6400 362224 6452
rect 362276 6440 362282 6452
rect 371602 6440 371608 6452
rect 362276 6412 371608 6440
rect 362276 6400 362282 6412
rect 371602 6400 371608 6412
rect 371660 6400 371666 6452
rect 374730 6400 374736 6452
rect 374788 6440 374794 6452
rect 384666 6440 384672 6452
rect 374788 6412 384672 6440
rect 374788 6400 374794 6412
rect 384666 6400 384672 6412
rect 384724 6400 384730 6452
rect 387242 6400 387248 6452
rect 387300 6440 387306 6452
rect 397822 6440 397828 6452
rect 387300 6412 397828 6440
rect 387300 6400 387306 6412
rect 397822 6400 397828 6412
rect 397880 6400 397886 6452
rect 398558 6400 398564 6452
rect 398616 6440 398622 6452
rect 409690 6440 409696 6452
rect 398616 6412 409696 6440
rect 398616 6400 398622 6412
rect 409690 6400 409696 6412
rect 409748 6400 409754 6452
rect 409800 6440 409828 6480
rect 412174 6468 412180 6520
rect 412232 6508 412238 6520
rect 423582 6508 423588 6520
rect 412232 6480 423588 6508
rect 412232 6468 412238 6480
rect 423582 6468 423588 6480
rect 423640 6468 423646 6520
rect 424594 6468 424600 6520
rect 424652 6508 424658 6520
rect 434530 6508 434536 6520
rect 424652 6480 434536 6508
rect 424652 6468 424658 6480
rect 434530 6468 434536 6480
rect 434588 6468 434594 6520
rect 437106 6468 437112 6520
rect 437164 6508 437170 6520
rect 447134 6508 447140 6520
rect 437164 6480 447140 6508
rect 437164 6468 437170 6480
rect 447134 6468 447140 6480
rect 447192 6468 447198 6520
rect 457530 6468 457536 6520
rect 457588 6508 457594 6520
rect 467834 6508 467840 6520
rect 457588 6480 467840 6508
rect 457588 6468 457594 6480
rect 467834 6468 467840 6480
rect 467892 6468 467898 6520
rect 472250 6468 472256 6520
rect 472308 6508 472314 6520
rect 483290 6508 483296 6520
rect 472308 6480 483296 6508
rect 472308 6468 472314 6480
rect 483290 6468 483296 6480
rect 483348 6468 483354 6520
rect 484670 6468 484676 6520
rect 484728 6508 484734 6520
rect 500126 6508 500132 6520
rect 484728 6480 500132 6508
rect 484728 6468 484734 6480
rect 500126 6468 500132 6480
rect 500184 6468 500190 6520
rect 503990 6468 503996 6520
rect 504048 6508 504054 6520
rect 514754 6508 514760 6520
rect 504048 6480 514760 6508
rect 504048 6468 504054 6480
rect 514754 6468 514760 6480
rect 514812 6468 514818 6520
rect 517606 6468 517612 6520
rect 517664 6508 517670 6520
rect 534534 6508 534540 6520
rect 517664 6480 534540 6508
rect 517664 6468 517670 6480
rect 534534 6468 534540 6480
rect 534592 6468 534598 6520
rect 578000 6480 582820 6576
rect 412545 6443 412603 6449
rect 412545 6440 412557 6443
rect 409800 6412 412557 6440
rect 412545 6409 412557 6412
rect 412591 6409 412603 6443
rect 412545 6403 412603 6409
rect 417786 6400 417792 6452
rect 417844 6440 417850 6452
rect 427814 6440 427820 6452
rect 417844 6412 427820 6440
rect 417844 6400 417850 6412
rect 427814 6400 427820 6412
rect 427872 6400 427878 6452
rect 435910 6400 435916 6452
rect 435968 6440 435974 6452
rect 445754 6440 445760 6452
rect 435968 6412 445760 6440
rect 435968 6400 435974 6412
rect 445754 6400 445760 6412
rect 445812 6400 445818 6452
rect 448422 6400 448428 6452
rect 448480 6440 448486 6452
rect 458174 6440 458180 6452
rect 448480 6412 458180 6440
rect 448480 6400 448486 6412
rect 458174 6400 458180 6412
rect 458232 6400 458238 6452
rect 466546 6400 466552 6452
rect 466604 6440 466610 6452
rect 477494 6440 477500 6452
rect 466604 6412 477500 6440
rect 466604 6400 466610 6412
rect 477494 6400 477500 6412
rect 477552 6400 477558 6452
rect 481266 6400 481272 6452
rect 481324 6440 481330 6452
rect 496538 6440 496544 6452
rect 481324 6412 496544 6440
rect 481324 6400 481330 6412
rect 496538 6400 496544 6412
rect 496596 6400 496602 6452
rect 497182 6400 497188 6452
rect 497240 6440 497246 6452
rect 513190 6440 513196 6452
rect 497240 6412 513196 6440
rect 497240 6400 497246 6412
rect 513190 6400 513196 6412
rect 513248 6400 513254 6452
rect 93302 6332 93308 6384
rect 93360 6372 93366 6384
rect 96982 6372 96988 6384
rect 93360 6344 96988 6372
rect 93360 6332 93366 6344
rect 96982 6332 96988 6344
rect 97040 6332 97046 6384
rect 272702 6332 272708 6384
rect 272760 6372 272766 6384
rect 275094 6372 275100 6384
rect 272760 6344 275100 6372
rect 272760 6332 272766 6344
rect 275094 6332 275100 6344
rect 275152 6332 275158 6384
rect 284018 6332 284024 6384
rect 284076 6372 284082 6384
rect 285674 6372 285680 6384
rect 284076 6344 285680 6372
rect 284076 6332 284082 6344
rect 285674 6332 285680 6344
rect 285732 6332 285738 6384
rect 319162 6332 319168 6384
rect 319220 6372 319226 6384
rect 322474 6372 322480 6384
rect 319220 6344 322480 6372
rect 319220 6332 319226 6344
rect 322474 6332 322480 6344
rect 322532 6332 322538 6384
rect 328270 6332 328276 6384
rect 328328 6372 328334 6384
rect 330570 6372 330576 6384
rect 328328 6344 330576 6372
rect 328328 6332 328334 6344
rect 330570 6332 330576 6344
rect 330628 6332 330634 6384
rect 340690 6332 340696 6384
rect 340748 6372 340754 6384
rect 342714 6372 342720 6384
rect 340748 6344 342720 6372
rect 340748 6332 340754 6344
rect 342714 6332 342720 6344
rect 342772 6332 342778 6384
rect 347498 6332 347504 6384
rect 347556 6372 347562 6384
rect 356146 6372 356152 6384
rect 347556 6344 356152 6372
rect 347556 6332 347562 6344
rect 356146 6332 356152 6344
rect 356204 6332 356210 6384
rect 361114 6332 361120 6384
rect 361172 6372 361178 6384
rect 370406 6372 370412 6384
rect 361172 6344 370412 6372
rect 361172 6332 361178 6344
rect 370406 6332 370412 6344
rect 370464 6332 370470 6384
rect 379238 6332 379244 6384
rect 379296 6372 379302 6384
rect 389082 6372 389088 6384
rect 379296 6344 389088 6372
rect 379296 6332 379302 6344
rect 389082 6332 389088 6344
rect 389140 6332 389146 6384
rect 391750 6332 391756 6384
rect 391808 6372 391814 6384
rect 402514 6372 402520 6384
rect 391808 6344 402520 6372
rect 391808 6332 391814 6344
rect 402514 6332 402520 6344
rect 402572 6332 402578 6384
rect 406470 6332 406476 6384
rect 406528 6372 406534 6384
rect 417970 6372 417976 6384
rect 406528 6344 417976 6372
rect 406528 6332 406534 6344
rect 417970 6332 417976 6344
rect 418028 6332 418034 6384
rect 421190 6332 421196 6384
rect 421248 6372 421254 6384
rect 432690 6372 432696 6384
rect 421248 6344 432696 6372
rect 421248 6332 421254 6344
rect 432690 6332 432696 6344
rect 432748 6332 432754 6384
rect 438210 6332 438216 6384
rect 438268 6372 438274 6384
rect 448606 6372 448612 6384
rect 438268 6344 448612 6372
rect 438268 6332 438274 6344
rect 448606 6332 448612 6344
rect 448664 6332 448670 6384
rect 450722 6332 450728 6384
rect 450780 6372 450786 6384
rect 462222 6372 462228 6384
rect 450780 6344 462228 6372
rect 450780 6332 450786 6344
rect 462222 6332 462228 6344
rect 462280 6332 462286 6384
rect 468846 6332 468852 6384
rect 468904 6372 468910 6384
rect 478966 6372 478972 6384
rect 468904 6344 478972 6372
rect 468904 6332 468910 6344
rect 478966 6332 478972 6344
rect 479024 6332 479030 6384
rect 483566 6332 483572 6384
rect 483624 6372 483630 6384
rect 489457 6375 489515 6381
rect 489457 6372 489469 6375
rect 483624 6344 489469 6372
rect 483624 6332 483630 6344
rect 489457 6341 489469 6344
rect 489503 6341 489515 6375
rect 489457 6335 489515 6341
rect 491478 6332 491484 6384
rect 491536 6372 491542 6384
rect 507210 6372 507216 6384
rect 491536 6344 507216 6372
rect 491536 6332 491542 6344
rect 507210 6332 507216 6344
rect 507268 6332 507274 6384
rect 507394 6332 507400 6384
rect 507452 6372 507458 6384
rect 523862 6372 523868 6384
rect 507452 6344 523868 6372
rect 507452 6332 507458 6344
rect 523862 6332 523868 6344
rect 523920 6332 523926 6384
rect 353202 6264 353208 6316
rect 353260 6304 353266 6316
rect 362126 6304 362132 6316
rect 353260 6276 362132 6304
rect 353260 6264 353266 6276
rect 362126 6264 362132 6276
rect 362184 6264 362190 6316
rect 364518 6264 364524 6316
rect 364576 6304 364582 6316
rect 367462 6304 367468 6316
rect 364576 6276 367468 6304
rect 364576 6264 364582 6276
rect 367462 6264 367468 6276
rect 367520 6264 367526 6316
rect 367922 6264 367928 6316
rect 367980 6304 367986 6316
rect 377582 6304 377588 6316
rect 367980 6276 377588 6304
rect 367980 6264 367986 6276
rect 377582 6264 377588 6276
rect 377640 6264 377646 6316
rect 386046 6264 386052 6316
rect 386104 6304 386110 6316
rect 396626 6304 396632 6316
rect 386104 6276 396632 6304
rect 386104 6264 386110 6276
rect 396626 6264 396632 6276
rect 396684 6264 396690 6316
rect 397362 6264 397368 6316
rect 397420 6304 397426 6316
rect 408402 6304 408408 6316
rect 397420 6276 408408 6304
rect 397420 6264 397426 6276
rect 408402 6264 408408 6276
rect 408460 6264 408466 6316
rect 413186 6264 413192 6316
rect 413244 6304 413250 6316
rect 424962 6304 424968 6316
rect 413244 6276 424968 6304
rect 413244 6264 413250 6276
rect 424962 6264 424968 6276
rect 425020 6264 425026 6316
rect 429102 6264 429108 6316
rect 429160 6304 429166 6316
rect 438854 6304 438860 6316
rect 429160 6276 438860 6304
rect 429160 6264 429166 6276
rect 438854 6264 438860 6276
rect 438912 6264 438918 6316
rect 443914 6264 443920 6316
rect 443972 6304 443978 6316
rect 454126 6304 454132 6316
rect 443972 6276 454132 6304
rect 443972 6264 443978 6276
rect 454126 6264 454132 6276
rect 454184 6264 454190 6316
rect 458634 6264 458640 6316
rect 458692 6304 458698 6316
rect 469490 6304 469496 6316
rect 458692 6276 469496 6304
rect 458692 6264 458698 6276
rect 469490 6264 469496 6276
rect 469548 6264 469554 6316
rect 480162 6264 480168 6316
rect 480220 6304 480226 6316
rect 490742 6304 490748 6316
rect 480220 6276 490748 6304
rect 480220 6264 480226 6276
rect 490742 6264 490748 6276
rect 490800 6264 490806 6316
rect 494882 6264 494888 6316
rect 494940 6304 494946 6316
rect 510798 6304 510804 6316
rect 494940 6276 510804 6304
rect 494940 6264 494946 6276
rect 510798 6264 510804 6276
rect 510856 6264 510862 6316
rect 516410 6264 516416 6316
rect 516468 6304 516474 6316
rect 533338 6304 533344 6316
rect 516468 6276 533344 6304
rect 516468 6264 516474 6276
rect 533338 6264 533344 6276
rect 533396 6264 533402 6316
rect 83826 6196 83832 6248
rect 83884 6236 83890 6248
rect 87874 6236 87880 6248
rect 83884 6208 87880 6236
rect 83884 6196 83890 6208
rect 87874 6196 87880 6208
rect 87932 6196 87938 6248
rect 264790 6196 264796 6248
rect 264848 6236 264854 6248
rect 266354 6236 266360 6248
rect 264848 6208 266360 6236
rect 264848 6196 264854 6208
rect 266354 6196 266360 6208
rect 266412 6196 266418 6248
rect 273806 6196 273812 6248
rect 273864 6236 273870 6248
rect 276014 6236 276020 6248
rect 273864 6208 276020 6236
rect 273864 6196 273870 6208
rect 276014 6196 276020 6208
rect 276072 6196 276078 6248
rect 337286 6196 337292 6248
rect 337344 6236 337350 6248
rect 339678 6236 339684 6248
rect 337344 6208 339684 6236
rect 337344 6196 337350 6208
rect 339678 6196 339684 6208
rect 339736 6196 339742 6248
rect 354306 6196 354312 6248
rect 354364 6236 354370 6248
rect 363322 6236 363328 6248
rect 354364 6208 363328 6236
rect 354364 6196 354370 6208
rect 363322 6196 363328 6208
rect 363380 6196 363386 6248
rect 363414 6196 363420 6248
rect 363472 6236 363478 6248
rect 372798 6236 372804 6248
rect 363472 6208 372804 6236
rect 363472 6196 363478 6208
rect 372798 6196 372804 6208
rect 372856 6196 372862 6248
rect 375834 6196 375840 6248
rect 375892 6236 375898 6248
rect 385862 6236 385868 6248
rect 375892 6208 385868 6236
rect 375892 6196 375898 6208
rect 385862 6196 385868 6208
rect 385920 6196 385926 6248
rect 388346 6196 388352 6248
rect 388404 6236 388410 6248
rect 399018 6236 399024 6248
rect 388404 6208 399024 6236
rect 388404 6196 388410 6208
rect 399018 6196 399024 6208
rect 399076 6196 399082 6248
rect 404170 6196 404176 6248
rect 404228 6236 404234 6248
rect 414106 6236 414112 6248
rect 404228 6208 414112 6236
rect 404228 6196 404234 6208
rect 414106 6196 414112 6208
rect 414164 6196 414170 6248
rect 420086 6196 420092 6248
rect 420144 6236 420150 6248
rect 430574 6236 430580 6248
rect 420144 6208 430580 6236
rect 420144 6196 420150 6208
rect 430574 6196 430580 6208
rect 430632 6196 430638 6248
rect 432506 6196 432512 6248
rect 432564 6236 432570 6248
rect 443546 6236 443552 6248
rect 432564 6208 443552 6236
rect 432564 6196 432570 6208
rect 443546 6196 443552 6208
rect 443604 6196 443610 6248
rect 447318 6196 447324 6248
rect 447376 6236 447382 6248
rect 458266 6236 458272 6248
rect 447376 6208 458272 6236
rect 447376 6196 447382 6208
rect 458266 6196 458272 6208
rect 458324 6196 458330 6248
rect 463142 6196 463148 6248
rect 463200 6236 463206 6248
rect 474090 6236 474096 6248
rect 463200 6208 474096 6236
rect 463200 6196 463206 6208
rect 474090 6196 474096 6208
rect 474148 6196 474154 6248
rect 475654 6196 475660 6248
rect 475712 6236 475718 6248
rect 484670 6236 484676 6248
rect 475712 6208 484676 6236
rect 475712 6196 475718 6208
rect 484670 6196 484676 6208
rect 484728 6196 484734 6248
rect 486970 6196 486976 6248
rect 487028 6236 487034 6248
rect 502426 6236 502432 6248
rect 487028 6208 502432 6236
rect 487028 6196 487034 6208
rect 502426 6196 502432 6208
rect 502484 6196 502490 6248
rect 508498 6196 508504 6248
rect 508556 6236 508562 6248
rect 525058 6236 525064 6248
rect 508556 6208 525064 6236
rect 508556 6196 508562 6208
rect 525058 6196 525064 6208
rect 525116 6196 525122 6248
rect 530026 6196 530032 6248
rect 530084 6236 530090 6248
rect 541434 6236 541440 6248
rect 530084 6208 541440 6236
rect 530084 6196 530090 6208
rect 541434 6196 541440 6208
rect 541492 6196 541498 6248
rect 5534 6128 5540 6180
rect 5592 6168 5598 6180
rect 10778 6168 10784 6180
rect 5592 6140 10784 6168
rect 5592 6128 5598 6140
rect 10778 6128 10784 6140
rect 10836 6128 10842 6180
rect 63586 6128 63592 6180
rect 63644 6168 63650 6180
rect 68646 6168 68652 6180
rect 63644 6140 68652 6168
rect 63644 6128 63650 6140
rect 68646 6128 68652 6140
rect 68704 6128 68710 6180
rect 87322 6128 87328 6180
rect 87380 6168 87386 6180
rect 91278 6168 91284 6180
rect 87380 6140 91284 6168
rect 87380 6128 87386 6140
rect 91278 6128 91284 6140
rect 91336 6128 91342 6180
rect 199010 6128 199016 6180
rect 199068 6168 199074 6180
rect 200390 6168 200396 6180
rect 199068 6140 200396 6168
rect 199068 6128 199074 6140
rect 200390 6128 200396 6140
rect 200448 6128 200454 6180
rect 235258 6128 235264 6180
rect 235316 6168 235322 6180
rect 238386 6168 238392 6180
rect 235316 6140 238392 6168
rect 235316 6128 235322 6140
rect 238386 6128 238392 6140
rect 238444 6128 238450 6180
rect 342990 6128 342996 6180
rect 343048 6168 343054 6180
rect 345934 6168 345940 6180
rect 343048 6140 345940 6168
rect 343048 6128 343054 6140
rect 345934 6128 345940 6140
rect 345992 6128 345998 6180
rect 355410 6128 355416 6180
rect 355468 6168 355474 6180
rect 364518 6168 364524 6180
rect 355468 6140 364524 6168
rect 355468 6128 355474 6140
rect 364518 6128 364524 6140
rect 364576 6128 364582 6180
rect 372430 6128 372436 6180
rect 372488 6168 372494 6180
rect 382366 6168 382372 6180
rect 372488 6140 382372 6168
rect 372488 6128 372494 6140
rect 382366 6128 382372 6140
rect 382424 6128 382430 6180
rect 389450 6128 389456 6180
rect 389508 6168 389514 6180
rect 400214 6168 400220 6180
rect 389508 6140 400220 6168
rect 389508 6128 389514 6140
rect 400214 6128 400220 6140
rect 400272 6128 400278 6180
rect 405366 6128 405372 6180
rect 405424 6168 405430 6180
rect 416682 6168 416688 6180
rect 405424 6140 416688 6168
rect 405424 6128 405430 6140
rect 416682 6128 416688 6140
rect 416740 6128 416746 6180
rect 422386 6128 422392 6180
rect 422444 6168 422450 6180
rect 422444 6140 424456 6168
rect 422444 6128 422450 6140
rect 245470 6060 245476 6112
rect 245528 6100 245534 6112
rect 247034 6100 247040 6112
rect 245528 6072 247040 6100
rect 245528 6060 245534 6072
rect 247034 6060 247040 6072
rect 247092 6060 247098 6112
rect 254578 6060 254584 6112
rect 254636 6100 254642 6112
rect 256694 6100 256700 6112
rect 254636 6072 256700 6100
rect 254636 6060 254642 6072
rect 256694 6060 256700 6072
rect 256752 6060 256758 6112
rect 290826 6060 290832 6112
rect 290884 6100 290890 6112
rect 292574 6100 292580 6112
rect 290884 6072 292580 6100
rect 290884 6060 290890 6072
rect 292574 6060 292580 6072
rect 292632 6060 292638 6112
rect 293126 6060 293132 6112
rect 293184 6100 293190 6112
rect 295426 6100 295432 6112
rect 293184 6072 295432 6100
rect 293184 6060 293190 6072
rect 295426 6060 295432 6072
rect 295484 6060 295490 6112
rect 302142 6060 302148 6112
rect 302200 6100 302206 6112
rect 304258 6100 304264 6112
rect 302200 6072 304264 6100
rect 302200 6060 302206 6072
rect 304258 6060 304264 6072
rect 304316 6060 304322 6112
rect 314654 6060 314660 6112
rect 314712 6100 314718 6112
rect 318242 6100 318248 6112
rect 314712 6072 318248 6100
rect 314712 6060 314718 6072
rect 318242 6060 318248 6072
rect 318300 6060 318306 6112
rect 332778 6060 332784 6112
rect 332836 6100 332842 6112
rect 336274 6100 336280 6112
rect 332836 6072 336280 6100
rect 332836 6060 332842 6072
rect 336274 6060 336280 6072
rect 336332 6060 336338 6112
rect 393958 6060 393964 6112
rect 394016 6100 394022 6112
rect 403802 6100 403808 6112
rect 394016 6072 403808 6100
rect 394016 6060 394022 6072
rect 403802 6060 403808 6072
rect 403860 6060 403866 6112
rect 414382 6060 414388 6112
rect 414440 6100 414446 6112
rect 424318 6100 424324 6112
rect 414440 6072 424324 6100
rect 414440 6060 414446 6072
rect 424318 6060 424324 6072
rect 424376 6060 424382 6112
rect 424428 6100 424456 6140
rect 427998 6128 428004 6180
rect 428056 6168 428062 6180
rect 438946 6168 438952 6180
rect 428056 6140 438952 6168
rect 428056 6128 428062 6140
rect 438946 6128 438952 6140
rect 439004 6128 439010 6180
rect 452930 6128 452936 6180
rect 452988 6168 452994 6180
rect 463694 6168 463700 6180
rect 452988 6140 463700 6168
rect 452988 6128 452994 6140
rect 463694 6128 463700 6140
rect 463752 6128 463758 6180
rect 474458 6128 474464 6180
rect 474516 6168 474522 6180
rect 489178 6168 489184 6180
rect 474516 6140 489184 6168
rect 474516 6128 474522 6140
rect 489178 6128 489184 6140
rect 489236 6128 489242 6180
rect 489270 6128 489276 6180
rect 489328 6168 489334 6180
rect 500586 6168 500592 6180
rect 489328 6140 500592 6168
rect 489328 6128 489334 6140
rect 500586 6128 500592 6140
rect 500644 6128 500650 6180
rect 501690 6128 501696 6180
rect 501748 6168 501754 6180
rect 517882 6168 517888 6180
rect 501748 6140 517888 6168
rect 501748 6128 501754 6140
rect 517882 6128 517888 6140
rect 517940 6128 517946 6180
rect 522114 6128 522120 6180
rect 522172 6168 522178 6180
rect 539318 6168 539324 6180
rect 522172 6140 539324 6168
rect 522172 6128 522178 6140
rect 539318 6128 539324 6140
rect 539376 6128 539382 6180
rect 434622 6100 434628 6112
rect 424428 6072 434628 6100
rect 434622 6060 434628 6072
rect 434680 6060 434686 6112
rect 439314 6060 439320 6112
rect 439372 6100 439378 6112
rect 448514 6100 448520 6112
rect 439372 6072 448520 6100
rect 439372 6060 439378 6072
rect 448514 6060 448520 6072
rect 448572 6060 448578 6112
rect 455230 6060 455236 6112
rect 455288 6100 455294 6112
rect 464246 6100 464252 6112
rect 455288 6072 464252 6100
rect 455288 6060 455294 6072
rect 464246 6060 464252 6072
rect 464304 6060 464310 6112
rect 465442 6060 465448 6112
rect 465500 6100 465506 6112
rect 476114 6100 476120 6112
rect 465500 6072 476120 6100
rect 465500 6060 465506 6072
rect 476114 6060 476120 6072
rect 476172 6060 476178 6112
rect 489457 6103 489515 6109
rect 489457 6069 489469 6103
rect 489503 6100 489515 6103
rect 494146 6100 494152 6112
rect 489503 6072 494152 6100
rect 489503 6069 489515 6072
rect 489457 6063 489515 6069
rect 494146 6060 494152 6072
rect 494204 6060 494210 6112
rect 496078 6060 496084 6112
rect 496136 6100 496142 6112
rect 506474 6100 506480 6112
rect 496136 6072 506480 6100
rect 496136 6060 496142 6072
rect 506474 6060 506480 6072
rect 506532 6060 506538 6112
rect 509602 6060 509608 6112
rect 509660 6100 509666 6112
rect 521194 6100 521200 6112
rect 509660 6072 521200 6100
rect 509660 6060 509666 6072
rect 521194 6060 521200 6072
rect 521252 6060 521258 6112
rect 549346 6060 549352 6112
rect 549404 6100 549410 6112
rect 550542 6100 550548 6112
rect 549404 6072 550548 6100
rect 549404 6060 549410 6072
rect 550542 6060 550548 6072
rect 550600 6060 550606 6112
rect 1104 6010 582820 6032
rect 1104 5958 18822 6010
rect 18874 5958 18886 6010
rect 18938 5958 18950 6010
rect 19002 5958 19014 6010
rect 19066 5958 19078 6010
rect 19130 5958 19142 6010
rect 19194 5958 19206 6010
rect 19258 5958 19270 6010
rect 19322 5958 19334 6010
rect 19386 5958 54822 6010
rect 54874 5958 54886 6010
rect 54938 5958 54950 6010
rect 55002 5958 55014 6010
rect 55066 5958 55078 6010
rect 55130 5958 55142 6010
rect 55194 5958 55206 6010
rect 55258 5958 55270 6010
rect 55322 5958 55334 6010
rect 55386 5958 90822 6010
rect 90874 5958 90886 6010
rect 90938 5958 90950 6010
rect 91002 5958 91014 6010
rect 91066 5958 91078 6010
rect 91130 5958 91142 6010
rect 91194 5958 91206 6010
rect 91258 5958 91270 6010
rect 91322 5958 91334 6010
rect 91386 5958 126822 6010
rect 126874 5958 126886 6010
rect 126938 5958 126950 6010
rect 127002 5958 127014 6010
rect 127066 5958 127078 6010
rect 127130 5958 127142 6010
rect 127194 5958 127206 6010
rect 127258 5958 127270 6010
rect 127322 5958 127334 6010
rect 127386 5958 162822 6010
rect 162874 5958 162886 6010
rect 162938 5958 162950 6010
rect 163002 5958 163014 6010
rect 163066 5958 163078 6010
rect 163130 5958 163142 6010
rect 163194 5958 163206 6010
rect 163258 5958 163270 6010
rect 163322 5958 163334 6010
rect 163386 5958 198822 6010
rect 198874 5958 198886 6010
rect 198938 5958 198950 6010
rect 199002 5958 199014 6010
rect 199066 5958 199078 6010
rect 199130 5958 199142 6010
rect 199194 5958 199206 6010
rect 199258 5958 199270 6010
rect 199322 5958 199334 6010
rect 199386 5958 234822 6010
rect 234874 5958 234886 6010
rect 234938 5958 234950 6010
rect 235002 5958 235014 6010
rect 235066 5958 235078 6010
rect 235130 5958 235142 6010
rect 235194 5958 235206 6010
rect 235258 5958 235270 6010
rect 235322 5958 235334 6010
rect 235386 5958 270822 6010
rect 270874 5958 270886 6010
rect 270938 5958 270950 6010
rect 271002 5958 271014 6010
rect 271066 5958 271078 6010
rect 271130 5958 271142 6010
rect 271194 5958 271206 6010
rect 271258 5958 271270 6010
rect 271322 5958 271334 6010
rect 271386 5958 306822 6010
rect 306874 5958 306886 6010
rect 306938 5958 306950 6010
rect 307002 5958 307014 6010
rect 307066 5958 307078 6010
rect 307130 5958 307142 6010
rect 307194 5958 307206 6010
rect 307258 5958 307270 6010
rect 307322 5958 307334 6010
rect 307386 5958 342822 6010
rect 342874 5958 342886 6010
rect 342938 5958 342950 6010
rect 343002 5958 343014 6010
rect 343066 5958 343078 6010
rect 343130 5958 343142 6010
rect 343194 5958 343206 6010
rect 343258 5958 343270 6010
rect 343322 5958 343334 6010
rect 343386 5958 378822 6010
rect 378874 5958 378886 6010
rect 378938 5958 378950 6010
rect 379002 5958 379014 6010
rect 379066 5958 379078 6010
rect 379130 5958 379142 6010
rect 379194 5958 379206 6010
rect 379258 5958 379270 6010
rect 379322 5958 379334 6010
rect 379386 5958 414822 6010
rect 414874 5958 414886 6010
rect 414938 5958 414950 6010
rect 415002 5958 415014 6010
rect 415066 5958 415078 6010
rect 415130 5958 415142 6010
rect 415194 5958 415206 6010
rect 415258 5958 415270 6010
rect 415322 5958 415334 6010
rect 415386 5958 450822 6010
rect 450874 5958 450886 6010
rect 450938 5958 450950 6010
rect 451002 5958 451014 6010
rect 451066 5958 451078 6010
rect 451130 5958 451142 6010
rect 451194 5958 451206 6010
rect 451258 5958 451270 6010
rect 451322 5958 451334 6010
rect 451386 5958 486822 6010
rect 486874 5958 486886 6010
rect 486938 5958 486950 6010
rect 487002 5958 487014 6010
rect 487066 5958 487078 6010
rect 487130 5958 487142 6010
rect 487194 5958 487206 6010
rect 487258 5958 487270 6010
rect 487322 5958 487334 6010
rect 487386 5958 522822 6010
rect 522874 5958 522886 6010
rect 522938 5958 522950 6010
rect 523002 5958 523014 6010
rect 523066 5958 523078 6010
rect 523130 5958 523142 6010
rect 523194 5958 523206 6010
rect 523258 5958 523270 6010
rect 523322 5958 523334 6010
rect 523386 5958 558822 6010
rect 558874 5958 558886 6010
rect 558938 5958 558950 6010
rect 559002 5958 559014 6010
rect 559066 5958 559078 6010
rect 559130 5958 559142 6010
rect 559194 5958 559206 6010
rect 559258 5958 559270 6010
rect 559322 5958 559334 6010
rect 559386 5958 582820 6010
rect 1104 5936 582820 5958
rect 266998 5856 267004 5908
rect 267056 5896 267062 5908
rect 269666 5896 269672 5908
rect 267056 5868 269672 5896
rect 267056 5856 267062 5868
rect 269666 5856 269672 5868
rect 269724 5856 269730 5908
rect 315758 5856 315764 5908
rect 315816 5896 315822 5908
rect 318702 5896 318708 5908
rect 315816 5868 318708 5896
rect 315816 5856 315822 5868
rect 318702 5856 318708 5868
rect 318760 5856 318766 5908
rect 322566 5856 322572 5908
rect 322624 5896 322630 5908
rect 324314 5896 324320 5908
rect 322624 5868 324320 5896
rect 322624 5856 322630 5868
rect 324314 5856 324320 5868
rect 324372 5856 324378 5908
rect 324866 5856 324872 5908
rect 324924 5896 324930 5908
rect 328270 5896 328276 5908
rect 324924 5868 328276 5896
rect 324924 5856 324930 5868
rect 328270 5856 328276 5868
rect 328328 5856 328334 5908
rect 335078 5856 335084 5908
rect 335136 5896 335142 5908
rect 337378 5896 337384 5908
rect 335136 5868 337384 5896
rect 335136 5856 335142 5868
rect 337378 5856 337384 5868
rect 337436 5856 337442 5908
rect 408770 5856 408776 5908
rect 408828 5896 408834 5908
rect 418154 5896 418160 5908
rect 408828 5868 418160 5896
rect 408828 5856 408834 5868
rect 418154 5856 418160 5868
rect 418212 5856 418218 5908
rect 445018 5856 445024 5908
rect 445076 5896 445082 5908
rect 454678 5896 454684 5908
rect 445076 5868 454684 5896
rect 445076 5856 445082 5868
rect 454678 5856 454684 5868
rect 454736 5856 454742 5908
rect 459738 5856 459744 5908
rect 459796 5896 459802 5908
rect 469398 5896 469404 5908
rect 459796 5868 469404 5896
rect 459796 5856 459802 5868
rect 469398 5856 469404 5868
rect 469456 5856 469462 5908
rect 492674 5856 492680 5908
rect 492732 5896 492738 5908
rect 503990 5896 503996 5908
rect 492732 5868 503996 5896
rect 492732 5856 492738 5868
rect 503990 5856 503996 5868
rect 504048 5856 504054 5908
rect 510706 5856 510712 5908
rect 510764 5896 510770 5908
rect 522390 5896 522396 5908
rect 510764 5868 522396 5896
rect 510764 5856 510770 5868
rect 522390 5856 522396 5868
rect 522448 5856 522454 5908
rect 94498 5788 94504 5840
rect 94556 5828 94562 5840
rect 98086 5828 98092 5840
rect 94556 5800 98092 5828
rect 94556 5788 94562 5800
rect 98086 5788 98092 5800
rect 98144 5788 98150 5840
rect 238662 5788 238668 5840
rect 238720 5828 238726 5840
rect 240134 5828 240140 5840
rect 238720 5800 240140 5828
rect 238720 5788 238726 5800
rect 240134 5788 240140 5800
rect 240192 5788 240198 5840
rect 257982 5788 257988 5840
rect 258040 5828 258046 5840
rect 260098 5828 260104 5840
rect 258040 5800 260104 5828
rect 258040 5788 258046 5800
rect 260098 5788 260104 5800
rect 260156 5788 260162 5840
rect 265894 5788 265900 5840
rect 265952 5828 265958 5840
rect 269022 5828 269028 5840
rect 265952 5800 269028 5828
rect 265952 5788 265958 5800
rect 269022 5788 269028 5800
rect 269080 5788 269086 5840
rect 282914 5788 282920 5840
rect 282972 5828 282978 5840
rect 285766 5828 285772 5840
rect 282972 5800 285772 5828
rect 282972 5788 282978 5800
rect 285766 5788 285772 5800
rect 285824 5788 285830 5840
rect 286318 5788 286324 5840
rect 286376 5828 286382 5840
rect 289446 5828 289452 5840
rect 286376 5800 289452 5828
rect 286376 5788 286382 5800
rect 289446 5788 289452 5800
rect 289504 5788 289510 5840
rect 295334 5788 295340 5840
rect 295392 5828 295398 5840
rect 298922 5828 298928 5840
rect 295392 5800 298928 5828
rect 295392 5788 295398 5800
rect 298922 5788 298928 5800
rect 298980 5788 298986 5840
rect 301038 5788 301044 5840
rect 301096 5828 301102 5840
rect 303706 5828 303712 5840
rect 301096 5800 303712 5828
rect 301096 5788 301102 5800
rect 303706 5788 303712 5800
rect 303764 5788 303770 5840
rect 304442 5788 304448 5840
rect 304500 5828 304506 5840
rect 307662 5828 307668 5840
rect 304500 5800 307668 5828
rect 304500 5788 304506 5800
rect 307662 5788 307668 5800
rect 307720 5788 307726 5840
rect 321462 5788 321468 5840
rect 321520 5828 321526 5840
rect 323578 5828 323584 5840
rect 321520 5800 323584 5828
rect 321520 5788 321526 5800
rect 323578 5788 323584 5800
rect 323636 5788 323642 5840
rect 330478 5788 330484 5840
rect 330536 5828 330542 5840
rect 332962 5828 332968 5840
rect 330536 5800 332968 5828
rect 330536 5788 330542 5800
rect 332962 5788 332968 5800
rect 333020 5788 333026 5840
rect 344094 5788 344100 5840
rect 344152 5828 344158 5840
rect 347406 5828 347412 5840
rect 344152 5800 347412 5828
rect 344152 5788 344158 5800
rect 347406 5788 347412 5800
rect 347464 5788 347470 5840
rect 348694 5788 348700 5840
rect 348752 5828 348758 5840
rect 351730 5828 351736 5840
rect 348752 5800 351736 5828
rect 348752 5788 348758 5800
rect 351730 5788 351736 5800
rect 351788 5788 351794 5840
rect 380434 5788 380440 5840
rect 380492 5828 380498 5840
rect 382274 5828 382280 5840
rect 380492 5800 382280 5828
rect 380492 5788 380498 5800
rect 382274 5788 382280 5800
rect 382332 5788 382338 5840
rect 433702 5788 433708 5840
rect 433760 5828 433766 5840
rect 444374 5828 444380 5840
rect 433760 5800 444380 5828
rect 433760 5788 433766 5800
rect 444374 5788 444380 5800
rect 444432 5788 444438 5840
rect 469950 5788 469956 5840
rect 470008 5828 470014 5840
rect 478874 5828 478880 5840
rect 470008 5800 478880 5828
rect 470008 5788 470014 5800
rect 478874 5788 478880 5800
rect 478932 5788 478938 5840
rect 500494 5788 500500 5840
rect 500552 5828 500558 5840
rect 511902 5828 511908 5840
rect 500552 5800 511908 5828
rect 500552 5788 500558 5800
rect 511902 5788 511908 5800
rect 511960 5788 511966 5840
rect 513006 5788 513012 5840
rect 513064 5828 513070 5840
rect 529842 5828 529848 5840
rect 513064 5800 529848 5828
rect 513064 5788 513070 5800
rect 529842 5788 529848 5800
rect 529900 5788 529906 5840
rect 23842 5720 23848 5772
rect 23900 5760 23906 5772
rect 25498 5760 25504 5772
rect 23900 5732 25504 5760
rect 23900 5720 23906 5732
rect 25498 5720 25504 5732
rect 25556 5720 25562 5772
rect 79042 5720 79048 5772
rect 79100 5760 79106 5772
rect 83366 5760 83372 5772
rect 79100 5732 83372 5760
rect 79100 5720 79106 5732
rect 83366 5720 83372 5732
rect 83424 5720 83430 5772
rect 84930 5720 84936 5772
rect 84988 5760 84994 5772
rect 88978 5760 88984 5772
rect 84988 5732 88984 5760
rect 84988 5720 84994 5732
rect 88978 5720 88984 5732
rect 89036 5720 89042 5772
rect 89714 5720 89720 5772
rect 89772 5760 89778 5772
rect 93578 5760 93584 5772
rect 89772 5732 93584 5760
rect 89772 5720 89778 5732
rect 93578 5720 93584 5732
rect 93636 5720 93642 5772
rect 96890 5720 96896 5772
rect 96948 5760 96954 5772
rect 100386 5760 100392 5772
rect 96948 5732 100392 5760
rect 96948 5720 96954 5732
rect 100386 5720 100392 5732
rect 100444 5720 100450 5772
rect 105170 5720 105176 5772
rect 105228 5760 105234 5772
rect 108298 5760 108304 5772
rect 105228 5732 108304 5760
rect 105228 5720 105234 5732
rect 108298 5720 108304 5732
rect 108356 5720 108362 5772
rect 118234 5720 118240 5772
rect 118292 5760 118298 5772
rect 120810 5760 120816 5772
rect 118292 5732 120816 5760
rect 118292 5720 118298 5732
rect 120810 5720 120816 5732
rect 120868 5720 120874 5772
rect 226242 5720 226248 5772
rect 226300 5760 226306 5772
rect 228910 5760 228916 5772
rect 226300 5732 228916 5760
rect 226300 5720 226306 5732
rect 228910 5720 228916 5732
rect 228968 5720 228974 5772
rect 234154 5720 234160 5772
rect 234212 5760 234218 5772
rect 237190 5760 237196 5772
rect 234212 5732 237196 5760
rect 234212 5720 234218 5732
rect 237190 5720 237196 5732
rect 237248 5720 237254 5772
rect 243170 5720 243176 5772
rect 243228 5760 243234 5772
rect 246758 5760 246764 5772
rect 243228 5732 246764 5760
rect 243228 5720 243234 5732
rect 246758 5720 246764 5732
rect 246816 5720 246822 5772
rect 247770 5720 247776 5772
rect 247828 5760 247834 5772
rect 251082 5760 251088 5772
rect 247828 5732 251088 5760
rect 247828 5720 247834 5732
rect 251082 5720 251088 5732
rect 251140 5720 251146 5772
rect 252278 5720 252284 5772
rect 252336 5760 252342 5772
rect 254210 5760 254216 5772
rect 252336 5732 254216 5760
rect 252336 5720 252342 5732
rect 254210 5720 254216 5732
rect 254268 5720 254274 5772
rect 277210 5720 277216 5772
rect 277268 5760 277274 5772
rect 279786 5760 279792 5772
rect 277268 5732 279792 5760
rect 277268 5720 277274 5732
rect 279786 5720 279792 5732
rect 279844 5720 279850 5772
rect 280614 5720 280620 5772
rect 280672 5760 280678 5772
rect 283190 5760 283196 5772
rect 280672 5732 283196 5760
rect 280672 5720 280678 5732
rect 283190 5720 283196 5732
rect 283248 5720 283254 5772
rect 289722 5720 289728 5772
rect 289780 5760 289786 5772
rect 292482 5760 292488 5772
rect 289780 5732 292488 5760
rect 289780 5720 289786 5732
rect 292482 5720 292488 5732
rect 292540 5720 292546 5772
rect 308950 5720 308956 5772
rect 309008 5760 309014 5772
rect 311802 5760 311808 5772
rect 309008 5732 311808 5760
rect 309008 5720 309014 5732
rect 311802 5720 311808 5732
rect 311860 5720 311866 5772
rect 323670 5720 323676 5772
rect 323728 5760 323734 5772
rect 326982 5760 326988 5772
rect 323728 5732 326988 5760
rect 323728 5720 323734 5732
rect 326982 5720 326988 5732
rect 327040 5720 327046 5772
rect 410978 5720 410984 5772
rect 411036 5760 411042 5772
rect 413922 5760 413928 5772
rect 411036 5732 413928 5760
rect 411036 5720 411042 5732
rect 413922 5720 413928 5732
rect 413980 5720 413986 5772
rect 490374 5720 490380 5772
rect 490432 5760 490438 5772
rect 506014 5760 506020 5772
rect 490432 5732 506020 5760
rect 490432 5720 490438 5732
rect 506014 5720 506020 5732
rect 506072 5720 506078 5772
rect 15194 5652 15200 5704
rect 15252 5692 15258 5704
rect 17586 5692 17592 5704
rect 15252 5664 17592 5692
rect 15252 5652 15258 5664
rect 17586 5652 17592 5664
rect 17644 5652 17650 5704
rect 18598 5652 18604 5704
rect 18656 5692 18662 5704
rect 20990 5692 20996 5704
rect 18656 5664 20996 5692
rect 18656 5652 18662 5664
rect 20990 5652 20996 5664
rect 21048 5652 21054 5704
rect 23106 5652 23112 5704
rect 23164 5692 23170 5704
rect 24394 5692 24400 5704
rect 23164 5664 24400 5692
rect 23164 5652 23170 5664
rect 24394 5652 24400 5664
rect 24452 5652 24458 5704
rect 26234 5652 26240 5704
rect 26292 5692 26298 5704
rect 28902 5692 28908 5704
rect 26292 5664 28908 5692
rect 26292 5652 26298 5664
rect 28902 5652 28908 5664
rect 28960 5652 28966 5704
rect 75454 5652 75460 5704
rect 75512 5692 75518 5704
rect 79962 5692 79968 5704
rect 75512 5664 79968 5692
rect 75512 5652 75518 5664
rect 79962 5652 79968 5664
rect 80020 5652 80026 5704
rect 80238 5652 80244 5704
rect 80296 5692 80302 5704
rect 84470 5692 84476 5704
rect 80296 5664 84476 5692
rect 80296 5652 80302 5664
rect 84470 5652 84476 5664
rect 84528 5652 84534 5704
rect 88518 5652 88524 5704
rect 88576 5692 88582 5704
rect 92382 5692 92388 5704
rect 88576 5664 92388 5692
rect 88576 5652 88582 5664
rect 92382 5652 92388 5664
rect 92440 5652 92446 5704
rect 95694 5652 95700 5704
rect 95752 5692 95758 5704
rect 99190 5692 99196 5704
rect 95752 5664 99196 5692
rect 95752 5652 95758 5664
rect 99190 5652 99196 5664
rect 99248 5652 99254 5704
rect 100478 5652 100484 5704
rect 100536 5692 100542 5704
rect 103790 5692 103796 5704
rect 100536 5664 103796 5692
rect 100536 5652 100542 5664
rect 103790 5652 103796 5664
rect 103848 5652 103854 5704
rect 103974 5652 103980 5704
rect 104032 5692 104038 5704
rect 107194 5692 107200 5704
rect 104032 5664 107200 5692
rect 104032 5652 104038 5664
rect 107194 5652 107200 5664
rect 107252 5652 107258 5704
rect 107562 5652 107568 5704
rect 107620 5692 107626 5704
rect 110598 5692 110604 5704
rect 107620 5664 110604 5692
rect 107620 5652 107626 5664
rect 110598 5652 110604 5664
rect 110656 5652 110662 5704
rect 111150 5652 111156 5704
rect 111208 5692 111214 5704
rect 114002 5692 114008 5704
rect 111208 5664 114008 5692
rect 111208 5652 111214 5664
rect 114002 5652 114008 5664
rect 114060 5652 114066 5704
rect 114738 5652 114744 5704
rect 114796 5692 114802 5704
rect 117406 5692 117412 5704
rect 114796 5664 117412 5692
rect 114796 5652 114802 5664
rect 117406 5652 117412 5664
rect 117464 5652 117470 5704
rect 120626 5652 120632 5704
rect 120684 5692 120690 5704
rect 123018 5692 123024 5704
rect 120684 5664 123024 5692
rect 120684 5652 120690 5664
rect 123018 5652 123024 5664
rect 123076 5652 123082 5704
rect 132586 5652 132592 5704
rect 132644 5692 132650 5704
rect 134334 5692 134340 5704
rect 132644 5664 134340 5692
rect 132644 5652 132650 5664
rect 134334 5652 134340 5664
rect 134392 5652 134398 5704
rect 143258 5652 143264 5704
rect 143316 5692 143322 5704
rect 144546 5692 144552 5704
rect 143316 5664 144552 5692
rect 143316 5652 143322 5664
rect 144546 5652 144552 5664
rect 144604 5652 144610 5704
rect 145650 5652 145656 5704
rect 145708 5692 145714 5704
rect 146846 5692 146852 5704
rect 145708 5664 146852 5692
rect 145708 5652 145714 5664
rect 146846 5652 146852 5664
rect 146904 5652 146910 5704
rect 195606 5652 195612 5704
rect 195664 5692 195670 5704
rect 196802 5692 196808 5704
rect 195664 5664 196808 5692
rect 195664 5652 195670 5664
rect 196802 5652 196808 5664
rect 196860 5652 196866 5704
rect 206922 5652 206928 5704
rect 206980 5692 206986 5704
rect 208670 5692 208676 5704
rect 206980 5664 208676 5692
rect 206980 5652 206986 5664
rect 208670 5652 208676 5664
rect 208728 5652 208734 5704
rect 214834 5652 214840 5704
rect 214892 5692 214898 5704
rect 216674 5692 216680 5704
rect 214892 5664 216680 5692
rect 214892 5652 214898 5664
rect 216674 5652 216680 5664
rect 216732 5652 216738 5704
rect 220538 5652 220544 5704
rect 220596 5692 220602 5704
rect 222930 5692 222936 5704
rect 220596 5664 222936 5692
rect 220596 5652 220602 5664
rect 222930 5652 222936 5664
rect 222988 5652 222994 5704
rect 223942 5652 223948 5704
rect 224000 5692 224006 5704
rect 226518 5692 226524 5704
rect 224000 5664 226524 5692
rect 224000 5652 224006 5664
rect 226518 5652 226524 5664
rect 226576 5652 226582 5704
rect 228450 5652 228456 5704
rect 228508 5692 228514 5704
rect 231302 5692 231308 5704
rect 228508 5664 231308 5692
rect 228508 5652 228514 5664
rect 231302 5652 231308 5664
rect 231360 5652 231366 5704
rect 231854 5652 231860 5704
rect 231912 5692 231918 5704
rect 234706 5692 234712 5704
rect 231912 5664 234712 5692
rect 231912 5652 231918 5664
rect 234706 5652 234712 5664
rect 234764 5652 234770 5704
rect 242066 5652 242072 5704
rect 242124 5692 242130 5704
rect 245562 5692 245568 5704
rect 242124 5664 245568 5692
rect 242124 5652 242130 5664
rect 245562 5652 245568 5664
rect 245620 5652 245626 5704
rect 249978 5652 249984 5704
rect 250036 5692 250042 5704
rect 253842 5692 253848 5704
rect 250036 5664 253848 5692
rect 250036 5652 250042 5664
rect 253842 5652 253848 5664
rect 253900 5652 253906 5704
rect 260190 5652 260196 5704
rect 260248 5692 260254 5704
rect 262398 5692 262404 5704
rect 260248 5664 262404 5692
rect 260248 5652 260254 5664
rect 262398 5652 262404 5664
rect 262456 5652 262462 5704
rect 262490 5652 262496 5704
rect 262548 5692 262554 5704
rect 264974 5692 264980 5704
rect 262548 5664 264980 5692
rect 262548 5652 262554 5664
rect 264974 5652 264980 5664
rect 265032 5652 265038 5704
rect 270402 5652 270408 5704
rect 270460 5692 270466 5704
rect 272978 5692 272984 5704
rect 270460 5664 272984 5692
rect 270460 5652 270466 5664
rect 272978 5652 272984 5664
rect 273036 5652 273042 5704
rect 276106 5652 276112 5704
rect 276164 5692 276170 5704
rect 279326 5692 279332 5704
rect 276164 5664 279332 5692
rect 276164 5652 276170 5664
rect 279326 5652 279332 5664
rect 279384 5652 279390 5704
rect 281718 5652 281724 5704
rect 281776 5692 281782 5704
rect 284386 5692 284392 5704
rect 281776 5664 284392 5692
rect 281776 5652 281782 5664
rect 284386 5652 284392 5664
rect 284444 5652 284450 5704
rect 291930 5652 291936 5704
rect 291988 5692 291994 5704
rect 294322 5692 294328 5704
rect 291988 5664 294328 5692
rect 291988 5652 291994 5664
rect 294322 5652 294328 5664
rect 294380 5652 294386 5704
rect 296530 5652 296536 5704
rect 296588 5692 296594 5704
rect 299198 5692 299204 5704
rect 296588 5664 299204 5692
rect 296588 5652 296594 5664
rect 299198 5652 299204 5664
rect 299256 5652 299262 5704
rect 299934 5652 299940 5704
rect 299992 5692 299998 5704
rect 303062 5692 303068 5704
rect 299992 5664 303068 5692
rect 299992 5652 299998 5664
rect 303062 5652 303068 5664
rect 303120 5652 303126 5704
rect 303338 5652 303344 5704
rect 303396 5692 303402 5704
rect 304994 5692 305000 5704
rect 303396 5664 305000 5692
rect 303396 5652 303402 5664
rect 304994 5652 305000 5664
rect 305052 5652 305058 5704
rect 305546 5652 305552 5704
rect 305604 5692 305610 5704
rect 308214 5692 308220 5704
rect 305604 5664 308220 5692
rect 305604 5652 305610 5664
rect 308214 5652 308220 5664
rect 308272 5652 308278 5704
rect 310146 5652 310152 5704
rect 310204 5692 310210 5704
rect 313090 5692 313096 5704
rect 310204 5664 313096 5692
rect 310204 5652 310210 5664
rect 313090 5652 313096 5664
rect 313148 5652 313154 5704
rect 318058 5652 318064 5704
rect 318116 5692 318122 5704
rect 321462 5692 321468 5704
rect 318116 5664 321468 5692
rect 318116 5652 318122 5664
rect 321462 5652 321468 5664
rect 321520 5652 321526 5704
rect 329374 5652 329380 5704
rect 329432 5692 329438 5704
rect 332410 5692 332416 5704
rect 329432 5664 332416 5692
rect 329432 5652 329438 5664
rect 332410 5652 332416 5664
rect 332468 5652 332474 5704
rect 338482 5652 338488 5704
rect 338540 5692 338546 5704
rect 341794 5692 341800 5704
rect 338540 5664 341800 5692
rect 338540 5652 338546 5664
rect 341794 5652 341800 5664
rect 341852 5652 341858 5704
rect 341886 5652 341892 5704
rect 341944 5692 341950 5704
rect 343634 5692 343640 5704
rect 341944 5664 343640 5692
rect 341944 5652 341950 5664
rect 343634 5652 343640 5664
rect 343692 5652 343698 5704
rect 349798 5652 349804 5704
rect 349856 5692 349862 5704
rect 352282 5692 352288 5704
rect 349856 5664 352288 5692
rect 349856 5652 349862 5664
rect 352282 5652 352288 5664
rect 352340 5652 352346 5704
rect 357710 5652 357716 5704
rect 357768 5692 357774 5704
rect 360746 5692 360752 5704
rect 357768 5664 360752 5692
rect 357768 5652 357774 5664
rect 360746 5652 360752 5664
rect 360804 5652 360810 5704
rect 381538 5652 381544 5704
rect 381596 5692 381602 5704
rect 384942 5692 384948 5704
rect 381596 5664 384948 5692
rect 381596 5652 381602 5664
rect 384942 5652 384948 5664
rect 385000 5652 385006 5704
rect 409874 5652 409880 5704
rect 409932 5692 409938 5704
rect 413370 5692 413376 5704
rect 409932 5664 413376 5692
rect 409932 5652 409938 5664
rect 413370 5652 413376 5664
rect 413428 5652 413434 5704
rect 440510 5652 440516 5704
rect 440568 5692 440574 5704
rect 444282 5692 444288 5704
rect 440568 5664 444288 5692
rect 440568 5652 440574 5664
rect 444282 5652 444288 5664
rect 444340 5652 444346 5704
rect 13814 5584 13820 5636
rect 13872 5624 13878 5636
rect 16482 5624 16488 5636
rect 13872 5596 16488 5624
rect 13872 5584 13878 5596
rect 16482 5584 16488 5596
rect 16540 5584 16546 5636
rect 18046 5584 18052 5636
rect 18104 5624 18110 5636
rect 19886 5624 19892 5636
rect 18104 5596 19892 5624
rect 18104 5584 18110 5596
rect 19886 5584 19892 5596
rect 19944 5584 19950 5636
rect 20714 5584 20720 5636
rect 20772 5624 20778 5636
rect 23290 5624 23296 5636
rect 20772 5596 23296 5624
rect 20772 5584 20778 5596
rect 23290 5584 23296 5596
rect 23348 5584 23354 5636
rect 27706 5584 27712 5636
rect 27764 5624 27770 5636
rect 30098 5624 30104 5636
rect 27764 5596 30104 5624
rect 27764 5584 27770 5596
rect 30098 5584 30104 5596
rect 30156 5584 30162 5636
rect 34514 5584 34520 5636
rect 34572 5624 34578 5636
rect 36906 5624 36912 5636
rect 34572 5596 36912 5624
rect 34572 5584 34578 5596
rect 36906 5584 36912 5596
rect 36964 5584 36970 5636
rect 37458 5584 37464 5636
rect 37516 5624 37522 5636
rect 39114 5624 39120 5636
rect 37516 5596 39120 5624
rect 37516 5584 37522 5596
rect 39114 5584 39120 5596
rect 39172 5584 39178 5636
rect 69474 5584 69480 5636
rect 69532 5624 69538 5636
rect 74258 5624 74264 5636
rect 69532 5596 74264 5624
rect 69532 5584 69538 5596
rect 74258 5584 74264 5596
rect 74316 5584 74322 5636
rect 77846 5584 77852 5636
rect 77904 5624 77910 5636
rect 82262 5624 82268 5636
rect 77904 5596 82268 5624
rect 77904 5584 77910 5596
rect 82262 5584 82268 5596
rect 82320 5584 82326 5636
rect 82630 5584 82636 5636
rect 82688 5624 82694 5636
rect 86770 5624 86776 5636
rect 82688 5596 86776 5624
rect 82688 5584 82694 5596
rect 86770 5584 86776 5596
rect 86828 5584 86834 5636
rect 90726 5584 90732 5636
rect 90784 5624 90790 5636
rect 94682 5624 94688 5636
rect 90784 5596 94688 5624
rect 90784 5584 90790 5596
rect 94682 5584 94688 5596
rect 94740 5584 94746 5636
rect 98086 5584 98092 5636
rect 98144 5624 98150 5636
rect 101490 5624 101496 5636
rect 98144 5596 101496 5624
rect 98144 5584 98150 5596
rect 101490 5584 101496 5596
rect 101548 5584 101554 5636
rect 101582 5584 101588 5636
rect 101640 5624 101646 5636
rect 104894 5624 104900 5636
rect 101640 5596 104900 5624
rect 101640 5584 101646 5596
rect 104894 5584 104900 5596
rect 104952 5584 104958 5636
rect 106366 5584 106372 5636
rect 106424 5624 106430 5636
rect 109402 5624 109408 5636
rect 106424 5596 109408 5624
rect 106424 5584 106430 5596
rect 109402 5584 109408 5596
rect 109460 5584 109466 5636
rect 109954 5584 109960 5636
rect 110012 5624 110018 5636
rect 112806 5624 112812 5636
rect 110012 5596 112812 5624
rect 110012 5584 110018 5596
rect 112806 5584 112812 5596
rect 112864 5584 112870 5636
rect 113542 5584 113548 5636
rect 113600 5624 113606 5636
rect 116210 5624 116216 5636
rect 113600 5596 116216 5624
rect 113600 5584 113606 5596
rect 116210 5584 116216 5596
rect 116268 5584 116274 5636
rect 117130 5584 117136 5636
rect 117188 5624 117194 5636
rect 119614 5624 119620 5636
rect 117188 5596 119620 5624
rect 117188 5584 117194 5596
rect 119614 5584 119620 5596
rect 119672 5584 119678 5636
rect 121822 5584 121828 5636
rect 121880 5624 121886 5636
rect 124122 5624 124128 5636
rect 121880 5596 124128 5624
rect 121880 5584 121886 5596
rect 124122 5584 124128 5596
rect 124180 5584 124186 5636
rect 124214 5584 124220 5636
rect 124272 5624 124278 5636
rect 126422 5624 126428 5636
rect 124272 5596 126428 5624
rect 124272 5584 124278 5596
rect 126422 5584 126428 5596
rect 126480 5584 126486 5636
rect 126606 5584 126612 5636
rect 126664 5624 126670 5636
rect 128722 5624 128728 5636
rect 126664 5596 128728 5624
rect 126664 5584 126670 5596
rect 128722 5584 128728 5596
rect 128780 5584 128786 5636
rect 128998 5584 129004 5636
rect 129056 5624 129062 5636
rect 130930 5624 130936 5636
rect 129056 5596 130936 5624
rect 129056 5584 129062 5596
rect 130930 5584 130936 5596
rect 130988 5584 130994 5636
rect 131390 5584 131396 5636
rect 131448 5624 131454 5636
rect 133230 5624 133236 5636
rect 131448 5596 133236 5624
rect 131448 5584 131454 5596
rect 133230 5584 133236 5596
rect 133288 5584 133294 5636
rect 134886 5584 134892 5636
rect 134944 5624 134950 5636
rect 136634 5624 136640 5636
rect 134944 5596 136640 5624
rect 134944 5584 134950 5596
rect 136634 5584 136640 5596
rect 136692 5584 136698 5636
rect 137278 5584 137284 5636
rect 137336 5624 137342 5636
rect 138934 5624 138940 5636
rect 137336 5596 138940 5624
rect 137336 5584 137342 5596
rect 138934 5584 138940 5596
rect 138992 5584 138998 5636
rect 139670 5584 139676 5636
rect 139728 5624 139734 5636
rect 141142 5624 141148 5636
rect 139728 5596 141148 5624
rect 139728 5584 139734 5596
rect 141142 5584 141148 5596
rect 141200 5584 141206 5636
rect 142062 5584 142068 5636
rect 142120 5624 142126 5636
rect 143442 5624 143448 5636
rect 142120 5596 143448 5624
rect 142120 5584 142126 5596
rect 143442 5584 143448 5596
rect 143500 5584 143506 5636
rect 197906 5584 197912 5636
rect 197964 5624 197970 5636
rect 198734 5624 198740 5636
rect 197964 5596 198740 5624
rect 197964 5584 197970 5596
rect 198734 5584 198740 5596
rect 198792 5584 198798 5636
rect 201218 5584 201224 5636
rect 201276 5624 201282 5636
rect 202690 5624 202696 5636
rect 201276 5596 202696 5624
rect 201276 5584 201282 5596
rect 202690 5584 202696 5596
rect 202748 5584 202754 5636
rect 203518 5584 203524 5636
rect 203576 5624 203582 5636
rect 205082 5624 205088 5636
rect 203576 5596 205088 5624
rect 203576 5584 203582 5596
rect 205082 5584 205088 5596
rect 205140 5584 205146 5636
rect 205818 5584 205824 5636
rect 205876 5624 205882 5636
rect 207474 5624 207480 5636
rect 205876 5596 207480 5624
rect 205876 5584 205882 5596
rect 207474 5584 207480 5596
rect 207532 5584 207538 5636
rect 209222 5584 209228 5636
rect 209280 5624 209286 5636
rect 211062 5624 211068 5636
rect 209280 5596 211068 5624
rect 209280 5584 209286 5596
rect 211062 5584 211068 5596
rect 211120 5584 211126 5636
rect 211430 5584 211436 5636
rect 211488 5624 211494 5636
rect 213454 5624 213460 5636
rect 211488 5596 213460 5624
rect 211488 5584 211494 5596
rect 213454 5584 213460 5596
rect 213512 5584 213518 5636
rect 213730 5584 213736 5636
rect 213788 5624 213794 5636
rect 215846 5624 215852 5636
rect 213788 5596 215852 5624
rect 213788 5584 213794 5596
rect 215846 5584 215852 5596
rect 215904 5584 215910 5636
rect 217134 5584 217140 5636
rect 217192 5624 217198 5636
rect 219342 5624 219348 5636
rect 217192 5596 219348 5624
rect 217192 5584 217198 5596
rect 219342 5584 219348 5596
rect 219400 5584 219406 5636
rect 219434 5584 219440 5636
rect 219492 5624 219498 5636
rect 221734 5624 221740 5636
rect 219492 5596 221740 5624
rect 219492 5584 219498 5596
rect 221734 5584 221740 5596
rect 221792 5584 221798 5636
rect 222838 5584 222844 5636
rect 222896 5624 222902 5636
rect 225322 5624 225328 5636
rect 222896 5596 225328 5624
rect 222896 5584 222902 5596
rect 225322 5584 225328 5596
rect 225380 5584 225386 5636
rect 227346 5584 227352 5636
rect 227404 5624 227410 5636
rect 230106 5624 230112 5636
rect 227404 5596 230112 5624
rect 227404 5584 227410 5596
rect 230106 5584 230112 5596
rect 230164 5584 230170 5636
rect 230750 5584 230756 5636
rect 230808 5624 230814 5636
rect 233694 5624 233700 5636
rect 230808 5596 233700 5624
rect 230808 5584 230814 5596
rect 233694 5584 233700 5596
rect 233752 5584 233758 5636
rect 236362 5584 236368 5636
rect 236420 5624 236426 5636
rect 239582 5624 239588 5636
rect 236420 5596 239588 5624
rect 236420 5584 236426 5596
rect 239582 5584 239588 5596
rect 239640 5584 239646 5636
rect 239766 5584 239772 5636
rect 239824 5624 239830 5636
rect 242802 5624 242808 5636
rect 239824 5596 242808 5624
rect 239824 5584 239830 5596
rect 242802 5584 242808 5596
rect 242860 5584 242866 5636
rect 244366 5584 244372 5636
rect 244424 5624 244430 5636
rect 247954 5624 247960 5636
rect 244424 5596 247960 5624
rect 244424 5584 244430 5596
rect 247954 5584 247960 5596
rect 248012 5584 248018 5636
rect 248874 5584 248880 5636
rect 248932 5624 248938 5636
rect 252462 5624 252468 5636
rect 248932 5596 252468 5624
rect 248932 5584 248938 5596
rect 252462 5584 252468 5596
rect 252520 5584 252526 5636
rect 253382 5584 253388 5636
rect 253440 5624 253446 5636
rect 255406 5624 255412 5636
rect 253440 5596 255412 5624
rect 253440 5584 253446 5596
rect 255406 5584 255412 5596
rect 255464 5584 255470 5636
rect 256786 5584 256792 5636
rect 256844 5624 256850 5636
rect 260742 5624 260748 5636
rect 256844 5596 260748 5624
rect 256844 5584 256850 5596
rect 260742 5584 260748 5596
rect 260800 5584 260806 5636
rect 261386 5584 261392 5636
rect 261444 5624 261450 5636
rect 263686 5624 263692 5636
rect 261444 5596 263692 5624
rect 261444 5584 261450 5596
rect 263686 5584 263692 5596
rect 263744 5584 263750 5636
rect 269298 5584 269304 5636
rect 269356 5624 269362 5636
rect 271874 5624 271880 5636
rect 269356 5596 271880 5624
rect 269356 5584 269362 5596
rect 271874 5584 271880 5596
rect 271932 5584 271938 5636
rect 278314 5584 278320 5636
rect 278372 5624 278378 5636
rect 280890 5624 280896 5636
rect 278372 5596 280896 5624
rect 278372 5584 278378 5596
rect 280890 5584 280896 5596
rect 280948 5584 280954 5636
rect 287422 5584 287428 5636
rect 287480 5624 287486 5636
rect 290182 5624 290188 5636
rect 287480 5596 290188 5624
rect 287480 5584 287486 5596
rect 290182 5584 290188 5596
rect 290240 5584 290246 5636
rect 297634 5584 297640 5636
rect 297692 5624 297698 5636
rect 300670 5624 300676 5636
rect 297692 5596 300676 5624
rect 297692 5584 297698 5596
rect 300670 5584 300676 5596
rect 300728 5584 300734 5636
rect 307846 5584 307852 5636
rect 307904 5624 307910 5636
rect 311158 5624 311164 5636
rect 307904 5596 311164 5624
rect 307904 5584 307910 5596
rect 311158 5584 311164 5596
rect 311216 5584 311222 5636
rect 312354 5584 312360 5636
rect 312412 5624 312418 5636
rect 314654 5624 314660 5636
rect 312412 5596 314660 5624
rect 312412 5584 312418 5596
rect 314654 5584 314660 5596
rect 314712 5584 314718 5636
rect 316862 5584 316868 5636
rect 316920 5624 316926 5636
rect 320082 5624 320088 5636
rect 316920 5596 320088 5624
rect 316920 5584 316926 5596
rect 320082 5584 320088 5596
rect 320140 5584 320146 5636
rect 327074 5584 327080 5636
rect 327132 5624 327138 5636
rect 330846 5624 330852 5636
rect 327132 5596 330852 5624
rect 327132 5584 327138 5596
rect 330846 5584 330852 5596
rect 330904 5584 330910 5636
rect 333882 5584 333888 5636
rect 333940 5624 333946 5636
rect 336642 5624 336648 5636
rect 333940 5596 336648 5624
rect 333940 5584 333946 5596
rect 336642 5584 336648 5596
rect 336700 5584 336706 5636
rect 345290 5584 345296 5636
rect 345348 5624 345354 5636
rect 348970 5624 348976 5636
rect 345348 5596 348976 5624
rect 345348 5584 345354 5596
rect 348970 5584 348976 5596
rect 349028 5584 349034 5636
rect 350902 5584 350908 5636
rect 350960 5624 350966 5636
rect 353294 5624 353300 5636
rect 350960 5596 353300 5624
rect 350960 5584 350966 5596
rect 353294 5584 353300 5596
rect 353352 5584 353358 5636
rect 365622 5584 365628 5636
rect 365680 5624 365686 5636
rect 367094 5624 367100 5636
rect 365680 5596 367100 5624
rect 365680 5584 365686 5596
rect 367094 5584 367100 5596
rect 367152 5584 367158 5636
rect 488074 5584 488080 5636
rect 488132 5624 488138 5636
rect 491202 5624 491208 5636
rect 488132 5596 491208 5624
rect 488132 5584 488138 5596
rect 491202 5584 491208 5596
rect 491260 5584 491266 5636
rect 11054 5516 11060 5568
rect 11112 5556 11118 5568
rect 14182 5556 14188 5568
rect 11112 5528 14188 5556
rect 11112 5516 11118 5528
rect 14182 5516 14188 5528
rect 14240 5516 14246 5568
rect 16942 5516 16948 5568
rect 17000 5556 17006 5568
rect 18690 5556 18696 5568
rect 17000 5528 18696 5556
rect 17000 5516 17006 5528
rect 18690 5516 18696 5528
rect 18748 5516 18754 5568
rect 19426 5516 19432 5568
rect 19484 5556 19490 5568
rect 22094 5556 22100 5568
rect 19484 5528 22100 5556
rect 19484 5516 19490 5528
rect 22094 5516 22100 5528
rect 22152 5516 22158 5568
rect 28994 5516 29000 5568
rect 29052 5556 29058 5568
rect 31202 5556 31208 5568
rect 29052 5528 31208 5556
rect 29052 5516 29058 5528
rect 31202 5516 31208 5528
rect 31260 5516 31266 5568
rect 31754 5516 31760 5568
rect 31812 5556 31818 5568
rect 33134 5556 33140 5568
rect 31812 5528 33140 5556
rect 31812 5516 31818 5528
rect 33134 5516 33140 5528
rect 33192 5516 33198 5568
rect 36446 5516 36452 5568
rect 36504 5556 36510 5568
rect 38010 5556 38016 5568
rect 36504 5528 38016 5556
rect 36504 5516 36510 5528
rect 38010 5516 38016 5528
rect 38068 5516 38074 5568
rect 42794 5516 42800 5568
rect 42852 5556 42858 5568
rect 44818 5556 44824 5568
rect 42852 5528 44824 5556
rect 42852 5516 42858 5528
rect 44818 5516 44824 5528
rect 44876 5516 44882 5568
rect 55398 5516 55404 5568
rect 55456 5556 55462 5568
rect 60642 5556 60648 5568
rect 55456 5528 60648 5556
rect 55456 5516 55462 5528
rect 60642 5516 60648 5528
rect 60700 5516 60706 5568
rect 62390 5516 62396 5568
rect 62448 5556 62454 5568
rect 67450 5556 67456 5568
rect 62448 5528 67456 5556
rect 62448 5516 62454 5528
rect 67450 5516 67456 5528
rect 67508 5516 67514 5568
rect 71866 5516 71872 5568
rect 71924 5556 71930 5568
rect 76558 5556 76564 5568
rect 71924 5528 76564 5556
rect 71924 5516 71930 5528
rect 76558 5516 76564 5528
rect 76616 5516 76622 5568
rect 76650 5516 76656 5568
rect 76708 5556 76714 5568
rect 81066 5556 81072 5568
rect 76708 5528 81072 5556
rect 76708 5516 76714 5528
rect 81066 5516 81072 5528
rect 81124 5516 81130 5568
rect 81434 5516 81440 5568
rect 81492 5556 81498 5568
rect 85574 5556 85580 5568
rect 81492 5528 85580 5556
rect 81492 5516 81498 5528
rect 85574 5516 85580 5528
rect 85632 5516 85638 5568
rect 86126 5516 86132 5568
rect 86184 5556 86190 5568
rect 90174 5556 90180 5568
rect 86184 5528 90180 5556
rect 86184 5516 86190 5528
rect 90174 5516 90180 5528
rect 90232 5516 90238 5568
rect 92106 5516 92112 5568
rect 92164 5556 92170 5568
rect 95786 5556 95792 5568
rect 92164 5528 95792 5556
rect 92164 5516 92170 5528
rect 95786 5516 95792 5528
rect 95844 5516 95850 5568
rect 99282 5516 99288 5568
rect 99340 5556 99346 5568
rect 102594 5556 102600 5568
rect 99340 5528 102600 5556
rect 99340 5516 99346 5528
rect 102594 5516 102600 5528
rect 102652 5516 102658 5568
rect 102778 5516 102784 5568
rect 102836 5556 102842 5568
rect 105998 5556 106004 5568
rect 102836 5528 106004 5556
rect 102836 5516 102842 5528
rect 105998 5516 106004 5528
rect 106056 5516 106062 5568
rect 108666 5516 108672 5568
rect 108724 5556 108730 5568
rect 111702 5556 111708 5568
rect 108724 5528 111708 5556
rect 108724 5516 108730 5528
rect 111702 5516 111708 5528
rect 111760 5516 111766 5568
rect 112346 5516 112352 5568
rect 112404 5556 112410 5568
rect 115106 5556 115112 5568
rect 112404 5528 115112 5556
rect 112404 5516 112410 5528
rect 115106 5516 115112 5528
rect 115164 5516 115170 5568
rect 115934 5516 115940 5568
rect 115992 5556 115998 5568
rect 118510 5556 118516 5568
rect 115992 5528 118516 5556
rect 115992 5516 115998 5528
rect 118510 5516 118516 5528
rect 118568 5516 118574 5568
rect 119430 5516 119436 5568
rect 119488 5556 119494 5568
rect 121914 5556 121920 5568
rect 119488 5528 121920 5556
rect 119488 5516 119494 5528
rect 121914 5516 121920 5528
rect 121972 5516 121978 5568
rect 123018 5516 123024 5568
rect 123076 5556 123082 5568
rect 125318 5556 125324 5568
rect 123076 5528 125324 5556
rect 123076 5516 123082 5528
rect 125318 5516 125324 5528
rect 125376 5516 125382 5568
rect 125410 5516 125416 5568
rect 125468 5556 125474 5568
rect 127526 5556 127532 5568
rect 125468 5528 127532 5556
rect 125468 5516 125474 5528
rect 127526 5516 127532 5528
rect 127584 5516 127590 5568
rect 127802 5516 127808 5568
rect 127860 5556 127866 5568
rect 129826 5556 129832 5568
rect 127860 5528 129832 5556
rect 127860 5516 127866 5528
rect 129826 5516 129832 5528
rect 129884 5516 129890 5568
rect 130194 5516 130200 5568
rect 130252 5556 130258 5568
rect 132126 5556 132132 5568
rect 130252 5528 132132 5556
rect 130252 5516 130258 5528
rect 132126 5516 132132 5528
rect 132184 5516 132190 5568
rect 133782 5516 133788 5568
rect 133840 5556 133846 5568
rect 135530 5556 135536 5568
rect 133840 5528 135536 5556
rect 133840 5516 133846 5528
rect 135530 5516 135536 5528
rect 135588 5516 135594 5568
rect 136082 5516 136088 5568
rect 136140 5556 136146 5568
rect 137738 5556 137744 5568
rect 136140 5528 137744 5556
rect 136140 5516 136146 5528
rect 137738 5516 137744 5528
rect 137796 5516 137802 5568
rect 138474 5516 138480 5568
rect 138532 5556 138538 5568
rect 140038 5556 140044 5568
rect 138532 5528 140044 5556
rect 138532 5516 138538 5528
rect 140038 5516 140044 5528
rect 140096 5516 140102 5568
rect 140866 5516 140872 5568
rect 140924 5556 140930 5568
rect 142338 5556 142344 5568
rect 140924 5528 142344 5556
rect 140924 5516 140930 5528
rect 142338 5516 142344 5528
rect 142396 5516 142402 5568
rect 144454 5516 144460 5568
rect 144512 5556 144518 5568
rect 145742 5556 145748 5568
rect 144512 5528 145748 5556
rect 144512 5516 144518 5528
rect 145742 5516 145748 5528
rect 145800 5516 145806 5568
rect 146846 5516 146852 5568
rect 146904 5556 146910 5568
rect 147950 5556 147956 5568
rect 146904 5528 147956 5556
rect 146904 5516 146910 5528
rect 147950 5516 147956 5528
rect 148008 5516 148014 5568
rect 148042 5516 148048 5568
rect 148100 5556 148106 5568
rect 149146 5556 149152 5568
rect 148100 5528 149152 5556
rect 148100 5516 148106 5528
rect 149146 5516 149152 5528
rect 149204 5516 149210 5568
rect 151538 5516 151544 5568
rect 151596 5556 151602 5568
rect 152550 5556 152556 5568
rect 151596 5528 152556 5556
rect 151596 5516 151602 5528
rect 152550 5516 152556 5528
rect 152608 5516 152614 5568
rect 152734 5516 152740 5568
rect 152792 5556 152798 5568
rect 153654 5556 153660 5568
rect 152792 5528 153660 5556
rect 152792 5516 152798 5528
rect 153654 5516 153660 5528
rect 153712 5516 153718 5568
rect 153930 5516 153936 5568
rect 153988 5556 153994 5568
rect 154758 5556 154764 5568
rect 153988 5528 154764 5556
rect 153988 5516 153994 5528
rect 154758 5516 154764 5528
rect 154816 5516 154822 5568
rect 155126 5516 155132 5568
rect 155184 5556 155190 5568
rect 155954 5556 155960 5568
rect 155184 5528 155960 5556
rect 155184 5516 155190 5528
rect 155954 5516 155960 5528
rect 156012 5516 156018 5568
rect 181990 5516 181996 5568
rect 182048 5556 182054 5568
rect 182542 5556 182548 5568
rect 182048 5528 182548 5556
rect 182048 5516 182054 5528
rect 182542 5516 182548 5528
rect 182600 5516 182606 5568
rect 183094 5516 183100 5568
rect 183152 5556 183158 5568
rect 183738 5556 183744 5568
rect 183152 5528 183744 5556
rect 183152 5516 183158 5528
rect 183738 5516 183744 5528
rect 183796 5516 183802 5568
rect 188798 5516 188804 5568
rect 188856 5556 188862 5568
rect 189626 5556 189632 5568
rect 188856 5528 189632 5556
rect 188856 5516 188862 5528
rect 189626 5516 189632 5528
rect 189684 5516 189690 5568
rect 189902 5516 189908 5568
rect 189960 5556 189966 5568
rect 190822 5556 190828 5568
rect 189960 5528 190828 5556
rect 189960 5516 189966 5528
rect 190822 5516 190828 5528
rect 190880 5516 190886 5568
rect 191098 5516 191104 5568
rect 191156 5556 191162 5568
rect 192018 5556 192024 5568
rect 191156 5528 192024 5556
rect 191156 5516 191162 5528
rect 192018 5516 192024 5528
rect 192076 5516 192082 5568
rect 192202 5516 192208 5568
rect 192260 5556 192266 5568
rect 193214 5556 193220 5568
rect 192260 5528 193220 5556
rect 192260 5516 192266 5528
rect 193214 5516 193220 5528
rect 193272 5516 193278 5568
rect 194502 5516 194508 5568
rect 194560 5556 194566 5568
rect 195606 5556 195612 5568
rect 194560 5528 195612 5556
rect 194560 5516 194566 5528
rect 195606 5516 195612 5528
rect 195664 5516 195670 5568
rect 196710 5516 196716 5568
rect 196768 5556 196774 5568
rect 197998 5556 198004 5568
rect 196768 5528 198004 5556
rect 196768 5516 196774 5528
rect 197998 5516 198004 5528
rect 198056 5516 198062 5568
rect 200114 5516 200120 5568
rect 200172 5556 200178 5568
rect 201494 5556 201500 5568
rect 200172 5528 201500 5556
rect 200172 5516 200178 5528
rect 201494 5516 201500 5528
rect 201552 5516 201558 5568
rect 202414 5516 202420 5568
rect 202472 5556 202478 5568
rect 203886 5556 203892 5568
rect 202472 5528 203892 5556
rect 202472 5516 202478 5528
rect 203886 5516 203892 5528
rect 203944 5516 203950 5568
rect 204622 5516 204628 5568
rect 204680 5556 204686 5568
rect 206278 5556 206284 5568
rect 204680 5528 206284 5556
rect 204680 5516 204686 5528
rect 206278 5516 206284 5528
rect 206336 5516 206342 5568
rect 208026 5516 208032 5568
rect 208084 5556 208090 5568
rect 209866 5556 209872 5568
rect 208084 5528 209872 5556
rect 208084 5516 208090 5528
rect 209866 5516 209872 5528
rect 209924 5516 209930 5568
rect 210326 5516 210332 5568
rect 210384 5556 210390 5568
rect 212258 5556 212264 5568
rect 210384 5528 212264 5556
rect 210384 5516 210390 5528
rect 212258 5516 212264 5528
rect 212316 5516 212322 5568
rect 212626 5516 212632 5568
rect 212684 5556 212690 5568
rect 214650 5556 214656 5568
rect 212684 5528 214656 5556
rect 212684 5516 212690 5528
rect 214650 5516 214656 5528
rect 214708 5516 214714 5568
rect 216030 5516 216036 5568
rect 216088 5556 216094 5568
rect 218146 5556 218152 5568
rect 216088 5528 218152 5556
rect 216088 5516 216094 5528
rect 218146 5516 218152 5528
rect 218204 5516 218210 5568
rect 218238 5516 218244 5568
rect 218296 5556 218302 5568
rect 220538 5556 220544 5568
rect 218296 5528 220544 5556
rect 218296 5516 218302 5528
rect 220538 5516 220544 5528
rect 220596 5516 220602 5568
rect 221642 5516 221648 5568
rect 221700 5556 221706 5568
rect 224126 5556 224132 5568
rect 221700 5528 224132 5556
rect 221700 5516 221706 5528
rect 224126 5516 224132 5528
rect 224184 5516 224190 5568
rect 225046 5516 225052 5568
rect 225104 5556 225110 5568
rect 227714 5556 227720 5568
rect 225104 5528 227720 5556
rect 225104 5516 225110 5528
rect 227714 5516 227720 5528
rect 227772 5516 227778 5568
rect 229646 5516 229652 5568
rect 229704 5556 229710 5568
rect 232498 5556 232504 5568
rect 229704 5528 232504 5556
rect 229704 5516 229710 5528
rect 232498 5516 232504 5528
rect 232556 5516 232562 5568
rect 233050 5516 233056 5568
rect 233108 5556 233114 5568
rect 235902 5556 235908 5568
rect 233108 5528 235908 5556
rect 233108 5516 233114 5528
rect 235902 5516 235908 5528
rect 235960 5516 235966 5568
rect 237558 5516 237564 5568
rect 237616 5556 237622 5568
rect 240778 5556 240784 5568
rect 237616 5528 240784 5556
rect 237616 5516 237622 5528
rect 240778 5516 240784 5528
rect 240836 5516 240842 5568
rect 240962 5516 240968 5568
rect 241020 5556 241026 5568
rect 244182 5556 244188 5568
rect 241020 5528 244188 5556
rect 241020 5516 241026 5528
rect 244182 5516 244188 5528
rect 244240 5516 244246 5568
rect 246574 5516 246580 5568
rect 246632 5556 246638 5568
rect 249242 5556 249248 5568
rect 246632 5528 249248 5556
rect 246632 5516 246638 5528
rect 249242 5516 249248 5528
rect 249300 5516 249306 5568
rect 251174 5516 251180 5568
rect 251232 5556 251238 5568
rect 255038 5556 255044 5568
rect 251232 5528 255044 5556
rect 251232 5516 251238 5528
rect 255038 5516 255044 5528
rect 255096 5516 255102 5568
rect 255682 5516 255688 5568
rect 255740 5556 255746 5568
rect 258994 5556 259000 5568
rect 255740 5528 259000 5556
rect 255740 5516 255746 5528
rect 258994 5516 259000 5528
rect 259052 5516 259058 5568
rect 259086 5516 259092 5568
rect 259144 5556 259150 5568
rect 261202 5556 261208 5568
rect 259144 5528 261208 5556
rect 259144 5516 259150 5528
rect 261202 5516 261208 5528
rect 261260 5516 261266 5568
rect 263594 5516 263600 5568
rect 263652 5556 263658 5568
rect 266446 5556 266452 5568
rect 263652 5528 266452 5556
rect 263652 5516 263658 5528
rect 266446 5516 266452 5528
rect 266504 5516 266510 5568
rect 268194 5516 268200 5568
rect 268252 5556 268258 5568
rect 270494 5556 270500 5568
rect 268252 5528 270500 5556
rect 268252 5516 268258 5528
rect 270494 5516 270500 5528
rect 270552 5516 270558 5568
rect 271598 5516 271604 5568
rect 271656 5556 271662 5568
rect 273990 5556 273996 5568
rect 271656 5528 273996 5556
rect 271656 5516 271662 5528
rect 273990 5516 273996 5528
rect 274048 5516 274054 5568
rect 274910 5516 274916 5568
rect 274968 5556 274974 5568
rect 278406 5556 278412 5568
rect 274968 5528 278412 5556
rect 274968 5516 274974 5528
rect 278406 5516 278412 5528
rect 278464 5516 278470 5568
rect 279510 5516 279516 5568
rect 279568 5556 279574 5568
rect 282086 5556 282092 5568
rect 279568 5528 282092 5556
rect 279568 5516 279574 5528
rect 282086 5516 282092 5528
rect 282144 5516 282150 5568
rect 285122 5516 285128 5568
rect 285180 5556 285186 5568
rect 288250 5556 288256 5568
rect 285180 5528 288256 5556
rect 285180 5516 285186 5528
rect 288250 5516 288256 5528
rect 288308 5516 288314 5568
rect 288526 5516 288532 5568
rect 288584 5556 288590 5568
rect 291378 5556 291384 5568
rect 288584 5528 291384 5556
rect 288584 5516 288590 5528
rect 291378 5516 291384 5528
rect 291436 5516 291442 5568
rect 294230 5516 294236 5568
rect 294288 5556 294294 5568
rect 297818 5556 297824 5568
rect 294288 5528 297824 5556
rect 294288 5516 294294 5528
rect 297818 5516 297824 5528
rect 297876 5516 297882 5568
rect 298738 5516 298744 5568
rect 298796 5556 298802 5568
rect 301774 5556 301780 5568
rect 298796 5528 301780 5556
rect 298796 5516 298802 5528
rect 301774 5516 301780 5528
rect 301832 5516 301838 5568
rect 306742 5516 306748 5568
rect 306800 5556 306806 5568
rect 309962 5556 309968 5568
rect 306800 5528 309968 5556
rect 306800 5516 306806 5528
rect 309962 5516 309968 5528
rect 310020 5516 310026 5568
rect 311250 5516 311256 5568
rect 311308 5556 311314 5568
rect 313366 5556 313372 5568
rect 311308 5528 313372 5556
rect 311308 5516 311314 5528
rect 313366 5516 313372 5528
rect 313424 5516 313430 5568
rect 313458 5516 313464 5568
rect 313516 5556 313522 5568
rect 317230 5556 317236 5568
rect 313516 5528 317236 5556
rect 313516 5516 313522 5528
rect 317230 5516 317236 5528
rect 317288 5516 317294 5568
rect 320266 5516 320272 5568
rect 320324 5556 320330 5568
rect 323026 5556 323032 5568
rect 320324 5528 323032 5556
rect 320324 5516 320330 5528
rect 323026 5516 323032 5528
rect 323084 5516 323090 5568
rect 325970 5516 325976 5568
rect 326028 5556 326034 5568
rect 329742 5556 329748 5568
rect 326028 5528 329748 5556
rect 326028 5516 326034 5528
rect 329742 5516 329748 5528
rect 329800 5516 329806 5568
rect 336182 5516 336188 5568
rect 336240 5556 336246 5568
rect 339402 5556 339408 5568
rect 336240 5528 339408 5556
rect 336240 5516 336246 5528
rect 339402 5516 339408 5528
rect 339460 5516 339466 5568
rect 339586 5516 339592 5568
rect 339644 5556 339650 5568
rect 342254 5556 342260 5568
rect 339644 5528 342260 5556
rect 339644 5516 339650 5528
rect 342254 5516 342260 5528
rect 342312 5516 342318 5568
rect 346394 5516 346400 5568
rect 346452 5556 346458 5568
rect 350350 5556 350356 5568
rect 346452 5528 350356 5556
rect 346452 5516 346458 5528
rect 350350 5516 350356 5528
rect 350408 5516 350414 5568
rect 352006 5516 352012 5568
rect 352064 5556 352070 5568
rect 355502 5556 355508 5568
rect 352064 5528 355508 5556
rect 352064 5516 352070 5528
rect 355502 5516 355508 5528
rect 355560 5516 355566 5568
rect 358814 5516 358820 5568
rect 358872 5556 358878 5568
rect 361574 5556 361580 5568
rect 358872 5528 361580 5556
rect 358872 5516 358878 5528
rect 361574 5516 361580 5528
rect 361632 5516 361638 5568
rect 366818 5516 366824 5568
rect 366876 5556 366882 5568
rect 368474 5556 368480 5568
rect 366876 5528 368480 5556
rect 366876 5516 366882 5528
rect 368474 5516 368480 5528
rect 368532 5516 368538 5568
rect 395154 5516 395160 5568
rect 395212 5556 395218 5568
rect 398650 5556 398656 5568
rect 395212 5528 398656 5556
rect 395212 5516 395218 5528
rect 398650 5516 398656 5528
rect 398708 5516 398714 5568
rect 425698 5516 425704 5568
rect 425756 5556 425762 5568
rect 428826 5556 428832 5568
rect 425756 5528 428832 5556
rect 425756 5516 425762 5528
rect 428826 5516 428832 5528
rect 428884 5516 428890 5568
rect 456334 5516 456340 5568
rect 456392 5556 456398 5568
rect 458634 5556 458640 5568
rect 456392 5528 458640 5556
rect 456392 5516 456398 5528
rect 458634 5516 458640 5528
rect 458692 5516 458698 5568
rect 471054 5516 471060 5568
rect 471112 5556 471118 5568
rect 474642 5556 474648 5568
rect 471112 5528 474648 5556
rect 471112 5516 471118 5528
rect 474642 5516 474648 5528
rect 474700 5516 474706 5568
rect 1104 5466 582820 5488
rect 1104 5414 36822 5466
rect 36874 5414 36886 5466
rect 36938 5414 36950 5466
rect 37002 5414 37014 5466
rect 37066 5414 37078 5466
rect 37130 5414 37142 5466
rect 37194 5414 37206 5466
rect 37258 5414 37270 5466
rect 37322 5414 37334 5466
rect 37386 5414 72822 5466
rect 72874 5414 72886 5466
rect 72938 5414 72950 5466
rect 73002 5414 73014 5466
rect 73066 5414 73078 5466
rect 73130 5414 73142 5466
rect 73194 5414 73206 5466
rect 73258 5414 73270 5466
rect 73322 5414 73334 5466
rect 73386 5414 108822 5466
rect 108874 5414 108886 5466
rect 108938 5414 108950 5466
rect 109002 5414 109014 5466
rect 109066 5414 109078 5466
rect 109130 5414 109142 5466
rect 109194 5414 109206 5466
rect 109258 5414 109270 5466
rect 109322 5414 109334 5466
rect 109386 5414 144822 5466
rect 144874 5414 144886 5466
rect 144938 5414 144950 5466
rect 145002 5414 145014 5466
rect 145066 5414 145078 5466
rect 145130 5414 145142 5466
rect 145194 5414 145206 5466
rect 145258 5414 145270 5466
rect 145322 5414 145334 5466
rect 145386 5414 180822 5466
rect 180874 5414 180886 5466
rect 180938 5414 180950 5466
rect 181002 5414 181014 5466
rect 181066 5414 181078 5466
rect 181130 5414 181142 5466
rect 181194 5414 181206 5466
rect 181258 5414 181270 5466
rect 181322 5414 181334 5466
rect 181386 5414 216822 5466
rect 216874 5414 216886 5466
rect 216938 5414 216950 5466
rect 217002 5414 217014 5466
rect 217066 5414 217078 5466
rect 217130 5414 217142 5466
rect 217194 5414 217206 5466
rect 217258 5414 217270 5466
rect 217322 5414 217334 5466
rect 217386 5414 252822 5466
rect 252874 5414 252886 5466
rect 252938 5414 252950 5466
rect 253002 5414 253014 5466
rect 253066 5414 253078 5466
rect 253130 5414 253142 5466
rect 253194 5414 253206 5466
rect 253258 5414 253270 5466
rect 253322 5414 253334 5466
rect 253386 5414 288822 5466
rect 288874 5414 288886 5466
rect 288938 5414 288950 5466
rect 289002 5414 289014 5466
rect 289066 5414 289078 5466
rect 289130 5414 289142 5466
rect 289194 5414 289206 5466
rect 289258 5414 289270 5466
rect 289322 5414 289334 5466
rect 289386 5414 324822 5466
rect 324874 5414 324886 5466
rect 324938 5414 324950 5466
rect 325002 5414 325014 5466
rect 325066 5414 325078 5466
rect 325130 5414 325142 5466
rect 325194 5414 325206 5466
rect 325258 5414 325270 5466
rect 325322 5414 325334 5466
rect 325386 5414 360822 5466
rect 360874 5414 360886 5466
rect 360938 5414 360950 5466
rect 361002 5414 361014 5466
rect 361066 5414 361078 5466
rect 361130 5414 361142 5466
rect 361194 5414 361206 5466
rect 361258 5414 361270 5466
rect 361322 5414 361334 5466
rect 361386 5414 396822 5466
rect 396874 5414 396886 5466
rect 396938 5414 396950 5466
rect 397002 5414 397014 5466
rect 397066 5414 397078 5466
rect 397130 5414 397142 5466
rect 397194 5414 397206 5466
rect 397258 5414 397270 5466
rect 397322 5414 397334 5466
rect 397386 5414 432822 5466
rect 432874 5414 432886 5466
rect 432938 5414 432950 5466
rect 433002 5414 433014 5466
rect 433066 5414 433078 5466
rect 433130 5414 433142 5466
rect 433194 5414 433206 5466
rect 433258 5414 433270 5466
rect 433322 5414 433334 5466
rect 433386 5414 468822 5466
rect 468874 5414 468886 5466
rect 468938 5414 468950 5466
rect 469002 5414 469014 5466
rect 469066 5414 469078 5466
rect 469130 5414 469142 5466
rect 469194 5414 469206 5466
rect 469258 5414 469270 5466
rect 469322 5414 469334 5466
rect 469386 5414 504822 5466
rect 504874 5414 504886 5466
rect 504938 5414 504950 5466
rect 505002 5414 505014 5466
rect 505066 5414 505078 5466
rect 505130 5414 505142 5466
rect 505194 5414 505206 5466
rect 505258 5414 505270 5466
rect 505322 5414 505334 5466
rect 505386 5414 540822 5466
rect 540874 5414 540886 5466
rect 540938 5414 540950 5466
rect 541002 5414 541014 5466
rect 541066 5414 541078 5466
rect 541130 5414 541142 5466
rect 541194 5414 541206 5466
rect 541258 5414 541270 5466
rect 541322 5414 541334 5466
rect 541386 5414 576822 5466
rect 576874 5414 576886 5466
rect 576938 5414 576950 5466
rect 577002 5414 577014 5466
rect 577066 5414 577078 5466
rect 577130 5414 577142 5466
rect 577194 5414 577206 5466
rect 577258 5414 577270 5466
rect 577322 5414 577334 5466
rect 577386 5414 582820 5466
rect 1104 5392 582820 5414
rect 1104 4922 582820 4944
rect 1104 4870 18822 4922
rect 18874 4870 18886 4922
rect 18938 4870 18950 4922
rect 19002 4870 19014 4922
rect 19066 4870 19078 4922
rect 19130 4870 19142 4922
rect 19194 4870 19206 4922
rect 19258 4870 19270 4922
rect 19322 4870 19334 4922
rect 19386 4870 54822 4922
rect 54874 4870 54886 4922
rect 54938 4870 54950 4922
rect 55002 4870 55014 4922
rect 55066 4870 55078 4922
rect 55130 4870 55142 4922
rect 55194 4870 55206 4922
rect 55258 4870 55270 4922
rect 55322 4870 55334 4922
rect 55386 4870 90822 4922
rect 90874 4870 90886 4922
rect 90938 4870 90950 4922
rect 91002 4870 91014 4922
rect 91066 4870 91078 4922
rect 91130 4870 91142 4922
rect 91194 4870 91206 4922
rect 91258 4870 91270 4922
rect 91322 4870 91334 4922
rect 91386 4870 126822 4922
rect 126874 4870 126886 4922
rect 126938 4870 126950 4922
rect 127002 4870 127014 4922
rect 127066 4870 127078 4922
rect 127130 4870 127142 4922
rect 127194 4870 127206 4922
rect 127258 4870 127270 4922
rect 127322 4870 127334 4922
rect 127386 4870 162822 4922
rect 162874 4870 162886 4922
rect 162938 4870 162950 4922
rect 163002 4870 163014 4922
rect 163066 4870 163078 4922
rect 163130 4870 163142 4922
rect 163194 4870 163206 4922
rect 163258 4870 163270 4922
rect 163322 4870 163334 4922
rect 163386 4870 198822 4922
rect 198874 4870 198886 4922
rect 198938 4870 198950 4922
rect 199002 4870 199014 4922
rect 199066 4870 199078 4922
rect 199130 4870 199142 4922
rect 199194 4870 199206 4922
rect 199258 4870 199270 4922
rect 199322 4870 199334 4922
rect 199386 4870 234822 4922
rect 234874 4870 234886 4922
rect 234938 4870 234950 4922
rect 235002 4870 235014 4922
rect 235066 4870 235078 4922
rect 235130 4870 235142 4922
rect 235194 4870 235206 4922
rect 235258 4870 235270 4922
rect 235322 4870 235334 4922
rect 235386 4870 270822 4922
rect 270874 4870 270886 4922
rect 270938 4870 270950 4922
rect 271002 4870 271014 4922
rect 271066 4870 271078 4922
rect 271130 4870 271142 4922
rect 271194 4870 271206 4922
rect 271258 4870 271270 4922
rect 271322 4870 271334 4922
rect 271386 4870 306822 4922
rect 306874 4870 306886 4922
rect 306938 4870 306950 4922
rect 307002 4870 307014 4922
rect 307066 4870 307078 4922
rect 307130 4870 307142 4922
rect 307194 4870 307206 4922
rect 307258 4870 307270 4922
rect 307322 4870 307334 4922
rect 307386 4870 342822 4922
rect 342874 4870 342886 4922
rect 342938 4870 342950 4922
rect 343002 4870 343014 4922
rect 343066 4870 343078 4922
rect 343130 4870 343142 4922
rect 343194 4870 343206 4922
rect 343258 4870 343270 4922
rect 343322 4870 343334 4922
rect 343386 4870 378822 4922
rect 378874 4870 378886 4922
rect 378938 4870 378950 4922
rect 379002 4870 379014 4922
rect 379066 4870 379078 4922
rect 379130 4870 379142 4922
rect 379194 4870 379206 4922
rect 379258 4870 379270 4922
rect 379322 4870 379334 4922
rect 379386 4870 414822 4922
rect 414874 4870 414886 4922
rect 414938 4870 414950 4922
rect 415002 4870 415014 4922
rect 415066 4870 415078 4922
rect 415130 4870 415142 4922
rect 415194 4870 415206 4922
rect 415258 4870 415270 4922
rect 415322 4870 415334 4922
rect 415386 4870 450822 4922
rect 450874 4870 450886 4922
rect 450938 4870 450950 4922
rect 451002 4870 451014 4922
rect 451066 4870 451078 4922
rect 451130 4870 451142 4922
rect 451194 4870 451206 4922
rect 451258 4870 451270 4922
rect 451322 4870 451334 4922
rect 451386 4870 486822 4922
rect 486874 4870 486886 4922
rect 486938 4870 486950 4922
rect 487002 4870 487014 4922
rect 487066 4870 487078 4922
rect 487130 4870 487142 4922
rect 487194 4870 487206 4922
rect 487258 4870 487270 4922
rect 487322 4870 487334 4922
rect 487386 4870 522822 4922
rect 522874 4870 522886 4922
rect 522938 4870 522950 4922
rect 523002 4870 523014 4922
rect 523066 4870 523078 4922
rect 523130 4870 523142 4922
rect 523194 4870 523206 4922
rect 523258 4870 523270 4922
rect 523322 4870 523334 4922
rect 523386 4870 558822 4922
rect 558874 4870 558886 4922
rect 558938 4870 558950 4922
rect 559002 4870 559014 4922
rect 559066 4870 559078 4922
rect 559130 4870 559142 4922
rect 559194 4870 559206 4922
rect 559258 4870 559270 4922
rect 559322 4870 559334 4922
rect 559386 4870 582820 4922
rect 1104 4848 582820 4870
rect 1104 4378 582820 4400
rect 1104 4326 36822 4378
rect 36874 4326 36886 4378
rect 36938 4326 36950 4378
rect 37002 4326 37014 4378
rect 37066 4326 37078 4378
rect 37130 4326 37142 4378
rect 37194 4326 37206 4378
rect 37258 4326 37270 4378
rect 37322 4326 37334 4378
rect 37386 4326 72822 4378
rect 72874 4326 72886 4378
rect 72938 4326 72950 4378
rect 73002 4326 73014 4378
rect 73066 4326 73078 4378
rect 73130 4326 73142 4378
rect 73194 4326 73206 4378
rect 73258 4326 73270 4378
rect 73322 4326 73334 4378
rect 73386 4326 108822 4378
rect 108874 4326 108886 4378
rect 108938 4326 108950 4378
rect 109002 4326 109014 4378
rect 109066 4326 109078 4378
rect 109130 4326 109142 4378
rect 109194 4326 109206 4378
rect 109258 4326 109270 4378
rect 109322 4326 109334 4378
rect 109386 4326 144822 4378
rect 144874 4326 144886 4378
rect 144938 4326 144950 4378
rect 145002 4326 145014 4378
rect 145066 4326 145078 4378
rect 145130 4326 145142 4378
rect 145194 4326 145206 4378
rect 145258 4326 145270 4378
rect 145322 4326 145334 4378
rect 145386 4326 180822 4378
rect 180874 4326 180886 4378
rect 180938 4326 180950 4378
rect 181002 4326 181014 4378
rect 181066 4326 181078 4378
rect 181130 4326 181142 4378
rect 181194 4326 181206 4378
rect 181258 4326 181270 4378
rect 181322 4326 181334 4378
rect 181386 4326 216822 4378
rect 216874 4326 216886 4378
rect 216938 4326 216950 4378
rect 217002 4326 217014 4378
rect 217066 4326 217078 4378
rect 217130 4326 217142 4378
rect 217194 4326 217206 4378
rect 217258 4326 217270 4378
rect 217322 4326 217334 4378
rect 217386 4326 252822 4378
rect 252874 4326 252886 4378
rect 252938 4326 252950 4378
rect 253002 4326 253014 4378
rect 253066 4326 253078 4378
rect 253130 4326 253142 4378
rect 253194 4326 253206 4378
rect 253258 4326 253270 4378
rect 253322 4326 253334 4378
rect 253386 4326 288822 4378
rect 288874 4326 288886 4378
rect 288938 4326 288950 4378
rect 289002 4326 289014 4378
rect 289066 4326 289078 4378
rect 289130 4326 289142 4378
rect 289194 4326 289206 4378
rect 289258 4326 289270 4378
rect 289322 4326 289334 4378
rect 289386 4326 324822 4378
rect 324874 4326 324886 4378
rect 324938 4326 324950 4378
rect 325002 4326 325014 4378
rect 325066 4326 325078 4378
rect 325130 4326 325142 4378
rect 325194 4326 325206 4378
rect 325258 4326 325270 4378
rect 325322 4326 325334 4378
rect 325386 4326 360822 4378
rect 360874 4326 360886 4378
rect 360938 4326 360950 4378
rect 361002 4326 361014 4378
rect 361066 4326 361078 4378
rect 361130 4326 361142 4378
rect 361194 4326 361206 4378
rect 361258 4326 361270 4378
rect 361322 4326 361334 4378
rect 361386 4326 396822 4378
rect 396874 4326 396886 4378
rect 396938 4326 396950 4378
rect 397002 4326 397014 4378
rect 397066 4326 397078 4378
rect 397130 4326 397142 4378
rect 397194 4326 397206 4378
rect 397258 4326 397270 4378
rect 397322 4326 397334 4378
rect 397386 4326 432822 4378
rect 432874 4326 432886 4378
rect 432938 4326 432950 4378
rect 433002 4326 433014 4378
rect 433066 4326 433078 4378
rect 433130 4326 433142 4378
rect 433194 4326 433206 4378
rect 433258 4326 433270 4378
rect 433322 4326 433334 4378
rect 433386 4326 468822 4378
rect 468874 4326 468886 4378
rect 468938 4326 468950 4378
rect 469002 4326 469014 4378
rect 469066 4326 469078 4378
rect 469130 4326 469142 4378
rect 469194 4326 469206 4378
rect 469258 4326 469270 4378
rect 469322 4326 469334 4378
rect 469386 4326 504822 4378
rect 504874 4326 504886 4378
rect 504938 4326 504950 4378
rect 505002 4326 505014 4378
rect 505066 4326 505078 4378
rect 505130 4326 505142 4378
rect 505194 4326 505206 4378
rect 505258 4326 505270 4378
rect 505322 4326 505334 4378
rect 505386 4326 540822 4378
rect 540874 4326 540886 4378
rect 540938 4326 540950 4378
rect 541002 4326 541014 4378
rect 541066 4326 541078 4378
rect 541130 4326 541142 4378
rect 541194 4326 541206 4378
rect 541258 4326 541270 4378
rect 541322 4326 541334 4378
rect 541386 4326 576822 4378
rect 576874 4326 576886 4378
rect 576938 4326 576950 4378
rect 577002 4326 577014 4378
rect 577066 4326 577078 4378
rect 577130 4326 577142 4378
rect 577194 4326 577206 4378
rect 577258 4326 577270 4378
rect 577322 4326 577334 4378
rect 577386 4326 582820 4378
rect 1104 4304 582820 4326
rect 547693 4199 547751 4205
rect 547693 4165 547705 4199
rect 547739 4196 547751 4199
rect 547969 4199 548027 4205
rect 547969 4196 547981 4199
rect 547739 4168 547981 4196
rect 547739 4165 547751 4168
rect 547693 4159 547751 4165
rect 547969 4165 547981 4168
rect 548015 4165 548027 4199
rect 563241 4199 563299 4205
rect 563241 4196 563253 4199
rect 547969 4159 548027 4165
rect 557184 4168 563253 4196
rect 20806 4088 20812 4140
rect 20864 4128 20870 4140
rect 27522 4128 27528 4140
rect 20864 4100 27528 4128
rect 20864 4088 20870 4100
rect 27522 4088 27528 4100
rect 27580 4088 27586 4140
rect 42150 4088 42156 4140
rect 42208 4128 42214 4140
rect 48222 4128 48228 4140
rect 42208 4100 48228 4128
rect 42208 4088 42214 4100
rect 48222 4088 48228 4100
rect 48280 4088 48286 4140
rect 61194 4088 61200 4140
rect 61252 4128 61258 4140
rect 66346 4128 66352 4140
rect 61252 4100 66352 4128
rect 61252 4088 61258 4100
rect 66346 4088 66352 4100
rect 66404 4088 66410 4140
rect 279786 4088 279792 4140
rect 279844 4128 279850 4140
rect 282454 4128 282460 4140
rect 279844 4100 282460 4128
rect 279844 4088 279850 4100
rect 282454 4088 282460 4100
rect 282512 4088 282518 4140
rect 285674 4088 285680 4140
rect 285732 4128 285738 4140
rect 289538 4128 289544 4140
rect 285732 4100 289544 4128
rect 285732 4088 285738 4100
rect 289538 4088 289544 4100
rect 289596 4088 289602 4140
rect 295426 4088 295432 4140
rect 295484 4128 295490 4140
rect 299106 4128 299112 4140
rect 295484 4100 299112 4128
rect 295484 4088 295490 4100
rect 299106 4088 299112 4100
rect 299164 4088 299170 4140
rect 303706 4088 303712 4140
rect 303764 4128 303770 4140
rect 307478 4128 307484 4140
rect 303764 4100 307484 4128
rect 303764 4088 303770 4100
rect 307478 4088 307484 4100
rect 307536 4088 307542 4140
rect 313366 4088 313372 4140
rect 313424 4128 313430 4140
rect 318058 4128 318064 4140
rect 313424 4100 318064 4128
rect 313424 4088 313430 4100
rect 318058 4088 318064 4100
rect 318116 4088 318122 4140
rect 322474 4088 322480 4140
rect 322532 4128 322538 4140
rect 326430 4128 326436 4140
rect 322532 4100 326436 4128
rect 322532 4088 322538 4100
rect 326430 4088 326436 4100
rect 326488 4088 326494 4140
rect 351730 4088 351736 4140
rect 351788 4128 351794 4140
rect 357342 4128 357348 4140
rect 351788 4100 357348 4128
rect 351788 4088 351794 4100
rect 357342 4088 357348 4100
rect 357400 4088 357406 4140
rect 408494 4088 408500 4140
rect 408552 4128 408558 4140
rect 410886 4128 410892 4140
rect 408552 4100 410892 4128
rect 408552 4088 408558 4100
rect 410886 4088 410892 4100
rect 410944 4088 410950 4140
rect 434530 4088 434536 4140
rect 434588 4128 434594 4140
rect 437014 4128 437020 4140
rect 434588 4100 437020 4128
rect 434588 4088 434594 4100
rect 437014 4088 437020 4100
rect 437072 4088 437078 4140
rect 448514 4088 448520 4140
rect 448572 4128 448578 4140
rect 452470 4128 452476 4140
rect 448572 4100 452476 4128
rect 448572 4088 448578 4100
rect 452470 4088 452476 4100
rect 452528 4088 452534 4140
rect 453666 4088 453672 4140
rect 453724 4128 453730 4140
rect 456058 4128 456064 4140
rect 453724 4100 456064 4128
rect 453724 4088 453730 4100
rect 456058 4088 456064 4100
rect 456116 4088 456122 4140
rect 459554 4088 459560 4140
rect 459612 4128 459618 4140
rect 463234 4128 463240 4140
rect 459612 4100 463240 4128
rect 459612 4088 459618 4100
rect 463234 4088 463240 4100
rect 463292 4088 463298 4140
rect 472526 4088 472532 4140
rect 472584 4128 472590 4140
rect 475102 4128 475108 4140
rect 472584 4100 475108 4128
rect 472584 4088 472590 4100
rect 475102 4088 475108 4100
rect 475160 4088 475166 4140
rect 477494 4088 477500 4140
rect 477552 4128 477558 4140
rect 481082 4128 481088 4140
rect 477552 4100 481088 4128
rect 477552 4088 477558 4100
rect 481082 4088 481088 4100
rect 481140 4088 481146 4140
rect 484394 4088 484400 4140
rect 484452 4128 484458 4140
rect 488166 4128 488172 4140
rect 484452 4100 488172 4128
rect 484452 4088 484458 4100
rect 488166 4088 488172 4100
rect 488224 4088 488230 4140
rect 535730 4088 535736 4140
rect 535788 4128 535794 4140
rect 553578 4128 553584 4140
rect 535788 4100 553584 4128
rect 535788 4088 535794 4100
rect 553578 4088 553584 4100
rect 553636 4088 553642 4140
rect 553854 4088 553860 4140
rect 553912 4128 553918 4140
rect 557184 4128 557212 4168
rect 563241 4165 563253 4168
rect 563287 4165 563299 4199
rect 563241 4159 563299 4165
rect 553912 4100 557212 4128
rect 553912 4088 553918 4100
rect 557258 4088 557264 4140
rect 557316 4128 557322 4140
rect 576210 4128 576216 4140
rect 557316 4100 576216 4128
rect 557316 4088 557322 4100
rect 576210 4088 576216 4100
rect 576268 4088 576274 4140
rect 566 4020 572 4072
rect 624 4060 630 4072
rect 8570 4060 8576 4072
rect 624 4032 8576 4060
rect 624 4020 630 4032
rect 8570 4020 8576 4032
rect 8628 4020 8634 4072
rect 11238 4020 11244 4072
rect 11296 4060 11302 4072
rect 16942 4060 16948 4072
rect 11296 4032 16948 4060
rect 11296 4020 11302 4032
rect 16942 4020 16948 4032
rect 17000 4020 17006 4072
rect 21910 4020 21916 4072
rect 21968 4060 21974 4072
rect 26234 4060 26240 4072
rect 21968 4032 26240 4060
rect 21968 4020 21974 4032
rect 26234 4020 26240 4032
rect 26292 4020 26298 4072
rect 31478 4020 31484 4072
rect 31536 4060 31542 4072
rect 36446 4060 36452 4072
rect 31536 4032 36452 4060
rect 31536 4020 31542 4032
rect 36446 4020 36452 4032
rect 36504 4020 36510 4072
rect 40954 4020 40960 4072
rect 41012 4060 41018 4072
rect 46842 4060 46848 4072
rect 41012 4032 46848 4060
rect 41012 4020 41018 4032
rect 46842 4020 46848 4032
rect 46900 4020 46906 4072
rect 50522 4020 50528 4072
rect 50580 4060 50586 4072
rect 56134 4060 56140 4072
rect 50580 4032 56140 4060
rect 50580 4020 50586 4032
rect 56134 4020 56140 4032
rect 56192 4020 56198 4072
rect 247034 4020 247040 4072
rect 247092 4060 247098 4072
rect 249150 4060 249156 4072
rect 247092 4032 249156 4060
rect 247092 4020 247098 4032
rect 249150 4020 249156 4032
rect 249208 4020 249214 4072
rect 256694 4020 256700 4072
rect 256752 4060 256758 4072
rect 258626 4060 258632 4072
rect 256752 4032 258632 4060
rect 256752 4020 256758 4032
rect 258626 4020 258632 4032
rect 258684 4020 258690 4072
rect 276014 4020 276020 4072
rect 276072 4060 276078 4072
rect 278866 4060 278872 4072
rect 276072 4032 278872 4060
rect 276072 4020 276078 4032
rect 278866 4020 278872 4032
rect 278924 4020 278930 4072
rect 285766 4020 285772 4072
rect 285824 4060 285830 4072
rect 288342 4060 288348 4072
rect 285824 4032 288348 4060
rect 285824 4020 285830 4032
rect 288342 4020 288348 4032
rect 288400 4020 288406 4072
rect 289446 4020 289452 4072
rect 289504 4060 289510 4072
rect 291930 4060 291936 4072
rect 289504 4032 291936 4060
rect 289504 4020 289510 4032
rect 291930 4020 291936 4032
rect 291988 4020 291994 4072
rect 294322 4020 294328 4072
rect 294380 4060 294386 4072
rect 297910 4060 297916 4072
rect 294380 4032 297916 4060
rect 294380 4020 294386 4032
rect 297910 4020 297916 4032
rect 297968 4020 297974 4072
rect 313090 4020 313096 4072
rect 313148 4060 313154 4072
rect 316954 4060 316960 4072
rect 313148 4032 316960 4060
rect 313148 4020 313154 4032
rect 316954 4020 316960 4032
rect 317012 4020 317018 4072
rect 332410 4020 332416 4072
rect 332468 4060 332474 4072
rect 337102 4060 337108 4072
rect 332468 4032 337108 4060
rect 332468 4020 332474 4032
rect 337102 4020 337108 4032
rect 337160 4020 337166 4072
rect 341794 4020 341800 4072
rect 341852 4060 341858 4072
rect 346670 4060 346676 4072
rect 341852 4032 346676 4060
rect 341852 4020 341858 4032
rect 346670 4020 346676 4032
rect 346728 4020 346734 4072
rect 360746 4020 360752 4072
rect 360804 4060 360810 4072
rect 366910 4060 366916 4072
rect 360804 4032 366916 4060
rect 360804 4020 360810 4032
rect 366910 4020 366916 4032
rect 366968 4020 366974 4072
rect 432690 4020 432696 4072
rect 432748 4060 432754 4072
rect 433518 4060 433524 4072
rect 432748 4032 433524 4060
rect 432748 4020 432754 4032
rect 433518 4020 433524 4032
rect 433576 4020 433582 4072
rect 445754 4020 445760 4072
rect 445812 4060 445818 4072
rect 448974 4060 448980 4072
rect 445812 4032 448980 4060
rect 445812 4020 445818 4032
rect 448974 4020 448980 4032
rect 449032 4020 449038 4072
rect 458174 4020 458180 4072
rect 458232 4060 458238 4072
rect 462038 4060 462044 4072
rect 458232 4032 462044 4060
rect 458232 4020 458238 4032
rect 462038 4020 462044 4032
rect 462096 4020 462102 4072
rect 467834 4020 467840 4072
rect 467892 4060 467898 4072
rect 471514 4060 471520 4072
rect 467892 4032 471520 4060
rect 467892 4020 467898 4032
rect 471514 4020 471520 4032
rect 471572 4020 471578 4072
rect 476114 4020 476120 4072
rect 476172 4060 476178 4072
rect 479886 4060 479892 4072
rect 476172 4032 479892 4060
rect 476172 4020 476178 4032
rect 479886 4020 479892 4032
rect 479944 4020 479950 4072
rect 490742 4020 490748 4072
rect 490800 4060 490806 4072
rect 495342 4060 495348 4072
rect 490800 4032 495348 4060
rect 490800 4020 490806 4032
rect 495342 4020 495348 4032
rect 495400 4020 495406 4072
rect 538493 4063 538551 4069
rect 538493 4060 538505 4063
rect 533356 4032 538505 4060
rect 25498 3952 25504 4004
rect 25556 3992 25562 4004
rect 31662 3992 31668 4004
rect 25556 3964 31668 3992
rect 25556 3952 25562 3964
rect 31662 3952 31668 3964
rect 31720 3952 31726 4004
rect 59998 3952 60004 4004
rect 60056 3992 60062 4004
rect 65242 3992 65248 4004
rect 60056 3964 65248 3992
rect 60056 3952 60062 3964
rect 65242 3952 65248 3964
rect 65300 3952 65306 4004
rect 266446 3952 266452 4004
rect 266504 3992 266510 4004
rect 268102 3992 268108 4004
rect 266504 3964 268108 3992
rect 266504 3952 266510 3964
rect 268102 3952 268108 3964
rect 268160 3952 268166 4004
rect 284386 3952 284392 4004
rect 284444 3992 284450 4004
rect 287146 3992 287152 4004
rect 284444 3964 287152 3992
rect 284444 3952 284450 3964
rect 287146 3952 287152 3964
rect 287204 3952 287210 4004
rect 304258 3952 304264 4004
rect 304316 3992 304322 4004
rect 308582 3992 308588 4004
rect 304316 3964 308588 3992
rect 304316 3952 304322 3964
rect 308582 3952 308588 3964
rect 308640 3952 308646 4004
rect 323026 3952 323032 4004
rect 323084 3992 323090 4004
rect 327626 3992 327632 4004
rect 323084 3964 327632 3992
rect 323084 3952 323090 3964
rect 327626 3952 327632 3964
rect 327684 3952 327690 4004
rect 336274 3952 336280 4004
rect 336332 3992 336338 4004
rect 340690 3992 340696 4004
rect 336332 3964 340696 3992
rect 336332 3952 336338 3964
rect 340690 3952 340696 3964
rect 340748 3952 340754 4004
rect 525794 3952 525800 4004
rect 525852 3992 525858 4004
rect 532234 3992 532240 4004
rect 525852 3964 532240 3992
rect 525852 3952 525858 3964
rect 532234 3952 532240 3964
rect 532292 3952 532298 4004
rect 6454 3884 6460 3936
rect 6512 3924 6518 3936
rect 11054 3924 11060 3936
rect 6512 3896 11060 3924
rect 6512 3884 6518 3896
rect 11054 3884 11060 3896
rect 11112 3884 11118 3936
rect 24302 3884 24308 3936
rect 24360 3924 24366 3936
rect 28994 3924 29000 3936
rect 24360 3896 29000 3924
rect 24360 3884 24366 3896
rect 28994 3884 29000 3896
rect 29052 3884 29058 3936
rect 43346 3884 43352 3936
rect 43404 3924 43410 3936
rect 49326 3924 49332 3936
rect 43404 3896 49332 3924
rect 43404 3884 43410 3896
rect 49326 3884 49332 3896
rect 49384 3884 49390 3936
rect 342714 3884 342720 3936
rect 342772 3924 342778 3936
rect 349062 3924 349068 3936
rect 342772 3896 349068 3924
rect 342772 3884 342778 3896
rect 349062 3884 349068 3896
rect 349120 3884 349126 3936
rect 525518 3884 525524 3936
rect 525576 3924 525582 3936
rect 533356 3924 533384 4032
rect 538493 4029 538505 4032
rect 538539 4029 538551 4063
rect 538493 4023 538551 4029
rect 541434 4020 541440 4072
rect 541492 4060 541498 4072
rect 545393 4063 545451 4069
rect 545393 4060 545405 4063
rect 541492 4032 545405 4060
rect 541492 4020 541498 4032
rect 545393 4029 545405 4032
rect 545439 4029 545451 4063
rect 545393 4023 545451 4029
rect 545942 4020 545948 4072
rect 546000 4060 546006 4072
rect 558181 4063 558239 4069
rect 558181 4060 558193 4063
rect 546000 4032 558193 4060
rect 546000 4020 546006 4032
rect 558181 4029 558193 4032
rect 558227 4029 558239 4063
rect 558181 4023 558239 4029
rect 558273 4063 558331 4069
rect 558273 4029 558285 4063
rect 558319 4060 558331 4063
rect 560570 4060 560576 4072
rect 558319 4032 560576 4060
rect 558319 4029 558331 4032
rect 558273 4023 558331 4029
rect 560570 4020 560576 4032
rect 560628 4020 560634 4072
rect 560662 4020 560668 4072
rect 560720 4060 560726 4072
rect 579798 4060 579804 4072
rect 560720 4032 579804 4060
rect 560720 4020 560726 4032
rect 579798 4020 579804 4032
rect 579856 4020 579862 4072
rect 533430 3952 533436 4004
rect 533488 3992 533494 4004
rect 551186 3992 551192 4004
rect 533488 3964 551192 3992
rect 533488 3952 533494 3964
rect 551186 3952 551192 3964
rect 551244 3952 551250 4004
rect 551554 3952 551560 4004
rect 551612 3992 551618 4004
rect 570230 3992 570236 4004
rect 551612 3964 570236 3992
rect 551612 3952 551618 3964
rect 570230 3952 570236 3964
rect 570288 3952 570294 4004
rect 525576 3896 533384 3924
rect 525576 3884 525582 3896
rect 535914 3884 535920 3936
rect 535972 3924 535978 3936
rect 538122 3924 538128 3936
rect 535972 3896 538128 3924
rect 535972 3884 535978 3896
rect 538122 3884 538128 3896
rect 538180 3884 538186 3936
rect 541618 3884 541624 3936
rect 541676 3924 541682 3936
rect 547693 3927 547751 3933
rect 547693 3924 547705 3927
rect 541676 3896 547705 3924
rect 541676 3884 541682 3896
rect 547693 3893 547705 3896
rect 547739 3893 547751 3927
rect 547693 3887 547751 3893
rect 547785 3927 547843 3933
rect 547785 3893 547797 3927
rect 547831 3924 547843 3927
rect 558273 3927 558331 3933
rect 558273 3924 558285 3927
rect 547831 3896 558285 3924
rect 547831 3893 547843 3896
rect 547785 3887 547843 3893
rect 558273 3893 558285 3896
rect 558319 3893 558331 3927
rect 558273 3887 558331 3893
rect 558362 3884 558368 3936
rect 558420 3924 558426 3936
rect 562045 3927 562103 3933
rect 562045 3924 562057 3927
rect 558420 3896 562057 3924
rect 558420 3884 558426 3896
rect 562045 3893 562057 3896
rect 562091 3893 562103 3927
rect 562045 3887 562103 3893
rect 562962 3884 562968 3936
rect 563020 3924 563026 3936
rect 582190 3924 582196 3936
rect 563020 3896 582196 3924
rect 563020 3884 563026 3896
rect 582190 3884 582196 3896
rect 582248 3884 582254 3936
rect 1104 3834 582820 3856
rect 1104 3782 18822 3834
rect 18874 3782 18886 3834
rect 18938 3782 18950 3834
rect 19002 3782 19014 3834
rect 19066 3782 19078 3834
rect 19130 3782 19142 3834
rect 19194 3782 19206 3834
rect 19258 3782 19270 3834
rect 19322 3782 19334 3834
rect 19386 3782 54822 3834
rect 54874 3782 54886 3834
rect 54938 3782 54950 3834
rect 55002 3782 55014 3834
rect 55066 3782 55078 3834
rect 55130 3782 55142 3834
rect 55194 3782 55206 3834
rect 55258 3782 55270 3834
rect 55322 3782 55334 3834
rect 55386 3782 90822 3834
rect 90874 3782 90886 3834
rect 90938 3782 90950 3834
rect 91002 3782 91014 3834
rect 91066 3782 91078 3834
rect 91130 3782 91142 3834
rect 91194 3782 91206 3834
rect 91258 3782 91270 3834
rect 91322 3782 91334 3834
rect 91386 3782 126822 3834
rect 126874 3782 126886 3834
rect 126938 3782 126950 3834
rect 127002 3782 127014 3834
rect 127066 3782 127078 3834
rect 127130 3782 127142 3834
rect 127194 3782 127206 3834
rect 127258 3782 127270 3834
rect 127322 3782 127334 3834
rect 127386 3782 162822 3834
rect 162874 3782 162886 3834
rect 162938 3782 162950 3834
rect 163002 3782 163014 3834
rect 163066 3782 163078 3834
rect 163130 3782 163142 3834
rect 163194 3782 163206 3834
rect 163258 3782 163270 3834
rect 163322 3782 163334 3834
rect 163386 3782 198822 3834
rect 198874 3782 198886 3834
rect 198938 3782 198950 3834
rect 199002 3782 199014 3834
rect 199066 3782 199078 3834
rect 199130 3782 199142 3834
rect 199194 3782 199206 3834
rect 199258 3782 199270 3834
rect 199322 3782 199334 3834
rect 199386 3782 234822 3834
rect 234874 3782 234886 3834
rect 234938 3782 234950 3834
rect 235002 3782 235014 3834
rect 235066 3782 235078 3834
rect 235130 3782 235142 3834
rect 235194 3782 235206 3834
rect 235258 3782 235270 3834
rect 235322 3782 235334 3834
rect 235386 3782 270822 3834
rect 270874 3782 270886 3834
rect 270938 3782 270950 3834
rect 271002 3782 271014 3834
rect 271066 3782 271078 3834
rect 271130 3782 271142 3834
rect 271194 3782 271206 3834
rect 271258 3782 271270 3834
rect 271322 3782 271334 3834
rect 271386 3782 306822 3834
rect 306874 3782 306886 3834
rect 306938 3782 306950 3834
rect 307002 3782 307014 3834
rect 307066 3782 307078 3834
rect 307130 3782 307142 3834
rect 307194 3782 307206 3834
rect 307258 3782 307270 3834
rect 307322 3782 307334 3834
rect 307386 3782 342822 3834
rect 342874 3782 342886 3834
rect 342938 3782 342950 3834
rect 343002 3782 343014 3834
rect 343066 3782 343078 3834
rect 343130 3782 343142 3834
rect 343194 3782 343206 3834
rect 343258 3782 343270 3834
rect 343322 3782 343334 3834
rect 343386 3782 378822 3834
rect 378874 3782 378886 3834
rect 378938 3782 378950 3834
rect 379002 3782 379014 3834
rect 379066 3782 379078 3834
rect 379130 3782 379142 3834
rect 379194 3782 379206 3834
rect 379258 3782 379270 3834
rect 379322 3782 379334 3834
rect 379386 3782 414822 3834
rect 414874 3782 414886 3834
rect 414938 3782 414950 3834
rect 415002 3782 415014 3834
rect 415066 3782 415078 3834
rect 415130 3782 415142 3834
rect 415194 3782 415206 3834
rect 415258 3782 415270 3834
rect 415322 3782 415334 3834
rect 415386 3782 450822 3834
rect 450874 3782 450886 3834
rect 450938 3782 450950 3834
rect 451002 3782 451014 3834
rect 451066 3782 451078 3834
rect 451130 3782 451142 3834
rect 451194 3782 451206 3834
rect 451258 3782 451270 3834
rect 451322 3782 451334 3834
rect 451386 3782 486822 3834
rect 486874 3782 486886 3834
rect 486938 3782 486950 3834
rect 487002 3782 487014 3834
rect 487066 3782 487078 3834
rect 487130 3782 487142 3834
rect 487194 3782 487206 3834
rect 487258 3782 487270 3834
rect 487322 3782 487334 3834
rect 487386 3782 522822 3834
rect 522874 3782 522886 3834
rect 522938 3782 522950 3834
rect 523002 3782 523014 3834
rect 523066 3782 523078 3834
rect 523130 3782 523142 3834
rect 523194 3782 523206 3834
rect 523258 3782 523270 3834
rect 523322 3782 523334 3834
rect 523386 3782 558822 3834
rect 558874 3782 558886 3834
rect 558938 3782 558950 3834
rect 559002 3782 559014 3834
rect 559066 3782 559078 3834
rect 559130 3782 559142 3834
rect 559194 3782 559206 3834
rect 559258 3782 559270 3834
rect 559322 3782 559334 3834
rect 559386 3782 582820 3834
rect 1104 3760 582820 3782
rect 266354 3680 266360 3732
rect 266412 3720 266418 3732
rect 269298 3720 269304 3732
rect 266412 3692 269304 3720
rect 266412 3680 266418 3692
rect 269298 3680 269304 3692
rect 269356 3680 269362 3732
rect 275094 3680 275100 3732
rect 275152 3720 275158 3732
rect 277670 3720 277676 3732
rect 275152 3692 277676 3720
rect 275152 3680 275158 3692
rect 277670 3680 277676 3692
rect 277728 3680 277734 3732
rect 292574 3680 292580 3732
rect 292632 3720 292638 3732
rect 296714 3720 296720 3732
rect 292632 3692 296720 3720
rect 292632 3680 292638 3692
rect 296714 3680 296720 3692
rect 296772 3680 296778 3732
rect 464430 3680 464436 3732
rect 464488 3720 464494 3732
rect 467926 3720 467932 3732
rect 464488 3692 467932 3720
rect 464488 3680 464494 3692
rect 467926 3680 467932 3692
rect 467984 3680 467990 3732
rect 469490 3680 469496 3732
rect 469548 3720 469554 3732
rect 472710 3720 472716 3732
rect 469548 3692 472716 3720
rect 469548 3680 469554 3692
rect 472710 3680 472716 3692
rect 472768 3680 472774 3732
rect 474090 3680 474096 3732
rect 474148 3720 474154 3732
rect 477494 3720 477500 3732
rect 474148 3692 477500 3720
rect 474148 3680 474154 3692
rect 477494 3680 477500 3692
rect 477552 3680 477558 3732
rect 510430 3680 510436 3732
rect 510488 3720 510494 3732
rect 515582 3720 515588 3732
rect 510488 3692 515588 3720
rect 510488 3680 510494 3692
rect 515582 3680 515588 3692
rect 515640 3680 515646 3732
rect 524506 3680 524512 3732
rect 524564 3720 524570 3732
rect 531038 3720 531044 3732
rect 524564 3692 531044 3720
rect 524564 3680 524570 3692
rect 531038 3680 531044 3692
rect 531096 3680 531102 3732
rect 531222 3680 531228 3732
rect 531280 3720 531286 3732
rect 548886 3720 548892 3732
rect 531280 3692 548892 3720
rect 531280 3680 531286 3692
rect 548886 3680 548892 3692
rect 548944 3680 548950 3732
rect 550450 3680 550456 3732
rect 550508 3720 550514 3732
rect 552661 3723 552719 3729
rect 552661 3720 552673 3723
rect 550508 3692 552673 3720
rect 550508 3680 550514 3692
rect 552661 3689 552673 3692
rect 552707 3689 552719 3723
rect 552661 3683 552719 3689
rect 552750 3680 552756 3732
rect 552808 3720 552814 3732
rect 571426 3720 571432 3732
rect 552808 3692 571432 3720
rect 552808 3680 552814 3692
rect 571426 3680 571432 3692
rect 571484 3680 571490 3732
rect 29086 3612 29092 3664
rect 29144 3652 29150 3664
rect 35710 3652 35716 3664
rect 29144 3624 35716 3652
rect 29144 3612 29150 3624
rect 35710 3612 35716 3624
rect 35768 3612 35774 3664
rect 45738 3612 45744 3664
rect 45796 3652 45802 3664
rect 51626 3652 51632 3664
rect 45796 3624 51632 3652
rect 45796 3612 45802 3624
rect 51626 3612 51632 3624
rect 51684 3612 51690 3664
rect 64782 3612 64788 3664
rect 64840 3652 64846 3664
rect 69750 3652 69756 3664
rect 64840 3624 69756 3652
rect 64840 3612 64846 3624
rect 69750 3612 69756 3624
rect 69808 3612 69814 3664
rect 332962 3612 332968 3664
rect 333020 3652 333026 3664
rect 338298 3652 338304 3664
rect 333020 3624 338304 3652
rect 333020 3612 333026 3624
rect 338298 3612 338304 3624
rect 338356 3612 338362 3664
rect 342254 3612 342260 3664
rect 342312 3652 342318 3664
rect 347866 3652 347872 3664
rect 342312 3624 347872 3652
rect 342312 3612 342318 3624
rect 347866 3612 347872 3624
rect 347924 3612 347930 3664
rect 413370 3612 413376 3664
rect 413428 3652 413434 3664
rect 421558 3652 421564 3664
rect 413428 3624 421564 3652
rect 413428 3612 413434 3624
rect 421558 3612 421564 3624
rect 421616 3612 421622 3664
rect 472894 3612 472900 3664
rect 472952 3652 472958 3664
rect 476298 3652 476304 3664
rect 472952 3624 476304 3652
rect 472952 3612 472958 3624
rect 476298 3612 476304 3624
rect 476356 3612 476362 3664
rect 478966 3612 478972 3664
rect 479024 3652 479030 3664
rect 483474 3652 483480 3664
rect 479024 3624 483480 3652
rect 479024 3612 479030 3624
rect 483474 3612 483480 3624
rect 483532 3612 483538 3664
rect 518710 3612 518716 3664
rect 518768 3652 518774 3664
rect 535730 3652 535736 3664
rect 518768 3624 535736 3652
rect 518768 3612 518774 3624
rect 535730 3612 535736 3624
rect 535788 3612 535794 3664
rect 538030 3612 538036 3664
rect 538088 3652 538094 3664
rect 547877 3655 547935 3661
rect 547877 3652 547889 3655
rect 538088 3624 547889 3652
rect 538088 3612 538094 3624
rect 547877 3621 547889 3624
rect 547923 3621 547935 3655
rect 547877 3615 547935 3621
rect 547969 3655 548027 3661
rect 547969 3621 547981 3655
rect 548015 3652 548027 3655
rect 559466 3652 559472 3664
rect 548015 3624 559472 3652
rect 548015 3621 548027 3624
rect 547969 3615 548027 3621
rect 559466 3612 559472 3624
rect 559524 3612 559530 3664
rect 559558 3612 559564 3664
rect 559616 3652 559622 3664
rect 578602 3652 578608 3664
rect 559616 3624 578608 3652
rect 559616 3612 559622 3624
rect 578602 3612 578608 3624
rect 578660 3612 578666 3664
rect 5258 3544 5264 3596
rect 5316 3584 5322 3596
rect 12250 3584 12256 3596
rect 5316 3556 12256 3584
rect 5316 3544 5322 3556
rect 12250 3544 12256 3556
rect 12308 3544 12314 3596
rect 16022 3544 16028 3596
rect 16080 3584 16086 3596
rect 20714 3584 20720 3596
rect 16080 3556 20720 3584
rect 16080 3544 16086 3556
rect 20714 3544 20720 3556
rect 20772 3544 20778 3596
rect 34974 3544 34980 3596
rect 35032 3584 35038 3596
rect 41322 3584 41328 3596
rect 35032 3556 41328 3584
rect 35032 3544 35038 3556
rect 41322 3544 41328 3556
rect 41380 3544 41386 3596
rect 44542 3544 44548 3596
rect 44600 3584 44606 3596
rect 50430 3584 50436 3596
rect 44600 3556 50436 3584
rect 44600 3544 44606 3556
rect 50430 3544 50436 3556
rect 50488 3544 50494 3596
rect 52822 3544 52828 3596
rect 52880 3584 52886 3596
rect 58434 3584 58440 3596
rect 52880 3556 58440 3584
rect 52880 3544 52886 3556
rect 58434 3544 58440 3556
rect 58492 3544 58498 3596
rect 74258 3544 74264 3596
rect 74316 3584 74322 3596
rect 78858 3584 78864 3596
rect 74316 3556 78864 3584
rect 74316 3544 74322 3556
rect 78858 3544 78864 3556
rect 78916 3544 78922 3596
rect 292482 3544 292488 3596
rect 292540 3584 292546 3596
rect 295518 3584 295524 3596
rect 292540 3556 295524 3584
rect 292540 3544 292546 3556
rect 295518 3544 295524 3556
rect 295576 3544 295582 3596
rect 304994 3544 305000 3596
rect 305052 3584 305058 3596
rect 309778 3584 309784 3596
rect 305052 3556 309784 3584
rect 305052 3544 305058 3556
rect 309778 3544 309784 3556
rect 309836 3544 309842 3596
rect 311802 3544 311808 3596
rect 311860 3584 311866 3596
rect 315758 3584 315764 3596
rect 311860 3556 315764 3584
rect 311860 3544 311866 3556
rect 315758 3544 315764 3556
rect 315816 3544 315822 3596
rect 324314 3544 324320 3596
rect 324372 3584 324378 3596
rect 330018 3584 330024 3596
rect 324372 3556 330024 3584
rect 324372 3544 324378 3556
rect 330018 3544 330024 3556
rect 330076 3544 330082 3596
rect 333974 3544 333980 3596
rect 334032 3584 334038 3596
rect 339494 3584 339500 3596
rect 334032 3556 339500 3584
rect 334032 3544 334038 3556
rect 339494 3544 339500 3556
rect 339552 3544 339558 3596
rect 352282 3544 352288 3596
rect 352340 3584 352346 3596
rect 358538 3584 358544 3596
rect 352340 3556 358544 3584
rect 352340 3544 352346 3556
rect 358538 3544 358544 3556
rect 358596 3544 358602 3596
rect 367462 3544 367468 3596
rect 367520 3584 367526 3596
rect 373994 3584 374000 3596
rect 367520 3556 374000 3584
rect 367520 3544 367526 3556
rect 373994 3544 374000 3556
rect 374052 3544 374058 3596
rect 433886 3544 433892 3596
rect 433944 3584 433950 3596
rect 435818 3584 435824 3596
rect 433944 3556 435824 3584
rect 433944 3544 433950 3556
rect 435818 3544 435824 3556
rect 435876 3544 435882 3596
rect 456794 3544 456800 3596
rect 456852 3584 456858 3596
rect 459646 3584 459652 3596
rect 456852 3556 459652 3584
rect 456852 3544 456858 3556
rect 459646 3544 459652 3556
rect 459704 3544 459710 3596
rect 463326 3544 463332 3596
rect 463384 3584 463390 3596
rect 465626 3584 465632 3596
rect 463384 3556 465632 3584
rect 463384 3544 463390 3556
rect 465626 3544 465632 3556
rect 465684 3544 465690 3596
rect 488534 3544 488540 3596
rect 488592 3584 488598 3596
rect 492950 3584 492956 3596
rect 488592 3556 492956 3584
rect 488592 3544 488598 3556
rect 492950 3544 492956 3556
rect 493008 3544 493014 3596
rect 496814 3544 496820 3596
rect 496872 3584 496878 3596
rect 501230 3584 501236 3596
rect 496872 3556 501236 3584
rect 496872 3544 496878 3556
rect 501230 3544 501236 3556
rect 501288 3544 501294 3596
rect 510522 3544 510528 3596
rect 510580 3584 510586 3596
rect 514386 3584 514392 3596
rect 510580 3556 514392 3584
rect 510580 3544 510586 3556
rect 514386 3544 514392 3556
rect 514444 3544 514450 3596
rect 519814 3544 519820 3596
rect 519872 3584 519878 3596
rect 536926 3584 536932 3596
rect 519872 3556 536932 3584
rect 519872 3544 519878 3556
rect 536926 3544 536932 3556
rect 536984 3544 536990 3596
rect 541805 3587 541863 3593
rect 541805 3584 541817 3587
rect 539060 3556 541817 3584
rect 7650 3476 7656 3528
rect 7708 3516 7714 3528
rect 15010 3516 15016 3528
rect 7708 3488 15016 3516
rect 7708 3476 7714 3488
rect 15010 3476 15016 3488
rect 15068 3476 15074 3528
rect 17218 3476 17224 3528
rect 17276 3516 17282 3528
rect 23106 3516 23112 3528
rect 17276 3488 23112 3516
rect 17276 3476 17282 3488
rect 23106 3476 23112 3488
rect 23164 3476 23170 3528
rect 26694 3476 26700 3528
rect 26752 3516 26758 3528
rect 31754 3516 31760 3528
rect 26752 3488 31760 3516
rect 26752 3476 26758 3488
rect 31754 3476 31760 3488
rect 31812 3476 31818 3528
rect 33870 3476 33876 3528
rect 33928 3516 33934 3528
rect 39942 3516 39948 3528
rect 33928 3488 39948 3516
rect 33928 3476 33934 3488
rect 39942 3476 39948 3488
rect 40000 3476 40006 3528
rect 51626 3476 51632 3528
rect 51684 3516 51690 3528
rect 57238 3516 57244 3528
rect 51684 3488 57244 3516
rect 51684 3476 51690 3488
rect 57238 3476 57244 3488
rect 57296 3476 57302 3528
rect 57606 3476 57612 3528
rect 57664 3516 57670 3528
rect 62942 3516 62948 3528
rect 57664 3488 62948 3516
rect 57664 3476 57670 3488
rect 62942 3476 62948 3488
rect 63000 3476 63006 3528
rect 65978 3476 65984 3528
rect 66036 3516 66042 3528
rect 70854 3516 70860 3528
rect 66036 3488 70860 3516
rect 66036 3476 66042 3488
rect 70854 3476 70860 3488
rect 70912 3476 70918 3528
rect 72694 3476 72700 3528
rect 72752 3516 72758 3528
rect 77662 3516 77668 3528
rect 72752 3488 77668 3516
rect 72752 3476 72758 3488
rect 77662 3476 77668 3488
rect 77720 3476 77726 3528
rect 149238 3476 149244 3528
rect 149296 3516 149302 3528
rect 150250 3516 150256 3528
rect 149296 3488 150256 3516
rect 149296 3476 149302 3488
rect 150250 3476 150256 3488
rect 150308 3476 150314 3528
rect 150434 3476 150440 3528
rect 150492 3516 150498 3528
rect 151354 3516 151360 3528
rect 150492 3488 151360 3516
rect 150492 3476 150498 3488
rect 151354 3476 151360 3488
rect 151412 3476 151418 3528
rect 156322 3476 156328 3528
rect 156380 3516 156386 3528
rect 157058 3516 157064 3528
rect 156380 3488 157064 3516
rect 156380 3476 156386 3488
rect 157058 3476 157064 3488
rect 157116 3476 157122 3528
rect 187694 3476 187700 3528
rect 187752 3516 187758 3528
rect 188430 3516 188436 3528
rect 187752 3488 188436 3516
rect 187752 3476 187758 3488
rect 188430 3476 188436 3488
rect 188488 3476 188494 3528
rect 193306 3476 193312 3528
rect 193364 3516 193370 3528
rect 194410 3516 194416 3528
rect 193364 3488 194416 3516
rect 193364 3476 193370 3488
rect 194410 3476 194416 3488
rect 194468 3476 194474 3528
rect 255406 3476 255412 3528
rect 255464 3516 255470 3528
rect 257430 3516 257436 3528
rect 255464 3488 257436 3516
rect 255464 3476 255470 3488
rect 257430 3476 257436 3488
rect 257488 3476 257494 3528
rect 262398 3476 262404 3528
rect 262456 3516 262462 3528
rect 264606 3516 264612 3528
rect 262456 3488 264612 3516
rect 262456 3476 262462 3488
rect 264606 3476 264612 3488
rect 264664 3476 264670 3528
rect 264974 3476 264980 3528
rect 265032 3516 265038 3528
rect 266998 3516 267004 3528
rect 265032 3488 267004 3516
rect 265032 3476 265038 3488
rect 266998 3476 267004 3488
rect 267056 3476 267062 3528
rect 282086 3476 282092 3528
rect 282144 3516 282150 3528
rect 284754 3516 284760 3528
rect 282144 3488 284760 3516
rect 282144 3476 282150 3488
rect 284754 3476 284760 3488
rect 284812 3476 284818 3528
rect 290182 3476 290188 3528
rect 290240 3516 290246 3528
rect 293126 3516 293132 3528
rect 290240 3488 293132 3516
rect 290240 3476 290246 3488
rect 293126 3476 293132 3488
rect 293184 3476 293190 3528
rect 300670 3476 300676 3528
rect 300728 3516 300734 3528
rect 303798 3516 303804 3528
rect 300728 3488 303804 3516
rect 300728 3476 300734 3488
rect 303798 3476 303804 3488
rect 303856 3476 303862 3528
rect 311158 3476 311164 3528
rect 311216 3516 311222 3528
rect 314562 3516 314568 3528
rect 311216 3488 314568 3516
rect 311216 3476 311222 3488
rect 314562 3476 314568 3488
rect 314620 3476 314626 3528
rect 323578 3476 323584 3528
rect 323636 3516 323642 3528
rect 328822 3516 328828 3528
rect 323636 3488 328828 3516
rect 323636 3476 323642 3488
rect 328822 3476 328828 3488
rect 328880 3476 328886 3528
rect 329742 3476 329748 3528
rect 329800 3516 329806 3528
rect 333606 3516 333612 3528
rect 329800 3488 333612 3516
rect 329800 3476 329806 3488
rect 333606 3476 333612 3488
rect 333664 3476 333670 3528
rect 339402 3476 339408 3528
rect 339460 3516 339466 3528
rect 344278 3516 344284 3528
rect 339460 3488 344284 3516
rect 339460 3476 339466 3488
rect 344278 3476 344284 3488
rect 344336 3476 344342 3528
rect 353294 3476 353300 3528
rect 353352 3516 353358 3528
rect 359734 3516 359740 3528
rect 353352 3488 359740 3516
rect 353352 3476 353358 3488
rect 359734 3476 359740 3488
rect 359792 3476 359798 3528
rect 474642 3476 474648 3528
rect 474700 3516 474706 3528
rect 474700 3488 478828 3516
rect 474700 3476 474706 3488
rect 4062 3408 4068 3460
rect 4120 3448 4126 3460
rect 11606 3448 11612 3460
rect 4120 3420 11612 3448
rect 4120 3408 4126 3420
rect 11606 3408 11612 3420
rect 11664 3408 11670 3460
rect 14826 3408 14832 3460
rect 14884 3448 14890 3460
rect 19426 3448 19432 3460
rect 14884 3420 19432 3448
rect 14884 3408 14890 3420
rect 19426 3408 19432 3420
rect 19484 3408 19490 3460
rect 27890 3408 27896 3460
rect 27948 3448 27954 3460
rect 34330 3448 34336 3460
rect 27948 3420 34336 3448
rect 27948 3408 27954 3420
rect 34330 3408 34336 3420
rect 34388 3408 34394 3460
rect 38562 3408 38568 3460
rect 38620 3448 38626 3460
rect 42794 3448 42800 3460
rect 38620 3420 42800 3448
rect 38620 3408 38626 3420
rect 42794 3408 42800 3420
rect 42852 3408 42858 3460
rect 48130 3408 48136 3460
rect 48188 3448 48194 3460
rect 53650 3448 53656 3460
rect 48188 3420 53656 3448
rect 48188 3408 48194 3420
rect 53650 3408 53656 3420
rect 53708 3408 53714 3460
rect 54018 3408 54024 3460
rect 54076 3448 54082 3460
rect 59538 3448 59544 3460
rect 54076 3420 59544 3448
rect 54076 3408 54082 3420
rect 59538 3408 59544 3420
rect 59596 3408 59602 3460
rect 68278 3408 68284 3460
rect 68336 3448 68342 3460
rect 73430 3448 73436 3460
rect 68336 3420 73436 3448
rect 68336 3408 68342 3420
rect 73430 3408 73436 3420
rect 73488 3408 73494 3460
rect 254210 3408 254216 3460
rect 254268 3448 254274 3460
rect 256234 3448 256240 3460
rect 254268 3420 256240 3448
rect 254268 3408 254274 3420
rect 256234 3408 256240 3420
rect 256292 3408 256298 3460
rect 261202 3408 261208 3460
rect 261260 3448 261266 3460
rect 263410 3448 263416 3460
rect 261260 3420 263416 3448
rect 261260 3408 261266 3420
rect 263410 3408 263416 3420
rect 263468 3408 263474 3460
rect 263686 3408 263692 3460
rect 263744 3448 263750 3460
rect 265802 3448 265808 3460
rect 263744 3420 265808 3448
rect 263744 3408 263750 3420
rect 265802 3408 265808 3420
rect 265860 3408 265866 3460
rect 270494 3408 270500 3460
rect 270552 3448 270558 3460
rect 272886 3448 272892 3460
rect 270552 3420 272892 3448
rect 270552 3408 270558 3420
rect 272886 3408 272892 3420
rect 272944 3408 272950 3460
rect 272978 3408 272984 3460
rect 273036 3448 273042 3460
rect 275278 3448 275284 3460
rect 273036 3420 275284 3448
rect 273036 3408 273042 3420
rect 275278 3408 275284 3420
rect 275336 3408 275342 3460
rect 299198 3408 299204 3460
rect 299256 3448 299262 3460
rect 302602 3448 302608 3460
rect 299256 3420 302608 3448
rect 299256 3408 299262 3420
rect 302602 3408 302608 3420
rect 302660 3408 302666 3460
rect 303062 3408 303068 3460
rect 303120 3448 303126 3460
rect 306190 3448 306196 3460
rect 303120 3420 306196 3448
rect 303120 3408 303126 3420
rect 306190 3408 306196 3420
rect 306248 3408 306254 3460
rect 309962 3408 309968 3460
rect 310020 3448 310026 3460
rect 313366 3448 313372 3460
rect 310020 3420 313372 3448
rect 310020 3408 310026 3420
rect 313366 3408 313372 3420
rect 313424 3408 313430 3460
rect 314654 3408 314660 3460
rect 314712 3448 314718 3460
rect 319254 3448 319260 3460
rect 314712 3420 319260 3448
rect 314712 3408 314718 3420
rect 319254 3408 319260 3420
rect 319312 3408 319318 3460
rect 320082 3408 320088 3460
rect 320140 3448 320146 3460
rect 324038 3448 324044 3460
rect 320140 3420 324044 3448
rect 320140 3408 320146 3420
rect 324038 3408 324044 3420
rect 324096 3408 324102 3460
rect 330846 3408 330852 3460
rect 330904 3448 330910 3460
rect 334710 3448 334716 3460
rect 330904 3420 334716 3448
rect 330904 3408 330910 3420
rect 334710 3408 334716 3420
rect 334768 3408 334774 3460
rect 343634 3408 343640 3460
rect 343692 3448 343698 3460
rect 350258 3448 350264 3460
rect 343692 3420 350264 3448
rect 343692 3408 343698 3420
rect 350258 3408 350264 3420
rect 350316 3408 350322 3460
rect 350350 3408 350356 3460
rect 350408 3448 350414 3460
rect 354950 3448 354956 3460
rect 350408 3420 354956 3448
rect 350408 3408 350414 3420
rect 354950 3408 354956 3420
rect 355008 3408 355014 3460
rect 361574 3408 361580 3460
rect 361632 3448 361638 3460
rect 368014 3448 368020 3460
rect 361632 3420 368020 3448
rect 361632 3408 361638 3420
rect 368014 3408 368020 3420
rect 368072 3408 368078 3460
rect 382274 3408 382280 3460
rect 382332 3448 382338 3460
rect 390646 3448 390652 3460
rect 382332 3420 390652 3448
rect 382332 3408 382338 3420
rect 390646 3408 390652 3420
rect 390704 3408 390710 3460
rect 398650 3408 398656 3460
rect 398708 3448 398714 3460
rect 406102 3448 406108 3460
rect 398708 3420 406108 3448
rect 398708 3408 398714 3420
rect 406102 3408 406108 3420
rect 406160 3408 406166 3460
rect 413922 3408 413928 3460
rect 413980 3448 413986 3460
rect 422754 3448 422760 3460
rect 413980 3420 422760 3448
rect 413980 3408 413986 3420
rect 422754 3408 422760 3420
rect 422812 3408 422818 3460
rect 426434 3408 426440 3460
rect 426492 3448 426498 3460
rect 428734 3448 428740 3460
rect 426492 3420 428740 3448
rect 426492 3408 426498 3420
rect 428734 3408 428740 3420
rect 428792 3408 428798 3460
rect 428826 3408 428832 3460
rect 428884 3448 428890 3460
rect 438210 3448 438216 3460
rect 428884 3420 438216 3448
rect 428884 3408 428890 3420
rect 438210 3408 438216 3420
rect 438268 3408 438274 3460
rect 444282 3408 444288 3460
rect 444340 3448 444346 3460
rect 453666 3448 453672 3460
rect 444340 3420 453672 3448
rect 444340 3408 444346 3420
rect 453666 3408 453672 3420
rect 453724 3408 453730 3460
rect 458634 3408 458640 3460
rect 458692 3448 458698 3460
rect 458692 3420 462176 3448
rect 458692 3408 458698 3420
rect 8846 3340 8852 3392
rect 8904 3380 8910 3392
rect 13814 3380 13820 3392
rect 8904 3352 13820 3380
rect 8904 3340 8910 3352
rect 13814 3340 13820 3352
rect 13872 3340 13878 3392
rect 18322 3340 18328 3392
rect 18380 3380 18386 3392
rect 23842 3380 23848 3392
rect 18380 3352 23848 3380
rect 18380 3340 18386 3352
rect 23842 3340 23848 3352
rect 23900 3340 23906 3392
rect 36170 3340 36176 3392
rect 36228 3380 36234 3392
rect 42518 3380 42524 3392
rect 36228 3352 42524 3380
rect 36228 3340 36234 3352
rect 42518 3340 42524 3352
rect 42576 3340 42582 3392
rect 58802 3340 58808 3392
rect 58860 3380 58866 3392
rect 64046 3380 64052 3392
rect 58860 3352 64052 3380
rect 58860 3340 58866 3352
rect 64046 3340 64052 3352
rect 64104 3340 64110 3392
rect 280890 3340 280896 3392
rect 280948 3380 280954 3392
rect 283650 3380 283656 3392
rect 280948 3352 283656 3380
rect 280948 3340 280954 3352
rect 283650 3340 283656 3352
rect 283708 3340 283714 3392
rect 291378 3340 291384 3392
rect 291436 3380 291442 3392
rect 294322 3380 294328 3392
rect 291436 3352 294328 3380
rect 291436 3340 291442 3352
rect 294322 3340 294328 3352
rect 294380 3340 294386 3392
rect 301774 3340 301780 3392
rect 301832 3380 301838 3392
rect 304994 3380 305000 3392
rect 301832 3352 305000 3380
rect 301832 3340 301838 3352
rect 304994 3340 305000 3352
rect 305052 3340 305058 3392
rect 321462 3340 321468 3392
rect 321520 3380 321526 3392
rect 325418 3380 325424 3392
rect 321520 3352 325424 3380
rect 321520 3340 321526 3352
rect 325418 3340 325424 3352
rect 325476 3340 325482 3392
rect 348970 3340 348976 3392
rect 349028 3380 349034 3392
rect 353754 3380 353760 3392
rect 349028 3352 353760 3380
rect 349028 3340 349034 3352
rect 353754 3340 353760 3352
rect 353812 3340 353818 3392
rect 368474 3340 368480 3392
rect 368532 3380 368538 3392
rect 376386 3380 376392 3392
rect 368532 3352 376392 3380
rect 368532 3340 368538 3352
rect 376386 3340 376392 3352
rect 376444 3340 376450 3392
rect 394050 3340 394056 3392
rect 394108 3380 394114 3392
rect 395430 3380 395436 3392
rect 394108 3352 395436 3380
rect 394108 3340 394114 3352
rect 395430 3340 395436 3352
rect 395488 3340 395494 3392
rect 429194 3340 429200 3392
rect 429252 3380 429258 3392
rect 431126 3380 431132 3392
rect 429252 3352 431132 3380
rect 429252 3340 429258 3352
rect 431126 3340 431132 3352
rect 431184 3340 431190 3392
rect 437474 3340 437480 3392
rect 437532 3380 437538 3392
rect 439406 3380 439412 3392
rect 437532 3352 439412 3380
rect 437532 3340 437538 3352
rect 439406 3340 439412 3352
rect 439464 3340 439470 3392
rect 442350 3340 442356 3392
rect 442408 3380 442414 3392
rect 444190 3380 444196 3392
rect 442408 3352 444196 3380
rect 442408 3340 442414 3352
rect 444190 3340 444196 3352
rect 444248 3340 444254 3392
rect 445846 3340 445852 3392
rect 445904 3380 445910 3392
rect 447778 3380 447784 3392
rect 445904 3352 447784 3380
rect 445904 3340 445910 3352
rect 447778 3340 447784 3352
rect 447836 3340 447842 3392
rect 453114 3340 453120 3392
rect 453172 3380 453178 3392
rect 454862 3380 454868 3392
rect 453172 3352 454868 3380
rect 453172 3340 453178 3352
rect 454862 3340 454868 3352
rect 454920 3340 454926 3392
rect 462148 3380 462176 3420
rect 462222 3408 462228 3460
rect 462280 3448 462286 3460
rect 464430 3448 464436 3460
rect 462280 3420 464436 3448
rect 462280 3408 462286 3420
rect 464430 3408 464436 3420
rect 464488 3408 464494 3460
rect 469398 3408 469404 3460
rect 469456 3448 469462 3460
rect 473906 3448 473912 3460
rect 469456 3420 473912 3448
rect 469456 3408 469462 3420
rect 473906 3408 473912 3420
rect 473964 3408 473970 3460
rect 474734 3408 474740 3460
rect 474792 3448 474798 3460
rect 478690 3448 478696 3460
rect 474792 3420 478696 3448
rect 474792 3408 474798 3420
rect 478690 3408 478696 3420
rect 478748 3408 478754 3460
rect 478800 3448 478828 3488
rect 478874 3476 478880 3528
rect 478932 3516 478938 3528
rect 484578 3516 484584 3528
rect 478932 3488 484584 3516
rect 478932 3476 478938 3488
rect 484578 3476 484584 3488
rect 484636 3476 484642 3528
rect 506474 3476 506480 3528
rect 506532 3516 506538 3528
rect 511994 3516 512000 3528
rect 506532 3488 512000 3516
rect 506532 3476 506538 3488
rect 511994 3476 512000 3488
rect 512052 3476 512058 3528
rect 527818 3476 527824 3528
rect 527876 3516 527882 3528
rect 538953 3519 539011 3525
rect 538953 3516 538965 3519
rect 527876 3488 538965 3516
rect 527876 3476 527882 3488
rect 538953 3485 538965 3488
rect 538999 3485 539011 3519
rect 538953 3479 539011 3485
rect 485774 3448 485780 3460
rect 478800 3420 485780 3448
rect 485774 3408 485780 3420
rect 485832 3408 485838 3460
rect 491202 3408 491208 3460
rect 491260 3448 491266 3460
rect 503622 3448 503628 3460
rect 491260 3420 503628 3448
rect 491260 3408 491266 3420
rect 503622 3408 503628 3420
rect 503680 3408 503686 3460
rect 511718 3408 511724 3460
rect 511776 3448 511782 3460
rect 528646 3448 528652 3460
rect 511776 3420 528652 3448
rect 511776 3408 511782 3420
rect 528646 3408 528652 3420
rect 528704 3408 528710 3460
rect 534626 3408 534632 3460
rect 534684 3448 534690 3460
rect 539060 3448 539088 3556
rect 541805 3553 541817 3556
rect 541851 3553 541863 3587
rect 541805 3547 541863 3553
rect 542538 3544 542544 3596
rect 542596 3584 542602 3596
rect 547693 3587 547751 3593
rect 547693 3584 547705 3587
rect 542596 3556 547705 3584
rect 542596 3544 542602 3556
rect 547693 3553 547705 3556
rect 547739 3553 547751 3587
rect 547693 3547 547751 3553
rect 547782 3544 547788 3596
rect 547840 3584 547846 3596
rect 563146 3584 563152 3596
rect 547840 3556 563152 3584
rect 547840 3544 547846 3556
rect 563146 3544 563152 3556
rect 563204 3544 563210 3596
rect 563241 3587 563299 3593
rect 563241 3553 563253 3587
rect 563287 3584 563299 3587
rect 564437 3587 564495 3593
rect 564437 3584 564449 3587
rect 563287 3556 564449 3584
rect 563287 3553 563299 3556
rect 563241 3547 563299 3553
rect 564437 3553 564449 3556
rect 564483 3553 564495 3587
rect 564437 3547 564495 3553
rect 564526 3544 564532 3596
rect 564584 3584 564590 3596
rect 567105 3587 567163 3593
rect 567105 3584 567117 3587
rect 564584 3556 567117 3584
rect 564584 3544 564590 3556
rect 567105 3553 567117 3556
rect 567151 3553 567163 3587
rect 567105 3547 567163 3553
rect 539229 3519 539287 3525
rect 539229 3485 539241 3519
rect 539275 3516 539287 3519
rect 545298 3516 545304 3528
rect 539275 3488 545304 3516
rect 539275 3485 539287 3488
rect 539229 3479 539287 3485
rect 545298 3476 545304 3488
rect 545356 3476 545362 3528
rect 545393 3519 545451 3525
rect 545393 3485 545405 3519
rect 545439 3516 545451 3519
rect 546586 3516 546592 3528
rect 545439 3488 546592 3516
rect 545439 3485 545451 3488
rect 545393 3479 545451 3485
rect 546586 3476 546592 3488
rect 546644 3476 546650 3528
rect 547046 3476 547052 3528
rect 547104 3516 547110 3528
rect 552661 3519 552719 3525
rect 552661 3516 552673 3519
rect 547104 3488 552673 3516
rect 547104 3476 547110 3488
rect 552661 3485 552673 3488
rect 552707 3485 552719 3519
rect 552661 3479 552719 3485
rect 552753 3519 552811 3525
rect 552753 3485 552765 3519
rect 552799 3516 552811 3519
rect 569034 3516 569040 3528
rect 552799 3488 569040 3516
rect 552799 3485 552811 3488
rect 552753 3479 552811 3485
rect 569034 3476 569040 3488
rect 569092 3476 569098 3528
rect 534684 3420 539088 3448
rect 534684 3408 534690 3420
rect 539134 3408 539140 3460
rect 539192 3448 539198 3460
rect 544197 3451 544255 3457
rect 544197 3448 544209 3451
rect 539192 3420 544209 3448
rect 539192 3408 539198 3420
rect 544197 3417 544209 3420
rect 544243 3417 544255 3451
rect 544197 3411 544255 3417
rect 544746 3408 544752 3460
rect 544804 3448 544810 3460
rect 547598 3448 547604 3460
rect 544804 3420 547604 3448
rect 544804 3408 544810 3420
rect 547598 3408 547604 3420
rect 547656 3408 547662 3460
rect 559653 3451 559711 3457
rect 559653 3448 559665 3451
rect 547708 3420 559665 3448
rect 470318 3380 470324 3392
rect 462148 3352 470324 3380
rect 470318 3340 470324 3352
rect 470376 3340 470382 3392
rect 477586 3340 477592 3392
rect 477644 3380 477650 3392
rect 482278 3380 482284 3392
rect 477644 3352 482284 3380
rect 477644 3340 477650 3352
rect 482278 3340 482284 3352
rect 482336 3340 482342 3392
rect 487430 3340 487436 3392
rect 487488 3380 487494 3392
rect 491754 3380 491760 3392
rect 487488 3352 491760 3380
rect 487488 3340 487494 3352
rect 491754 3340 491760 3352
rect 491812 3340 491818 3392
rect 503898 3340 503904 3392
rect 503956 3380 503962 3392
rect 509602 3380 509608 3392
rect 503956 3352 509608 3380
rect 503956 3340 503962 3352
rect 509602 3340 509608 3352
rect 509660 3340 509666 3392
rect 520826 3340 520832 3392
rect 520884 3380 520890 3392
rect 522666 3380 522672 3392
rect 520884 3352 522672 3380
rect 520884 3340 520890 3352
rect 522666 3340 522672 3352
rect 522724 3340 522730 3392
rect 538493 3383 538551 3389
rect 538493 3349 538505 3383
rect 538539 3380 538551 3383
rect 542906 3380 542912 3392
rect 538539 3352 542912 3380
rect 538539 3349 538551 3352
rect 538493 3343 538551 3349
rect 542906 3340 542912 3352
rect 542964 3340 542970 3392
rect 543642 3340 543648 3392
rect 543700 3380 543706 3392
rect 547708 3380 547736 3420
rect 559653 3417 559665 3420
rect 559699 3417 559711 3451
rect 561674 3448 561680 3460
rect 559653 3411 559711 3417
rect 559760 3420 561680 3448
rect 543700 3352 547736 3380
rect 543700 3340 543706 3352
rect 547782 3340 547788 3392
rect 547840 3380 547846 3392
rect 558362 3380 558368 3392
rect 547840 3352 558368 3380
rect 547840 3340 547846 3352
rect 558362 3340 558368 3352
rect 558420 3340 558426 3392
rect 558457 3383 558515 3389
rect 558457 3349 558469 3383
rect 558503 3380 558515 3383
rect 559760 3380 559788 3420
rect 561674 3408 561680 3420
rect 561732 3408 561738 3460
rect 561766 3408 561772 3460
rect 561824 3448 561830 3460
rect 580994 3448 581000 3460
rect 561824 3420 581000 3448
rect 561824 3408 561830 3420
rect 580994 3408 581000 3420
rect 581052 3408 581058 3460
rect 558503 3352 559788 3380
rect 559837 3383 559895 3389
rect 558503 3349 558515 3352
rect 558457 3343 558515 3349
rect 559837 3349 559849 3383
rect 559883 3380 559895 3383
rect 561950 3380 561956 3392
rect 559883 3352 561956 3380
rect 559883 3349 559895 3352
rect 559837 3343 559895 3349
rect 561950 3340 561956 3352
rect 562008 3340 562014 3392
rect 562045 3383 562103 3389
rect 562045 3349 562057 3383
rect 562091 3380 562103 3383
rect 577406 3380 577412 3392
rect 562091 3352 577412 3380
rect 562091 3349 562103 3352
rect 562045 3343 562103 3349
rect 577406 3340 577412 3352
rect 577464 3340 577470 3392
rect 1104 3290 582820 3312
rect 1104 3238 36822 3290
rect 36874 3238 36886 3290
rect 36938 3238 36950 3290
rect 37002 3238 37014 3290
rect 37066 3238 37078 3290
rect 37130 3238 37142 3290
rect 37194 3238 37206 3290
rect 37258 3238 37270 3290
rect 37322 3238 37334 3290
rect 37386 3238 72822 3290
rect 72874 3238 72886 3290
rect 72938 3238 72950 3290
rect 73002 3238 73014 3290
rect 73066 3238 73078 3290
rect 73130 3238 73142 3290
rect 73194 3238 73206 3290
rect 73258 3238 73270 3290
rect 73322 3238 73334 3290
rect 73386 3238 108822 3290
rect 108874 3238 108886 3290
rect 108938 3238 108950 3290
rect 109002 3238 109014 3290
rect 109066 3238 109078 3290
rect 109130 3238 109142 3290
rect 109194 3238 109206 3290
rect 109258 3238 109270 3290
rect 109322 3238 109334 3290
rect 109386 3238 144822 3290
rect 144874 3238 144886 3290
rect 144938 3238 144950 3290
rect 145002 3238 145014 3290
rect 145066 3238 145078 3290
rect 145130 3238 145142 3290
rect 145194 3238 145206 3290
rect 145258 3238 145270 3290
rect 145322 3238 145334 3290
rect 145386 3238 180822 3290
rect 180874 3238 180886 3290
rect 180938 3238 180950 3290
rect 181002 3238 181014 3290
rect 181066 3238 181078 3290
rect 181130 3238 181142 3290
rect 181194 3238 181206 3290
rect 181258 3238 181270 3290
rect 181322 3238 181334 3290
rect 181386 3238 216822 3290
rect 216874 3238 216886 3290
rect 216938 3238 216950 3290
rect 217002 3238 217014 3290
rect 217066 3238 217078 3290
rect 217130 3238 217142 3290
rect 217194 3238 217206 3290
rect 217258 3238 217270 3290
rect 217322 3238 217334 3290
rect 217386 3238 252822 3290
rect 252874 3238 252886 3290
rect 252938 3238 252950 3290
rect 253002 3238 253014 3290
rect 253066 3238 253078 3290
rect 253130 3238 253142 3290
rect 253194 3238 253206 3290
rect 253258 3238 253270 3290
rect 253322 3238 253334 3290
rect 253386 3238 288822 3290
rect 288874 3238 288886 3290
rect 288938 3238 288950 3290
rect 289002 3238 289014 3290
rect 289066 3238 289078 3290
rect 289130 3238 289142 3290
rect 289194 3238 289206 3290
rect 289258 3238 289270 3290
rect 289322 3238 289334 3290
rect 289386 3238 324822 3290
rect 324874 3238 324886 3290
rect 324938 3238 324950 3290
rect 325002 3238 325014 3290
rect 325066 3238 325078 3290
rect 325130 3238 325142 3290
rect 325194 3238 325206 3290
rect 325258 3238 325270 3290
rect 325322 3238 325334 3290
rect 325386 3238 360822 3290
rect 360874 3238 360886 3290
rect 360938 3238 360950 3290
rect 361002 3238 361014 3290
rect 361066 3238 361078 3290
rect 361130 3238 361142 3290
rect 361194 3238 361206 3290
rect 361258 3238 361270 3290
rect 361322 3238 361334 3290
rect 361386 3238 396822 3290
rect 396874 3238 396886 3290
rect 396938 3238 396950 3290
rect 397002 3238 397014 3290
rect 397066 3238 397078 3290
rect 397130 3238 397142 3290
rect 397194 3238 397206 3290
rect 397258 3238 397270 3290
rect 397322 3238 397334 3290
rect 397386 3238 432822 3290
rect 432874 3238 432886 3290
rect 432938 3238 432950 3290
rect 433002 3238 433014 3290
rect 433066 3238 433078 3290
rect 433130 3238 433142 3290
rect 433194 3238 433206 3290
rect 433258 3238 433270 3290
rect 433322 3238 433334 3290
rect 433386 3238 468822 3290
rect 468874 3238 468886 3290
rect 468938 3238 468950 3290
rect 469002 3238 469014 3290
rect 469066 3238 469078 3290
rect 469130 3238 469142 3290
rect 469194 3238 469206 3290
rect 469258 3238 469270 3290
rect 469322 3238 469334 3290
rect 469386 3238 504822 3290
rect 504874 3238 504886 3290
rect 504938 3238 504950 3290
rect 505002 3238 505014 3290
rect 505066 3238 505078 3290
rect 505130 3238 505142 3290
rect 505194 3238 505206 3290
rect 505258 3238 505270 3290
rect 505322 3238 505334 3290
rect 505386 3238 540822 3290
rect 540874 3238 540886 3290
rect 540938 3238 540950 3290
rect 541002 3238 541014 3290
rect 541066 3238 541078 3290
rect 541130 3238 541142 3290
rect 541194 3238 541206 3290
rect 541258 3238 541270 3290
rect 541322 3238 541334 3290
rect 541386 3238 576822 3290
rect 576874 3238 576886 3290
rect 576938 3238 576950 3290
rect 577002 3238 577014 3290
rect 577066 3238 577078 3290
rect 577130 3238 577142 3290
rect 577194 3238 577206 3290
rect 577258 3238 577270 3290
rect 577322 3238 577334 3290
rect 577386 3238 582820 3290
rect 1104 3216 582820 3238
rect 13630 3136 13636 3188
rect 13688 3176 13694 3188
rect 18598 3176 18604 3188
rect 13688 3148 18604 3176
rect 13688 3136 13694 3148
rect 18598 3136 18604 3148
rect 18656 3136 18662 3188
rect 23106 3136 23112 3188
rect 23164 3176 23170 3188
rect 27706 3176 27712 3188
rect 23164 3148 27712 3176
rect 23164 3136 23170 3148
rect 27706 3136 27712 3148
rect 27764 3136 27770 3188
rect 49326 3136 49332 3188
rect 49384 3176 49390 3188
rect 54662 3176 54668 3188
rect 49384 3148 54668 3176
rect 49384 3136 49390 3148
rect 54662 3136 54668 3148
rect 54720 3136 54726 3188
rect 56410 3136 56416 3188
rect 56468 3176 56474 3188
rect 61838 3176 61844 3188
rect 56468 3148 61844 3176
rect 56468 3136 56474 3148
rect 61838 3136 61844 3148
rect 61896 3136 61902 3188
rect 67174 3136 67180 3188
rect 67232 3176 67238 3188
rect 72050 3176 72056 3188
rect 67232 3148 72056 3176
rect 67232 3136 67238 3148
rect 72050 3136 72056 3148
rect 72108 3136 72114 3188
rect 273990 3136 273996 3188
rect 274048 3176 274054 3188
rect 276474 3176 276480 3188
rect 274048 3148 276480 3176
rect 274048 3136 274054 3148
rect 276474 3136 276480 3148
rect 276532 3136 276538 3188
rect 283190 3136 283196 3188
rect 283248 3176 283254 3188
rect 285950 3176 285956 3188
rect 283248 3148 285956 3176
rect 283248 3136 283254 3148
rect 285950 3136 285956 3148
rect 286008 3136 286014 3188
rect 307662 3136 307668 3188
rect 307720 3176 307726 3188
rect 310974 3176 310980 3188
rect 307720 3148 310980 3176
rect 307720 3136 307726 3148
rect 310974 3136 310980 3148
rect 311032 3136 311038 3188
rect 317230 3136 317236 3188
rect 317288 3176 317294 3188
rect 320450 3176 320456 3188
rect 317288 3148 320456 3176
rect 317288 3136 317294 3148
rect 320450 3136 320456 3148
rect 320508 3136 320514 3188
rect 326982 3136 326988 3188
rect 327040 3176 327046 3188
rect 331214 3176 331220 3188
rect 327040 3148 331220 3176
rect 327040 3136 327046 3148
rect 331214 3136 331220 3148
rect 331272 3136 331278 3188
rect 336642 3136 336648 3188
rect 336700 3176 336706 3188
rect 341886 3176 341892 3188
rect 336700 3148 341892 3176
rect 336700 3136 336706 3148
rect 341886 3136 341892 3148
rect 341944 3136 341950 3188
rect 345934 3136 345940 3188
rect 345992 3176 345998 3188
rect 351362 3176 351368 3188
rect 345992 3148 351368 3176
rect 345992 3136 345998 3148
rect 351362 3136 351368 3148
rect 351420 3136 351426 3188
rect 367094 3136 367100 3188
rect 367152 3176 367158 3188
rect 375190 3176 375196 3188
rect 367152 3148 375196 3176
rect 367152 3136 367158 3148
rect 375190 3136 375196 3148
rect 375248 3136 375254 3188
rect 414106 3136 414112 3188
rect 414164 3176 414170 3188
rect 415670 3176 415676 3188
rect 414164 3148 415676 3176
rect 414164 3136 414170 3148
rect 415670 3136 415676 3148
rect 415728 3136 415734 3188
rect 418154 3136 418160 3188
rect 418212 3176 418218 3188
rect 420362 3176 420368 3188
rect 418212 3148 420368 3176
rect 418212 3136 418218 3148
rect 420362 3136 420368 3148
rect 420420 3136 420426 3188
rect 427814 3136 427820 3188
rect 427872 3176 427878 3188
rect 429930 3176 429936 3188
rect 427872 3148 429936 3176
rect 427872 3136 427878 3148
rect 429930 3136 429936 3148
rect 429988 3136 429994 3188
rect 430574 3136 430580 3188
rect 430632 3176 430638 3188
rect 432322 3176 432328 3188
rect 430632 3148 432328 3176
rect 430632 3136 430638 3148
rect 432322 3136 432328 3148
rect 432380 3136 432386 3188
rect 438946 3136 438952 3188
rect 439004 3176 439010 3188
rect 440602 3176 440608 3188
rect 439004 3148 440608 3176
rect 439004 3136 439010 3148
rect 440602 3136 440608 3148
rect 440660 3136 440666 3188
rect 443546 3136 443552 3188
rect 443604 3176 443610 3188
rect 445386 3176 445392 3188
rect 443604 3148 445392 3176
rect 443604 3136 443610 3148
rect 445386 3136 445392 3148
rect 445444 3136 445450 3188
rect 448606 3136 448612 3188
rect 448664 3176 448670 3188
rect 451458 3176 451464 3188
rect 448664 3148 451464 3176
rect 448664 3136 448670 3148
rect 451458 3136 451464 3148
rect 451516 3136 451522 3188
rect 454126 3136 454132 3188
rect 454184 3176 454190 3188
rect 457254 3176 457260 3188
rect 454184 3148 457260 3176
rect 454184 3136 454190 3148
rect 457254 3136 457260 3148
rect 457312 3136 457318 3188
rect 458266 3136 458272 3188
rect 458324 3176 458330 3188
rect 460842 3176 460848 3188
rect 458324 3148 460848 3176
rect 458324 3136 458330 3148
rect 460842 3136 460848 3148
rect 460900 3136 460906 3188
rect 483290 3136 483296 3188
rect 483348 3176 483354 3188
rect 486694 3176 486700 3188
rect 483348 3148 486700 3176
rect 483348 3136 483354 3148
rect 486694 3136 486700 3148
rect 486752 3136 486758 3188
rect 514754 3136 514760 3188
rect 514812 3176 514818 3188
rect 520274 3176 520280 3188
rect 514812 3148 520280 3176
rect 514812 3136 514818 3148
rect 520274 3136 520280 3148
rect 520332 3136 520338 3188
rect 540238 3136 540244 3188
rect 540296 3176 540302 3188
rect 547690 3176 547696 3188
rect 540296 3148 547696 3176
rect 540296 3136 540302 3148
rect 547690 3136 547696 3148
rect 547748 3136 547754 3188
rect 557166 3176 557172 3188
rect 547800 3148 557172 3176
rect 2866 3068 2872 3120
rect 2924 3108 2930 3120
rect 5534 3108 5540 3120
rect 2924 3080 5540 3108
rect 2924 3068 2930 3080
rect 5534 3068 5540 3080
rect 5592 3068 5598 3120
rect 32674 3068 32680 3120
rect 32732 3108 32738 3120
rect 37458 3108 37464 3120
rect 32732 3080 37464 3108
rect 32732 3068 32738 3080
rect 37458 3068 37464 3080
rect 37516 3068 37522 3120
rect 46934 3068 46940 3120
rect 46992 3108 46998 3120
rect 52730 3108 52736 3120
rect 46992 3080 52736 3108
rect 46992 3068 46998 3080
rect 52730 3068 52736 3080
rect 52788 3068 52794 3120
rect 318242 3068 318248 3120
rect 318300 3108 318306 3120
rect 321646 3108 321652 3120
rect 318300 3080 321652 3108
rect 318300 3068 318306 3080
rect 321646 3068 321652 3080
rect 321704 3068 321710 3120
rect 330570 3068 330576 3120
rect 330628 3108 330634 3120
rect 335906 3108 335912 3120
rect 330628 3080 335912 3108
rect 330628 3068 330634 3080
rect 335906 3068 335912 3080
rect 335964 3068 335970 3120
rect 339678 3068 339684 3120
rect 339736 3108 339742 3120
rect 345474 3108 345480 3120
rect 339736 3080 345480 3108
rect 339736 3068 339742 3080
rect 345474 3068 345480 3080
rect 345532 3068 345538 3120
rect 424318 3068 424324 3120
rect 424376 3108 424382 3120
rect 426342 3108 426348 3120
rect 424376 3080 426348 3108
rect 424376 3068 424382 3080
rect 426342 3068 426348 3080
rect 426400 3068 426406 3120
rect 438854 3068 438860 3120
rect 438912 3108 438918 3120
rect 441798 3108 441804 3120
rect 438912 3080 441804 3108
rect 438912 3068 438918 3080
rect 441798 3068 441804 3080
rect 441856 3068 441862 3120
rect 447134 3068 447140 3120
rect 447192 3108 447198 3120
rect 450170 3108 450176 3120
rect 447192 3080 450176 3108
rect 447192 3068 447198 3080
rect 450170 3068 450176 3080
rect 450228 3068 450234 3120
rect 454678 3068 454684 3120
rect 454736 3108 454742 3120
rect 458450 3108 458456 3120
rect 454736 3080 458456 3108
rect 454736 3068 454742 3080
rect 458450 3068 458456 3080
rect 458508 3068 458514 3120
rect 463694 3068 463700 3120
rect 463752 3108 463758 3120
rect 466822 3108 466828 3120
rect 463752 3080 466828 3108
rect 463752 3068 463758 3080
rect 466822 3068 466828 3080
rect 466880 3068 466886 3120
rect 484670 3068 484676 3120
rect 484728 3108 484734 3120
rect 490558 3108 490564 3120
rect 484728 3080 490564 3108
rect 484728 3068 484734 3080
rect 490558 3068 490564 3080
rect 490616 3068 490622 3120
rect 500586 3068 500592 3120
rect 500644 3108 500650 3120
rect 504726 3108 504732 3120
rect 500644 3080 504732 3108
rect 500644 3068 500650 3080
rect 504726 3068 504732 3080
rect 504784 3068 504790 3120
rect 526622 3068 526628 3120
rect 526680 3108 526686 3120
rect 544102 3108 544108 3120
rect 526680 3080 544108 3108
rect 526680 3068 526686 3080
rect 544102 3068 544108 3080
rect 544160 3068 544166 3120
rect 544197 3111 544255 3117
rect 544197 3077 544209 3111
rect 544243 3108 544255 3111
rect 547800 3108 547828 3148
rect 557166 3136 557172 3148
rect 557224 3136 557230 3188
rect 567105 3179 567163 3185
rect 567105 3145 567117 3179
rect 567151 3176 567163 3179
rect 575014 3176 575020 3188
rect 567151 3148 575020 3176
rect 567151 3145 567163 3148
rect 567105 3139 567163 3145
rect 575014 3136 575020 3148
rect 575072 3136 575078 3188
rect 544243 3080 547828 3108
rect 547877 3111 547935 3117
rect 544243 3077 544255 3080
rect 544197 3071 544255 3077
rect 547877 3077 547889 3111
rect 547923 3108 547935 3111
rect 555970 3108 555976 3120
rect 547923 3080 555976 3108
rect 547923 3077 547935 3080
rect 547877 3071 547935 3077
rect 555970 3068 555976 3080
rect 556028 3068 556034 3120
rect 556154 3068 556160 3120
rect 556212 3108 556218 3120
rect 558089 3111 558147 3117
rect 558089 3108 558101 3111
rect 556212 3080 558101 3108
rect 556212 3068 556218 3080
rect 558089 3077 558101 3080
rect 558135 3077 558147 3111
rect 558089 3071 558147 3077
rect 558181 3111 558239 3117
rect 558181 3077 558193 3111
rect 558227 3108 558239 3111
rect 560849 3111 560907 3117
rect 560849 3108 560861 3111
rect 558227 3080 560861 3108
rect 558227 3077 558239 3080
rect 558181 3071 558239 3077
rect 560849 3077 560861 3080
rect 560895 3077 560907 3111
rect 566734 3108 566740 3120
rect 560849 3071 560907 3077
rect 560956 3080 566740 3108
rect 12434 3000 12440 3052
rect 12492 3040 12498 3052
rect 18046 3040 18052 3052
rect 12492 3012 18052 3040
rect 12492 3000 12498 3012
rect 18046 3000 18052 3012
rect 18104 3000 18110 3052
rect 269666 3000 269672 3052
rect 269724 3040 269730 3052
rect 271690 3040 271696 3052
rect 269724 3012 271696 3040
rect 269724 3000 269730 3012
rect 271690 3000 271696 3012
rect 271748 3000 271754 3052
rect 271874 3000 271880 3052
rect 271932 3040 271938 3052
rect 274082 3040 274088 3052
rect 271932 3012 274088 3040
rect 271932 3000 271938 3012
rect 274082 3000 274088 3012
rect 274140 3000 274146 3052
rect 279326 3000 279332 3052
rect 279384 3040 279390 3052
rect 281258 3040 281264 3052
rect 279384 3012 281264 3040
rect 279384 3000 279390 3012
rect 281258 3000 281264 3012
rect 281316 3000 281322 3052
rect 298922 3000 298928 3052
rect 298980 3040 298986 3052
rect 301406 3040 301412 3052
rect 298980 3012 301412 3040
rect 298980 3000 298986 3012
rect 301406 3000 301412 3012
rect 301464 3000 301470 3052
rect 318702 3000 318708 3052
rect 318760 3040 318766 3052
rect 322842 3040 322848 3052
rect 318760 3012 322848 3040
rect 318760 3000 318766 3012
rect 322842 3000 322848 3012
rect 322900 3000 322906 3052
rect 328270 3000 328276 3052
rect 328328 3040 328334 3052
rect 332410 3040 332416 3052
rect 328328 3012 332416 3040
rect 328328 3000 328334 3012
rect 332410 3000 332416 3012
rect 332468 3000 332474 3052
rect 347406 3000 347412 3052
rect 347464 3040 347470 3052
rect 352558 3040 352564 3052
rect 347464 3012 352564 3040
rect 347464 3000 347470 3012
rect 352558 3000 352564 3012
rect 352616 3000 352622 3052
rect 403802 3000 403808 3052
rect 403860 3040 403866 3052
rect 404906 3040 404912 3052
rect 403860 3012 404912 3040
rect 403860 3000 403866 3012
rect 404906 3000 404912 3012
rect 404964 3000 404970 3052
rect 439038 3000 439044 3052
rect 439096 3040 439102 3052
rect 442994 3040 443000 3052
rect 439096 3012 443000 3040
rect 439096 3000 439102 3012
rect 442994 3000 443000 3012
rect 443052 3000 443058 3052
rect 444374 3000 444380 3052
rect 444432 3040 444438 3052
rect 446582 3040 446588 3052
rect 444432 3012 446588 3040
rect 444432 3000 444438 3012
rect 446582 3000 446588 3012
rect 446640 3000 446646 3052
rect 464246 3000 464252 3052
rect 464304 3040 464310 3052
rect 468662 3040 468668 3052
rect 464304 3012 468668 3040
rect 464304 3000 464310 3012
rect 468662 3000 468668 3012
rect 468720 3000 468726 3052
rect 494146 3000 494152 3052
rect 494204 3040 494210 3052
rect 498930 3040 498936 3052
rect 494204 3012 498936 3040
rect 494204 3000 494210 3012
rect 498930 3000 498936 3012
rect 498988 3000 498994 3052
rect 503990 3000 503996 3052
rect 504048 3040 504054 3052
rect 508406 3040 508412 3052
rect 504048 3012 508412 3040
rect 504048 3000 504054 3012
rect 508406 3000 508412 3012
rect 508464 3000 508470 3052
rect 521194 3000 521200 3052
rect 521252 3040 521258 3052
rect 526254 3040 526260 3052
rect 521252 3012 526260 3040
rect 521252 3000 521258 3012
rect 526254 3000 526260 3012
rect 526312 3000 526318 3052
rect 536834 3000 536840 3052
rect 536892 3040 536898 3052
rect 547969 3043 548027 3049
rect 547969 3040 547981 3043
rect 536892 3012 547981 3040
rect 536892 3000 536898 3012
rect 547969 3009 547981 3012
rect 548015 3009 548027 3043
rect 560956 3040 560984 3080
rect 566734 3068 566740 3080
rect 566792 3068 566798 3120
rect 566829 3111 566887 3117
rect 566829 3077 566841 3111
rect 566875 3108 566887 3111
rect 573818 3108 573824 3120
rect 566875 3080 573824 3108
rect 566875 3077 566887 3080
rect 566829 3071 566887 3077
rect 573818 3068 573824 3080
rect 573876 3068 573882 3120
rect 547969 3003 548027 3009
rect 554884 3012 560984 3040
rect 37458 2932 37464 2984
rect 37516 2972 37522 2984
rect 43714 2972 43720 2984
rect 37516 2944 43720 2972
rect 37516 2932 37522 2944
rect 43714 2932 43720 2944
rect 43772 2932 43778 2984
rect 260098 2932 260104 2984
rect 260156 2972 260162 2984
rect 262214 2972 262220 2984
rect 260156 2944 262220 2972
rect 260156 2932 260162 2944
rect 262214 2932 262220 2944
rect 262272 2932 262278 2984
rect 337378 2932 337384 2984
rect 337436 2972 337442 2984
rect 342714 2972 342720 2984
rect 337436 2944 342720 2972
rect 337436 2932 337442 2944
rect 342714 2932 342720 2944
rect 342772 2932 342778 2984
rect 511902 2932 511908 2984
rect 511960 2972 511966 2984
rect 516778 2972 516784 2984
rect 511960 2944 516784 2972
rect 511960 2932 511966 2944
rect 516778 2932 516784 2944
rect 516836 2932 516842 2984
rect 522390 2932 522396 2984
rect 522448 2972 522454 2984
rect 527450 2972 527456 2984
rect 522448 2944 527456 2972
rect 522448 2932 522454 2944
rect 527450 2932 527456 2944
rect 527508 2932 527514 2984
rect 536742 2932 536748 2984
rect 536800 2972 536806 2984
rect 541710 2972 541716 2984
rect 536800 2944 541716 2972
rect 536800 2932 536806 2944
rect 541710 2932 541716 2944
rect 541768 2932 541774 2984
rect 541805 2975 541863 2981
rect 541805 2941 541817 2975
rect 541851 2972 541863 2975
rect 552382 2972 552388 2984
rect 541851 2944 552388 2972
rect 541851 2941 541863 2944
rect 541805 2935 541863 2941
rect 552382 2932 552388 2944
rect 552440 2932 552446 2984
rect 554884 2972 554912 3012
rect 552492 2944 554912 2972
rect 1670 2864 1676 2916
rect 1728 2904 1734 2916
rect 9582 2904 9588 2916
rect 1728 2876 9588 2904
rect 1728 2864 1734 2876
rect 9582 2864 9588 2876
rect 9640 2864 9646 2916
rect 10042 2864 10048 2916
rect 10100 2904 10106 2916
rect 15194 2904 15200 2916
rect 10100 2876 15200 2904
rect 10100 2864 10106 2876
rect 15194 2864 15200 2876
rect 15252 2864 15258 2916
rect 240134 2864 240140 2916
rect 240192 2904 240198 2916
rect 241974 2904 241980 2916
rect 240192 2876 241980 2904
rect 240192 2864 240198 2876
rect 241974 2864 241980 2876
rect 242032 2864 242038 2916
rect 249242 2864 249248 2916
rect 249300 2904 249306 2916
rect 250346 2904 250352 2916
rect 249300 2876 250352 2904
rect 249300 2864 249306 2876
rect 250346 2864 250352 2876
rect 250404 2864 250410 2916
rect 258994 2864 259000 2916
rect 259052 2904 259058 2916
rect 259822 2904 259828 2916
rect 259052 2876 259828 2904
rect 259052 2864 259058 2876
rect 259822 2864 259828 2876
rect 259880 2864 259886 2916
rect 269022 2864 269028 2916
rect 269080 2904 269086 2916
rect 270494 2904 270500 2916
rect 269080 2876 270500 2904
rect 269080 2864 269086 2876
rect 270494 2864 270500 2876
rect 270552 2864 270558 2916
rect 288250 2864 288256 2916
rect 288308 2904 288314 2916
rect 290734 2904 290740 2916
rect 288308 2876 290740 2904
rect 288308 2864 288314 2876
rect 290734 2864 290740 2876
rect 290792 2864 290798 2916
rect 297818 2864 297824 2916
rect 297876 2904 297882 2916
rect 300302 2904 300308 2916
rect 297876 2876 300308 2904
rect 297876 2864 297882 2876
rect 300302 2864 300308 2876
rect 300360 2864 300366 2916
rect 384942 2864 384948 2916
rect 385000 2904 385006 2916
rect 391842 2904 391848 2916
rect 385000 2876 391848 2904
rect 385000 2864 385006 2876
rect 391842 2864 391848 2876
rect 391900 2864 391906 2916
rect 491110 2864 491116 2916
rect 491168 2904 491174 2916
rect 494146 2904 494152 2916
rect 491168 2876 494152 2904
rect 491168 2864 491174 2876
rect 494146 2864 494152 2876
rect 494204 2864 494210 2916
rect 528922 2864 528928 2916
rect 528980 2904 528986 2916
rect 546494 2904 546500 2916
rect 528980 2876 546500 2904
rect 528980 2864 528986 2876
rect 546494 2864 546500 2876
rect 546552 2864 546558 2916
rect 546586 2864 546592 2916
rect 546644 2904 546650 2916
rect 547690 2904 547696 2916
rect 546644 2876 547696 2904
rect 546644 2864 546650 2876
rect 547690 2864 547696 2876
rect 547748 2864 547754 2916
rect 548150 2864 548156 2916
rect 548208 2904 548214 2916
rect 552492 2904 552520 2944
rect 554958 2932 554964 2984
rect 555016 2972 555022 2984
rect 560757 2975 560815 2981
rect 560757 2972 560769 2975
rect 555016 2944 560769 2972
rect 555016 2932 555022 2944
rect 560757 2941 560769 2944
rect 560803 2941 560815 2975
rect 560757 2935 560815 2941
rect 561125 2975 561183 2981
rect 561125 2941 561137 2975
rect 561171 2972 561183 2975
rect 564342 2972 564348 2984
rect 561171 2944 564348 2972
rect 561171 2941 561183 2944
rect 561125 2935 561183 2941
rect 564342 2932 564348 2944
rect 564400 2932 564406 2984
rect 564437 2975 564495 2981
rect 564437 2941 564449 2975
rect 564483 2972 564495 2975
rect 572622 2972 572628 2984
rect 564483 2944 572628 2972
rect 564483 2941 564495 2944
rect 564437 2935 564495 2941
rect 572622 2932 572628 2944
rect 572680 2932 572686 2984
rect 548208 2876 552520 2904
rect 552661 2907 552719 2913
rect 548208 2864 548214 2876
rect 552661 2873 552673 2907
rect 552707 2904 552719 2907
rect 565538 2904 565544 2916
rect 552707 2876 565544 2904
rect 552707 2873 552719 2876
rect 552661 2867 552719 2873
rect 565538 2864 565544 2876
rect 565596 2864 565602 2916
rect 565633 2907 565691 2913
rect 565633 2873 565645 2907
rect 565679 2904 565691 2907
rect 566829 2907 566887 2913
rect 566829 2904 566841 2907
rect 565679 2876 566841 2904
rect 565679 2873 565691 2876
rect 565633 2867 565691 2873
rect 566829 2873 566841 2876
rect 566875 2873 566887 2907
rect 566829 2867 566887 2873
rect 19518 2796 19524 2848
rect 19576 2836 19582 2848
rect 26142 2836 26148 2848
rect 19576 2808 26148 2836
rect 19576 2796 19582 2808
rect 26142 2796 26148 2808
rect 26200 2796 26206 2848
rect 30282 2796 30288 2848
rect 30340 2836 30346 2848
rect 34514 2836 34520 2848
rect 30340 2808 34520 2836
rect 30340 2796 30346 2808
rect 34514 2796 34520 2808
rect 34572 2796 34578 2848
rect 39758 2796 39764 2848
rect 39816 2836 39822 2848
rect 45462 2836 45468 2848
rect 39816 2808 45468 2836
rect 39816 2796 39822 2808
rect 45462 2796 45468 2808
rect 45520 2796 45526 2848
rect 278406 2796 278412 2848
rect 278464 2836 278470 2848
rect 280062 2836 280068 2848
rect 278464 2808 280068 2836
rect 278464 2796 278470 2808
rect 280062 2796 280068 2808
rect 280120 2796 280126 2848
rect 308214 2796 308220 2848
rect 308272 2836 308278 2848
rect 312170 2836 312176 2848
rect 308272 2808 312176 2836
rect 308272 2796 308278 2808
rect 312170 2796 312176 2808
rect 312228 2796 312234 2848
rect 355502 2796 355508 2848
rect 355560 2836 355566 2848
rect 360746 2836 360752 2848
rect 355560 2808 360752 2836
rect 355560 2796 355566 2808
rect 360746 2796 360752 2808
rect 360804 2796 360810 2848
rect 532326 2796 532332 2848
rect 532384 2836 532390 2848
rect 550082 2836 550088 2848
rect 532384 2808 550088 2836
rect 532384 2796 532390 2808
rect 550082 2796 550088 2808
rect 550140 2796 550146 2848
rect 550542 2796 550548 2848
rect 550600 2836 550606 2848
rect 567838 2836 567844 2848
rect 550600 2808 567844 2836
rect 550600 2796 550606 2808
rect 567838 2796 567844 2808
rect 567896 2796 567902 2848
rect 1104 2746 582820 2768
rect 1104 2694 18822 2746
rect 18874 2694 18886 2746
rect 18938 2694 18950 2746
rect 19002 2694 19014 2746
rect 19066 2694 19078 2746
rect 19130 2694 19142 2746
rect 19194 2694 19206 2746
rect 19258 2694 19270 2746
rect 19322 2694 19334 2746
rect 19386 2694 54822 2746
rect 54874 2694 54886 2746
rect 54938 2694 54950 2746
rect 55002 2694 55014 2746
rect 55066 2694 55078 2746
rect 55130 2694 55142 2746
rect 55194 2694 55206 2746
rect 55258 2694 55270 2746
rect 55322 2694 55334 2746
rect 55386 2694 90822 2746
rect 90874 2694 90886 2746
rect 90938 2694 90950 2746
rect 91002 2694 91014 2746
rect 91066 2694 91078 2746
rect 91130 2694 91142 2746
rect 91194 2694 91206 2746
rect 91258 2694 91270 2746
rect 91322 2694 91334 2746
rect 91386 2694 126822 2746
rect 126874 2694 126886 2746
rect 126938 2694 126950 2746
rect 127002 2694 127014 2746
rect 127066 2694 127078 2746
rect 127130 2694 127142 2746
rect 127194 2694 127206 2746
rect 127258 2694 127270 2746
rect 127322 2694 127334 2746
rect 127386 2694 162822 2746
rect 162874 2694 162886 2746
rect 162938 2694 162950 2746
rect 163002 2694 163014 2746
rect 163066 2694 163078 2746
rect 163130 2694 163142 2746
rect 163194 2694 163206 2746
rect 163258 2694 163270 2746
rect 163322 2694 163334 2746
rect 163386 2694 198822 2746
rect 198874 2694 198886 2746
rect 198938 2694 198950 2746
rect 199002 2694 199014 2746
rect 199066 2694 199078 2746
rect 199130 2694 199142 2746
rect 199194 2694 199206 2746
rect 199258 2694 199270 2746
rect 199322 2694 199334 2746
rect 199386 2694 234822 2746
rect 234874 2694 234886 2746
rect 234938 2694 234950 2746
rect 235002 2694 235014 2746
rect 235066 2694 235078 2746
rect 235130 2694 235142 2746
rect 235194 2694 235206 2746
rect 235258 2694 235270 2746
rect 235322 2694 235334 2746
rect 235386 2694 270822 2746
rect 270874 2694 270886 2746
rect 270938 2694 270950 2746
rect 271002 2694 271014 2746
rect 271066 2694 271078 2746
rect 271130 2694 271142 2746
rect 271194 2694 271206 2746
rect 271258 2694 271270 2746
rect 271322 2694 271334 2746
rect 271386 2694 306822 2746
rect 306874 2694 306886 2746
rect 306938 2694 306950 2746
rect 307002 2694 307014 2746
rect 307066 2694 307078 2746
rect 307130 2694 307142 2746
rect 307194 2694 307206 2746
rect 307258 2694 307270 2746
rect 307322 2694 307334 2746
rect 307386 2694 342822 2746
rect 342874 2694 342886 2746
rect 342938 2694 342950 2746
rect 343002 2694 343014 2746
rect 343066 2694 343078 2746
rect 343130 2694 343142 2746
rect 343194 2694 343206 2746
rect 343258 2694 343270 2746
rect 343322 2694 343334 2746
rect 343386 2694 378822 2746
rect 378874 2694 378886 2746
rect 378938 2694 378950 2746
rect 379002 2694 379014 2746
rect 379066 2694 379078 2746
rect 379130 2694 379142 2746
rect 379194 2694 379206 2746
rect 379258 2694 379270 2746
rect 379322 2694 379334 2746
rect 379386 2694 414822 2746
rect 414874 2694 414886 2746
rect 414938 2694 414950 2746
rect 415002 2694 415014 2746
rect 415066 2694 415078 2746
rect 415130 2694 415142 2746
rect 415194 2694 415206 2746
rect 415258 2694 415270 2746
rect 415322 2694 415334 2746
rect 415386 2694 450822 2746
rect 450874 2694 450886 2746
rect 450938 2694 450950 2746
rect 451002 2694 451014 2746
rect 451066 2694 451078 2746
rect 451130 2694 451142 2746
rect 451194 2694 451206 2746
rect 451258 2694 451270 2746
rect 451322 2694 451334 2746
rect 451386 2694 486822 2746
rect 486874 2694 486886 2746
rect 486938 2694 486950 2746
rect 487002 2694 487014 2746
rect 487066 2694 487078 2746
rect 487130 2694 487142 2746
rect 487194 2694 487206 2746
rect 487258 2694 487270 2746
rect 487322 2694 487334 2746
rect 487386 2694 522822 2746
rect 522874 2694 522886 2746
rect 522938 2694 522950 2746
rect 523002 2694 523014 2746
rect 523066 2694 523078 2746
rect 523130 2694 523142 2746
rect 523194 2694 523206 2746
rect 523258 2694 523270 2746
rect 523322 2694 523334 2746
rect 523386 2694 558822 2746
rect 558874 2694 558886 2746
rect 558938 2694 558950 2746
rect 559002 2694 559014 2746
rect 559066 2694 559078 2746
rect 559130 2694 559142 2746
rect 559194 2694 559206 2746
rect 559258 2694 559270 2746
rect 559322 2694 559334 2746
rect 559386 2694 582820 2746
rect 1104 2672 582820 2694
rect 547969 2635 548027 2641
rect 547969 2601 547981 2635
rect 548015 2632 548027 2635
rect 554774 2632 554780 2644
rect 548015 2604 554780 2632
rect 548015 2601 548027 2604
rect 547969 2595 548027 2601
rect 554774 2592 554780 2604
rect 554832 2592 554838 2644
rect 560757 2635 560815 2641
rect 560757 2601 560769 2635
rect 560803 2632 560815 2635
rect 565633 2635 565691 2641
rect 565633 2632 565645 2635
rect 560803 2604 565645 2632
rect 560803 2601 560815 2604
rect 560757 2595 560815 2601
rect 565633 2601 565645 2604
rect 565679 2601 565691 2635
rect 565633 2595 565691 2601
rect 1104 2202 582820 2224
rect 1104 2150 36822 2202
rect 36874 2150 36886 2202
rect 36938 2150 36950 2202
rect 37002 2150 37014 2202
rect 37066 2150 37078 2202
rect 37130 2150 37142 2202
rect 37194 2150 37206 2202
rect 37258 2150 37270 2202
rect 37322 2150 37334 2202
rect 37386 2150 72822 2202
rect 72874 2150 72886 2202
rect 72938 2150 72950 2202
rect 73002 2150 73014 2202
rect 73066 2150 73078 2202
rect 73130 2150 73142 2202
rect 73194 2150 73206 2202
rect 73258 2150 73270 2202
rect 73322 2150 73334 2202
rect 73386 2150 108822 2202
rect 108874 2150 108886 2202
rect 108938 2150 108950 2202
rect 109002 2150 109014 2202
rect 109066 2150 109078 2202
rect 109130 2150 109142 2202
rect 109194 2150 109206 2202
rect 109258 2150 109270 2202
rect 109322 2150 109334 2202
rect 109386 2150 144822 2202
rect 144874 2150 144886 2202
rect 144938 2150 144950 2202
rect 145002 2150 145014 2202
rect 145066 2150 145078 2202
rect 145130 2150 145142 2202
rect 145194 2150 145206 2202
rect 145258 2150 145270 2202
rect 145322 2150 145334 2202
rect 145386 2150 180822 2202
rect 180874 2150 180886 2202
rect 180938 2150 180950 2202
rect 181002 2150 181014 2202
rect 181066 2150 181078 2202
rect 181130 2150 181142 2202
rect 181194 2150 181206 2202
rect 181258 2150 181270 2202
rect 181322 2150 181334 2202
rect 181386 2150 216822 2202
rect 216874 2150 216886 2202
rect 216938 2150 216950 2202
rect 217002 2150 217014 2202
rect 217066 2150 217078 2202
rect 217130 2150 217142 2202
rect 217194 2150 217206 2202
rect 217258 2150 217270 2202
rect 217322 2150 217334 2202
rect 217386 2150 252822 2202
rect 252874 2150 252886 2202
rect 252938 2150 252950 2202
rect 253002 2150 253014 2202
rect 253066 2150 253078 2202
rect 253130 2150 253142 2202
rect 253194 2150 253206 2202
rect 253258 2150 253270 2202
rect 253322 2150 253334 2202
rect 253386 2150 288822 2202
rect 288874 2150 288886 2202
rect 288938 2150 288950 2202
rect 289002 2150 289014 2202
rect 289066 2150 289078 2202
rect 289130 2150 289142 2202
rect 289194 2150 289206 2202
rect 289258 2150 289270 2202
rect 289322 2150 289334 2202
rect 289386 2150 324822 2202
rect 324874 2150 324886 2202
rect 324938 2150 324950 2202
rect 325002 2150 325014 2202
rect 325066 2150 325078 2202
rect 325130 2150 325142 2202
rect 325194 2150 325206 2202
rect 325258 2150 325270 2202
rect 325322 2150 325334 2202
rect 325386 2150 360822 2202
rect 360874 2150 360886 2202
rect 360938 2150 360950 2202
rect 361002 2150 361014 2202
rect 361066 2150 361078 2202
rect 361130 2150 361142 2202
rect 361194 2150 361206 2202
rect 361258 2150 361270 2202
rect 361322 2150 361334 2202
rect 361386 2150 396822 2202
rect 396874 2150 396886 2202
rect 396938 2150 396950 2202
rect 397002 2150 397014 2202
rect 397066 2150 397078 2202
rect 397130 2150 397142 2202
rect 397194 2150 397206 2202
rect 397258 2150 397270 2202
rect 397322 2150 397334 2202
rect 397386 2150 432822 2202
rect 432874 2150 432886 2202
rect 432938 2150 432950 2202
rect 433002 2150 433014 2202
rect 433066 2150 433078 2202
rect 433130 2150 433142 2202
rect 433194 2150 433206 2202
rect 433258 2150 433270 2202
rect 433322 2150 433334 2202
rect 433386 2150 468822 2202
rect 468874 2150 468886 2202
rect 468938 2150 468950 2202
rect 469002 2150 469014 2202
rect 469066 2150 469078 2202
rect 469130 2150 469142 2202
rect 469194 2150 469206 2202
rect 469258 2150 469270 2202
rect 469322 2150 469334 2202
rect 469386 2150 504822 2202
rect 504874 2150 504886 2202
rect 504938 2150 504950 2202
rect 505002 2150 505014 2202
rect 505066 2150 505078 2202
rect 505130 2150 505142 2202
rect 505194 2150 505206 2202
rect 505258 2150 505270 2202
rect 505322 2150 505334 2202
rect 505386 2150 540822 2202
rect 540874 2150 540886 2202
rect 540938 2150 540950 2202
rect 541002 2150 541014 2202
rect 541066 2150 541078 2202
rect 541130 2150 541142 2202
rect 541194 2150 541206 2202
rect 541258 2150 541270 2202
rect 541322 2150 541334 2202
rect 541386 2150 576822 2202
rect 576874 2150 576886 2202
rect 576938 2150 576950 2202
rect 577002 2150 577014 2202
rect 577066 2150 577078 2202
rect 577130 2150 577142 2202
rect 577194 2150 577206 2202
rect 577258 2150 577270 2202
rect 577322 2150 577334 2202
rect 577386 2150 582820 2202
rect 1104 2128 582820 2150
<< via1 >>
rect 251640 701972 251692 702024
rect 429844 701972 429896 702024
rect 237472 701904 237524 701956
rect 494796 701904 494848 701956
rect 223304 701836 223356 701888
rect 559656 701836 559708 701888
rect 36822 701734 36874 701786
rect 36886 701734 36938 701786
rect 36950 701734 37002 701786
rect 37014 701734 37066 701786
rect 37078 701734 37130 701786
rect 37142 701734 37194 701786
rect 37206 701734 37258 701786
rect 37270 701734 37322 701786
rect 37334 701734 37386 701786
rect 72822 701734 72874 701786
rect 72886 701734 72938 701786
rect 72950 701734 73002 701786
rect 73014 701734 73066 701786
rect 73078 701734 73130 701786
rect 73142 701734 73194 701786
rect 73206 701734 73258 701786
rect 73270 701734 73322 701786
rect 73334 701734 73386 701786
rect 108822 701734 108874 701786
rect 108886 701734 108938 701786
rect 108950 701734 109002 701786
rect 109014 701734 109066 701786
rect 109078 701734 109130 701786
rect 109142 701734 109194 701786
rect 109206 701734 109258 701786
rect 109270 701734 109322 701786
rect 109334 701734 109386 701786
rect 144822 701734 144874 701786
rect 144886 701734 144938 701786
rect 144950 701734 145002 701786
rect 145014 701734 145066 701786
rect 145078 701734 145130 701786
rect 145142 701734 145194 701786
rect 145206 701734 145258 701786
rect 145270 701734 145322 701786
rect 145334 701734 145386 701786
rect 180822 701734 180874 701786
rect 180886 701734 180938 701786
rect 180950 701734 181002 701786
rect 181014 701734 181066 701786
rect 181078 701734 181130 701786
rect 181142 701734 181194 701786
rect 181206 701734 181258 701786
rect 181270 701734 181322 701786
rect 181334 701734 181386 701786
rect 216822 701734 216874 701786
rect 216886 701734 216938 701786
rect 216950 701734 217002 701786
rect 217014 701734 217066 701786
rect 217078 701734 217130 701786
rect 217142 701734 217194 701786
rect 217206 701734 217258 701786
rect 217270 701734 217322 701786
rect 217334 701734 217386 701786
rect 252822 701734 252874 701786
rect 252886 701734 252938 701786
rect 252950 701734 253002 701786
rect 253014 701734 253066 701786
rect 253078 701734 253130 701786
rect 253142 701734 253194 701786
rect 253206 701734 253258 701786
rect 253270 701734 253322 701786
rect 253334 701734 253386 701786
rect 288822 701734 288874 701786
rect 288886 701734 288938 701786
rect 288950 701734 289002 701786
rect 289014 701734 289066 701786
rect 289078 701734 289130 701786
rect 289142 701734 289194 701786
rect 289206 701734 289258 701786
rect 289270 701734 289322 701786
rect 289334 701734 289386 701786
rect 324822 701734 324874 701786
rect 324886 701734 324938 701786
rect 324950 701734 325002 701786
rect 325014 701734 325066 701786
rect 325078 701734 325130 701786
rect 325142 701734 325194 701786
rect 325206 701734 325258 701786
rect 325270 701734 325322 701786
rect 325334 701734 325386 701786
rect 360822 701734 360874 701786
rect 360886 701734 360938 701786
rect 360950 701734 361002 701786
rect 361014 701734 361066 701786
rect 361078 701734 361130 701786
rect 361142 701734 361194 701786
rect 361206 701734 361258 701786
rect 361270 701734 361322 701786
rect 361334 701734 361386 701786
rect 396822 701734 396874 701786
rect 396886 701734 396938 701786
rect 396950 701734 397002 701786
rect 397014 701734 397066 701786
rect 397078 701734 397130 701786
rect 397142 701734 397194 701786
rect 397206 701734 397258 701786
rect 397270 701734 397322 701786
rect 397334 701734 397386 701786
rect 432822 701734 432874 701786
rect 432886 701734 432938 701786
rect 432950 701734 433002 701786
rect 433014 701734 433066 701786
rect 433078 701734 433130 701786
rect 433142 701734 433194 701786
rect 433206 701734 433258 701786
rect 433270 701734 433322 701786
rect 433334 701734 433386 701786
rect 468822 701734 468874 701786
rect 468886 701734 468938 701786
rect 468950 701734 469002 701786
rect 469014 701734 469066 701786
rect 469078 701734 469130 701786
rect 469142 701734 469194 701786
rect 469206 701734 469258 701786
rect 469270 701734 469322 701786
rect 469334 701734 469386 701786
rect 504822 701734 504874 701786
rect 504886 701734 504938 701786
rect 504950 701734 505002 701786
rect 505014 701734 505066 701786
rect 505078 701734 505130 701786
rect 505142 701734 505194 701786
rect 505206 701734 505258 701786
rect 505270 701734 505322 701786
rect 505334 701734 505386 701786
rect 540822 701734 540874 701786
rect 540886 701734 540938 701786
rect 540950 701734 541002 701786
rect 541014 701734 541066 701786
rect 541078 701734 541130 701786
rect 541142 701734 541194 701786
rect 541206 701734 541258 701786
rect 541270 701734 541322 701786
rect 541334 701734 541386 701786
rect 576822 701734 576874 701786
rect 576886 701734 576938 701786
rect 576950 701734 577002 701786
rect 577014 701734 577066 701786
rect 577078 701734 577130 701786
rect 577142 701734 577194 701786
rect 577206 701734 577258 701786
rect 577270 701734 577322 701786
rect 577334 701734 577386 701786
rect 235172 701632 235224 701684
rect 18822 701190 18874 701242
rect 18886 701190 18938 701242
rect 18950 701190 19002 701242
rect 19014 701190 19066 701242
rect 19078 701190 19130 701242
rect 19142 701190 19194 701242
rect 19206 701190 19258 701242
rect 19270 701190 19322 701242
rect 19334 701190 19386 701242
rect 54822 701190 54874 701242
rect 54886 701190 54938 701242
rect 54950 701190 55002 701242
rect 55014 701190 55066 701242
rect 55078 701190 55130 701242
rect 55142 701190 55194 701242
rect 55206 701190 55258 701242
rect 55270 701190 55322 701242
rect 55334 701190 55386 701242
rect 90822 701190 90874 701242
rect 90886 701190 90938 701242
rect 90950 701190 91002 701242
rect 91014 701190 91066 701242
rect 91078 701190 91130 701242
rect 91142 701190 91194 701242
rect 91206 701190 91258 701242
rect 91270 701190 91322 701242
rect 91334 701190 91386 701242
rect 126822 701190 126874 701242
rect 126886 701190 126938 701242
rect 126950 701190 127002 701242
rect 127014 701190 127066 701242
rect 127078 701190 127130 701242
rect 127142 701190 127194 701242
rect 127206 701190 127258 701242
rect 127270 701190 127322 701242
rect 127334 701190 127386 701242
rect 162822 701190 162874 701242
rect 162886 701190 162938 701242
rect 162950 701190 163002 701242
rect 163014 701190 163066 701242
rect 163078 701190 163130 701242
rect 163142 701190 163194 701242
rect 163206 701190 163258 701242
rect 163270 701190 163322 701242
rect 163334 701190 163386 701242
rect 198822 701190 198874 701242
rect 198886 701190 198938 701242
rect 198950 701190 199002 701242
rect 199014 701190 199066 701242
rect 199078 701190 199130 701242
rect 199142 701190 199194 701242
rect 199206 701190 199258 701242
rect 199270 701190 199322 701242
rect 199334 701190 199386 701242
rect 234822 701190 234874 701242
rect 234886 701190 234938 701242
rect 234950 701190 235002 701242
rect 235014 701190 235066 701242
rect 235078 701190 235130 701242
rect 235142 701190 235194 701242
rect 235206 701190 235258 701242
rect 235270 701190 235322 701242
rect 235334 701190 235386 701242
rect 270822 701190 270874 701242
rect 270886 701190 270938 701242
rect 270950 701190 271002 701242
rect 271014 701190 271066 701242
rect 271078 701190 271130 701242
rect 271142 701190 271194 701242
rect 271206 701190 271258 701242
rect 271270 701190 271322 701242
rect 271334 701190 271386 701242
rect 306822 701190 306874 701242
rect 306886 701190 306938 701242
rect 306950 701190 307002 701242
rect 307014 701190 307066 701242
rect 307078 701190 307130 701242
rect 307142 701190 307194 701242
rect 307206 701190 307258 701242
rect 307270 701190 307322 701242
rect 307334 701190 307386 701242
rect 342822 701190 342874 701242
rect 342886 701190 342938 701242
rect 342950 701190 343002 701242
rect 343014 701190 343066 701242
rect 343078 701190 343130 701242
rect 343142 701190 343194 701242
rect 343206 701190 343258 701242
rect 343270 701190 343322 701242
rect 343334 701190 343386 701242
rect 378822 701190 378874 701242
rect 378886 701190 378938 701242
rect 378950 701190 379002 701242
rect 379014 701190 379066 701242
rect 379078 701190 379130 701242
rect 379142 701190 379194 701242
rect 379206 701190 379258 701242
rect 379270 701190 379322 701242
rect 379334 701190 379386 701242
rect 414822 701190 414874 701242
rect 414886 701190 414938 701242
rect 414950 701190 415002 701242
rect 415014 701190 415066 701242
rect 415078 701190 415130 701242
rect 415142 701190 415194 701242
rect 415206 701190 415258 701242
rect 415270 701190 415322 701242
rect 415334 701190 415386 701242
rect 450822 701190 450874 701242
rect 450886 701190 450938 701242
rect 450950 701190 451002 701242
rect 451014 701190 451066 701242
rect 451078 701190 451130 701242
rect 451142 701190 451194 701242
rect 451206 701190 451258 701242
rect 451270 701190 451322 701242
rect 451334 701190 451386 701242
rect 486822 701190 486874 701242
rect 486886 701190 486938 701242
rect 486950 701190 487002 701242
rect 487014 701190 487066 701242
rect 487078 701190 487130 701242
rect 487142 701190 487194 701242
rect 487206 701190 487258 701242
rect 487270 701190 487322 701242
rect 487334 701190 487386 701242
rect 522822 701190 522874 701242
rect 522886 701190 522938 701242
rect 522950 701190 523002 701242
rect 523014 701190 523066 701242
rect 523078 701190 523130 701242
rect 523142 701190 523194 701242
rect 523206 701190 523258 701242
rect 523270 701190 523322 701242
rect 523334 701190 523386 701242
rect 558822 701190 558874 701242
rect 558886 701190 558938 701242
rect 558950 701190 559002 701242
rect 559014 701190 559066 701242
rect 559078 701190 559130 701242
rect 559142 701190 559194 701242
rect 559206 701190 559258 701242
rect 559270 701190 559322 701242
rect 559334 701190 559386 701242
rect 261116 700952 261168 701004
rect 413652 700952 413704 701004
rect 154120 700884 154172 700936
rect 317972 700884 318024 700936
rect 137836 700816 137888 700868
rect 313188 700816 313240 700868
rect 105452 700748 105504 700800
rect 322664 700748 322716 700800
rect 36822 700646 36874 700698
rect 36886 700646 36938 700698
rect 36950 700646 37002 700698
rect 37014 700646 37066 700698
rect 37078 700646 37130 700698
rect 37142 700646 37194 700698
rect 37206 700646 37258 700698
rect 37270 700646 37322 700698
rect 37334 700646 37386 700698
rect 72822 700646 72874 700698
rect 72886 700646 72938 700698
rect 72950 700646 73002 700698
rect 73014 700646 73066 700698
rect 73078 700646 73130 700698
rect 73142 700646 73194 700698
rect 73206 700646 73258 700698
rect 73270 700646 73322 700698
rect 73334 700646 73386 700698
rect 108822 700646 108874 700698
rect 108886 700646 108938 700698
rect 108950 700646 109002 700698
rect 109014 700646 109066 700698
rect 109078 700646 109130 700698
rect 109142 700646 109194 700698
rect 109206 700646 109258 700698
rect 109270 700646 109322 700698
rect 109334 700646 109386 700698
rect 144822 700646 144874 700698
rect 144886 700646 144938 700698
rect 144950 700646 145002 700698
rect 145014 700646 145066 700698
rect 145078 700646 145130 700698
rect 145142 700646 145194 700698
rect 145206 700646 145258 700698
rect 145270 700646 145322 700698
rect 145334 700646 145386 700698
rect 180822 700646 180874 700698
rect 180886 700646 180938 700698
rect 180950 700646 181002 700698
rect 181014 700646 181066 700698
rect 181078 700646 181130 700698
rect 181142 700646 181194 700698
rect 181206 700646 181258 700698
rect 181270 700646 181322 700698
rect 181334 700646 181386 700698
rect 216822 700646 216874 700698
rect 216886 700646 216938 700698
rect 216950 700646 217002 700698
rect 217014 700646 217066 700698
rect 217078 700646 217130 700698
rect 217142 700646 217194 700698
rect 217206 700646 217258 700698
rect 217270 700646 217322 700698
rect 217334 700646 217386 700698
rect 252822 700646 252874 700698
rect 252886 700646 252938 700698
rect 252950 700646 253002 700698
rect 253014 700646 253066 700698
rect 253078 700646 253130 700698
rect 253142 700646 253194 700698
rect 253206 700646 253258 700698
rect 253270 700646 253322 700698
rect 253334 700646 253386 700698
rect 288822 700646 288874 700698
rect 288886 700646 288938 700698
rect 288950 700646 289002 700698
rect 289014 700646 289066 700698
rect 289078 700646 289130 700698
rect 289142 700646 289194 700698
rect 289206 700646 289258 700698
rect 289270 700646 289322 700698
rect 289334 700646 289386 700698
rect 324822 700646 324874 700698
rect 324886 700646 324938 700698
rect 324950 700646 325002 700698
rect 325014 700646 325066 700698
rect 325078 700646 325130 700698
rect 325142 700646 325194 700698
rect 325206 700646 325258 700698
rect 325270 700646 325322 700698
rect 325334 700646 325386 700698
rect 360822 700646 360874 700698
rect 360886 700646 360938 700698
rect 360950 700646 361002 700698
rect 361014 700646 361066 700698
rect 361078 700646 361130 700698
rect 361142 700646 361194 700698
rect 361206 700646 361258 700698
rect 361270 700646 361322 700698
rect 361334 700646 361386 700698
rect 396822 700646 396874 700698
rect 396886 700646 396938 700698
rect 396950 700646 397002 700698
rect 397014 700646 397066 700698
rect 397078 700646 397130 700698
rect 397142 700646 397194 700698
rect 397206 700646 397258 700698
rect 397270 700646 397322 700698
rect 397334 700646 397386 700698
rect 432822 700646 432874 700698
rect 432886 700646 432938 700698
rect 432950 700646 433002 700698
rect 433014 700646 433066 700698
rect 433078 700646 433130 700698
rect 433142 700646 433194 700698
rect 433206 700646 433258 700698
rect 433270 700646 433322 700698
rect 433334 700646 433386 700698
rect 468822 700646 468874 700698
rect 468886 700646 468938 700698
rect 468950 700646 469002 700698
rect 469014 700646 469066 700698
rect 469078 700646 469130 700698
rect 469142 700646 469194 700698
rect 469206 700646 469258 700698
rect 469270 700646 469322 700698
rect 469334 700646 469386 700698
rect 504822 700646 504874 700698
rect 504886 700646 504938 700698
rect 504950 700646 505002 700698
rect 505014 700646 505066 700698
rect 505078 700646 505130 700698
rect 505142 700646 505194 700698
rect 505206 700646 505258 700698
rect 505270 700646 505322 700698
rect 505334 700646 505386 700698
rect 540822 700646 540874 700698
rect 540886 700646 540938 700698
rect 540950 700646 541002 700698
rect 541014 700646 541066 700698
rect 541078 700646 541130 700698
rect 541142 700646 541194 700698
rect 541206 700646 541258 700698
rect 541270 700646 541322 700698
rect 541334 700646 541386 700698
rect 576822 700646 576874 700698
rect 576886 700646 576938 700698
rect 576950 700646 577002 700698
rect 577014 700646 577066 700698
rect 577078 700646 577130 700698
rect 577142 700646 577194 700698
rect 577206 700646 577258 700698
rect 577270 700646 577322 700698
rect 577334 700646 577386 700698
rect 242256 700544 242308 700596
rect 462320 700544 462372 700596
rect 246948 700476 247000 700528
rect 478512 700476 478564 700528
rect 89168 700408 89220 700460
rect 332140 700408 332192 700460
rect 202788 700340 202840 700392
rect 296536 700340 296588 700392
rect 296628 700340 296680 700392
rect 543464 700340 543516 700392
rect 72700 700272 72752 700324
rect 327448 700272 327500 700324
rect 256424 700204 256476 700256
rect 397460 700204 397512 700256
rect 18822 700102 18874 700154
rect 18886 700102 18938 700154
rect 18950 700102 19002 700154
rect 19014 700102 19066 700154
rect 19078 700102 19130 700154
rect 19142 700102 19194 700154
rect 19206 700102 19258 700154
rect 19270 700102 19322 700154
rect 19334 700102 19386 700154
rect 54822 700102 54874 700154
rect 54886 700102 54938 700154
rect 54950 700102 55002 700154
rect 55014 700102 55066 700154
rect 55078 700102 55130 700154
rect 55142 700102 55194 700154
rect 55206 700102 55258 700154
rect 55270 700102 55322 700154
rect 55334 700102 55386 700154
rect 90822 700102 90874 700154
rect 90886 700102 90938 700154
rect 90950 700102 91002 700154
rect 91014 700102 91066 700154
rect 91078 700102 91130 700154
rect 91142 700102 91194 700154
rect 91206 700102 91258 700154
rect 91270 700102 91322 700154
rect 91334 700102 91386 700154
rect 126822 700102 126874 700154
rect 126886 700102 126938 700154
rect 126950 700102 127002 700154
rect 127014 700102 127066 700154
rect 127078 700102 127130 700154
rect 127142 700102 127194 700154
rect 127206 700102 127258 700154
rect 127270 700102 127322 700154
rect 127334 700102 127386 700154
rect 162822 700102 162874 700154
rect 162886 700102 162938 700154
rect 162950 700102 163002 700154
rect 163014 700102 163066 700154
rect 163078 700102 163130 700154
rect 163142 700102 163194 700154
rect 163206 700102 163258 700154
rect 163270 700102 163322 700154
rect 163334 700102 163386 700154
rect 198822 700102 198874 700154
rect 198886 700102 198938 700154
rect 198950 700102 199002 700154
rect 199014 700102 199066 700154
rect 199078 700102 199130 700154
rect 199142 700102 199194 700154
rect 199206 700102 199258 700154
rect 199270 700102 199322 700154
rect 199334 700102 199386 700154
rect 234822 700102 234874 700154
rect 234886 700102 234938 700154
rect 234950 700102 235002 700154
rect 235014 700102 235066 700154
rect 235078 700102 235130 700154
rect 235142 700102 235194 700154
rect 235206 700102 235258 700154
rect 235270 700102 235322 700154
rect 235334 700102 235386 700154
rect 270822 700102 270874 700154
rect 270886 700102 270938 700154
rect 270950 700102 271002 700154
rect 271014 700102 271066 700154
rect 271078 700102 271130 700154
rect 271142 700102 271194 700154
rect 271206 700102 271258 700154
rect 271270 700102 271322 700154
rect 271334 700102 271386 700154
rect 306822 700102 306874 700154
rect 306886 700102 306938 700154
rect 306950 700102 307002 700154
rect 307014 700102 307066 700154
rect 307078 700102 307130 700154
rect 307142 700102 307194 700154
rect 307206 700102 307258 700154
rect 307270 700102 307322 700154
rect 307334 700102 307386 700154
rect 342822 700102 342874 700154
rect 342886 700102 342938 700154
rect 342950 700102 343002 700154
rect 343014 700102 343066 700154
rect 343078 700102 343130 700154
rect 343142 700102 343194 700154
rect 343206 700102 343258 700154
rect 343270 700102 343322 700154
rect 343334 700102 343386 700154
rect 378822 700102 378874 700154
rect 378886 700102 378938 700154
rect 378950 700102 379002 700154
rect 379014 700102 379066 700154
rect 379078 700102 379130 700154
rect 379142 700102 379194 700154
rect 379206 700102 379258 700154
rect 379270 700102 379322 700154
rect 379334 700102 379386 700154
rect 414822 700102 414874 700154
rect 414886 700102 414938 700154
rect 414950 700102 415002 700154
rect 415014 700102 415066 700154
rect 415078 700102 415130 700154
rect 415142 700102 415194 700154
rect 415206 700102 415258 700154
rect 415270 700102 415322 700154
rect 415334 700102 415386 700154
rect 450822 700102 450874 700154
rect 450886 700102 450938 700154
rect 450950 700102 451002 700154
rect 451014 700102 451066 700154
rect 451078 700102 451130 700154
rect 451142 700102 451194 700154
rect 451206 700102 451258 700154
rect 451270 700102 451322 700154
rect 451334 700102 451386 700154
rect 486822 700102 486874 700154
rect 486886 700102 486938 700154
rect 486950 700102 487002 700154
rect 487014 700102 487066 700154
rect 487078 700102 487130 700154
rect 487142 700102 487194 700154
rect 487206 700102 487258 700154
rect 487270 700102 487322 700154
rect 487334 700102 487386 700154
rect 522822 700102 522874 700154
rect 522886 700102 522938 700154
rect 522950 700102 523002 700154
rect 523014 700102 523066 700154
rect 523078 700102 523130 700154
rect 523142 700102 523194 700154
rect 523206 700102 523258 700154
rect 523270 700102 523322 700154
rect 523334 700102 523386 700154
rect 558822 700102 558874 700154
rect 558886 700102 558938 700154
rect 558950 700102 559002 700154
rect 559014 700102 559066 700154
rect 559078 700102 559130 700154
rect 559142 700102 559194 700154
rect 559206 700102 559258 700154
rect 559270 700102 559322 700154
rect 559334 700102 559386 700154
rect 170312 700000 170364 700052
rect 308496 700000 308548 700052
rect 308588 700000 308640 700052
rect 265900 699932 265952 699984
rect 364984 699932 365036 699984
rect 218980 699864 219032 699916
rect 296720 699864 296772 699916
rect 298008 699864 298060 699916
rect 251088 699796 251140 699848
rect 267648 699796 267700 699848
rect 273260 699796 273312 699848
rect 331312 699864 331364 699916
rect 348792 699864 348844 699916
rect 259460 699728 259512 699780
rect 270592 699728 270644 699780
rect 332508 699796 332560 699848
rect 273904 699728 273956 699780
rect 283748 699728 283800 699780
rect 283840 699728 283892 699780
rect 288532 699728 288584 699780
rect 251088 699660 251140 699712
rect 282920 699660 282972 699712
rect 283012 699660 283064 699712
rect 296904 699728 296956 699780
rect 288716 699660 288768 699712
rect 292396 699660 292448 699712
rect 292488 699660 292540 699712
rect 302332 699660 302384 699712
rect 311992 699660 312044 699712
rect 36822 699558 36874 699610
rect 36886 699558 36938 699610
rect 36950 699558 37002 699610
rect 37014 699558 37066 699610
rect 37078 699558 37130 699610
rect 37142 699558 37194 699610
rect 37206 699558 37258 699610
rect 37270 699558 37322 699610
rect 37334 699558 37386 699610
rect 72822 699558 72874 699610
rect 72886 699558 72938 699610
rect 72950 699558 73002 699610
rect 73014 699558 73066 699610
rect 73078 699558 73130 699610
rect 73142 699558 73194 699610
rect 73206 699558 73258 699610
rect 73270 699558 73322 699610
rect 73334 699558 73386 699610
rect 108822 699558 108874 699610
rect 108886 699558 108938 699610
rect 108950 699558 109002 699610
rect 109014 699558 109066 699610
rect 109078 699558 109130 699610
rect 109142 699558 109194 699610
rect 109206 699558 109258 699610
rect 109270 699558 109322 699610
rect 109334 699558 109386 699610
rect 144822 699558 144874 699610
rect 144886 699558 144938 699610
rect 144950 699558 145002 699610
rect 145014 699558 145066 699610
rect 145078 699558 145130 699610
rect 145142 699558 145194 699610
rect 145206 699558 145258 699610
rect 145270 699558 145322 699610
rect 145334 699558 145386 699610
rect 180822 699558 180874 699610
rect 180886 699558 180938 699610
rect 180950 699558 181002 699610
rect 181014 699558 181066 699610
rect 181078 699558 181130 699610
rect 181142 699558 181194 699610
rect 181206 699558 181258 699610
rect 181270 699558 181322 699610
rect 181334 699558 181386 699610
rect 216822 699558 216874 699610
rect 216886 699558 216938 699610
rect 216950 699558 217002 699610
rect 217014 699558 217066 699610
rect 217078 699558 217130 699610
rect 217142 699558 217194 699610
rect 217206 699558 217258 699610
rect 217270 699558 217322 699610
rect 217334 699558 217386 699610
rect 252822 699558 252874 699610
rect 252886 699558 252938 699610
rect 252950 699558 253002 699610
rect 253014 699558 253066 699610
rect 253078 699558 253130 699610
rect 253142 699558 253194 699610
rect 253206 699558 253258 699610
rect 253270 699558 253322 699610
rect 253334 699558 253386 699610
rect 288822 699558 288874 699610
rect 288886 699558 288938 699610
rect 288950 699558 289002 699610
rect 289014 699558 289066 699610
rect 289078 699558 289130 699610
rect 289142 699558 289194 699610
rect 289206 699558 289258 699610
rect 289270 699558 289322 699610
rect 289334 699558 289386 699610
rect 324822 699558 324874 699610
rect 324886 699558 324938 699610
rect 324950 699558 325002 699610
rect 325014 699558 325066 699610
rect 325078 699558 325130 699610
rect 325142 699558 325194 699610
rect 325206 699558 325258 699610
rect 325270 699558 325322 699610
rect 325334 699558 325386 699610
rect 360822 699558 360874 699610
rect 360886 699558 360938 699610
rect 360950 699558 361002 699610
rect 361014 699558 361066 699610
rect 361078 699558 361130 699610
rect 361142 699558 361194 699610
rect 361206 699558 361258 699610
rect 361270 699558 361322 699610
rect 361334 699558 361386 699610
rect 396822 699558 396874 699610
rect 396886 699558 396938 699610
rect 396950 699558 397002 699610
rect 397014 699558 397066 699610
rect 397078 699558 397130 699610
rect 397142 699558 397194 699610
rect 397206 699558 397258 699610
rect 397270 699558 397322 699610
rect 397334 699558 397386 699610
rect 432822 699558 432874 699610
rect 432886 699558 432938 699610
rect 432950 699558 433002 699610
rect 433014 699558 433066 699610
rect 433078 699558 433130 699610
rect 433142 699558 433194 699610
rect 433206 699558 433258 699610
rect 433270 699558 433322 699610
rect 433334 699558 433386 699610
rect 468822 699558 468874 699610
rect 468886 699558 468938 699610
rect 468950 699558 469002 699610
rect 469014 699558 469066 699610
rect 469078 699558 469130 699610
rect 469142 699558 469194 699610
rect 469206 699558 469258 699610
rect 469270 699558 469322 699610
rect 469334 699558 469386 699610
rect 504822 699558 504874 699610
rect 504886 699558 504938 699610
rect 504950 699558 505002 699610
rect 505014 699558 505066 699610
rect 505078 699558 505130 699610
rect 505142 699558 505194 699610
rect 505206 699558 505258 699610
rect 505270 699558 505322 699610
rect 505334 699558 505386 699610
rect 540822 699558 540874 699610
rect 540886 699558 540938 699610
rect 540950 699558 541002 699610
rect 541014 699558 541066 699610
rect 541078 699558 541130 699610
rect 541142 699558 541194 699610
rect 541206 699558 541258 699610
rect 541270 699558 541322 699610
rect 541334 699558 541386 699610
rect 576822 699558 576874 699610
rect 576886 699558 576938 699610
rect 576950 699558 577002 699610
rect 577014 699558 577066 699610
rect 577078 699558 577130 699610
rect 577142 699558 577194 699610
rect 577206 699558 577258 699610
rect 577270 699558 577322 699610
rect 577334 699558 577386 699610
rect 142804 699456 142856 699508
rect 403348 699456 403400 699508
rect 71780 699388 71832 699440
rect 417332 699388 417384 699440
rect 100208 699320 100260 699372
rect 273352 699320 273404 699372
rect 283012 699320 283064 699372
rect 296536 699320 296588 699372
rect 296628 699320 296680 699372
rect 445760 699320 445812 699372
rect 133328 699252 133380 699304
rect 146944 699252 146996 699304
rect 161756 699252 161808 699304
rect 579344 699252 579396 699304
rect 48136 699184 48188 699236
rect 142712 699184 142764 699236
rect 147588 699184 147640 699236
rect 186136 699184 186188 699236
rect 267648 699184 267700 699236
rect 302332 699184 302384 699236
rect 5080 699116 5132 699168
rect 311716 699184 311768 699236
rect 364340 699184 364392 699236
rect 373908 699184 373960 699236
rect 374000 699184 374052 699236
rect 383568 699184 383620 699236
rect 579252 699184 579304 699236
rect 321652 699116 321704 699168
rect 331036 699116 331088 699168
rect 331128 699116 331180 699168
rect 340696 699116 340748 699168
rect 459928 699116 459980 699168
rect 18822 699014 18874 699066
rect 18886 699014 18938 699066
rect 18950 699014 19002 699066
rect 19014 699014 19066 699066
rect 19078 699014 19130 699066
rect 19142 699014 19194 699066
rect 19206 699014 19258 699066
rect 19270 699014 19322 699066
rect 19334 699014 19386 699066
rect 54822 699014 54874 699066
rect 54886 699014 54938 699066
rect 54950 699014 55002 699066
rect 55014 699014 55066 699066
rect 55078 699014 55130 699066
rect 55142 699014 55194 699066
rect 55206 699014 55258 699066
rect 55270 699014 55322 699066
rect 55334 699014 55386 699066
rect 90822 699014 90874 699066
rect 90886 699014 90938 699066
rect 90950 699014 91002 699066
rect 91014 699014 91066 699066
rect 91078 699014 91130 699066
rect 91142 699014 91194 699066
rect 91206 699014 91258 699066
rect 91270 699014 91322 699066
rect 91334 699014 91386 699066
rect 126822 699014 126874 699066
rect 126886 699014 126938 699066
rect 126950 699014 127002 699066
rect 127014 699014 127066 699066
rect 127078 699014 127130 699066
rect 127142 699014 127194 699066
rect 127206 699014 127258 699066
rect 127270 699014 127322 699066
rect 127334 699014 127386 699066
rect 162822 699014 162874 699066
rect 162886 699014 162938 699066
rect 162950 699014 163002 699066
rect 163014 699014 163066 699066
rect 163078 699014 163130 699066
rect 163142 699014 163194 699066
rect 163206 699014 163258 699066
rect 163270 699014 163322 699066
rect 163334 699014 163386 699066
rect 198822 699014 198874 699066
rect 198886 699014 198938 699066
rect 198950 699014 199002 699066
rect 199014 699014 199066 699066
rect 199078 699014 199130 699066
rect 199142 699014 199194 699066
rect 199206 699014 199258 699066
rect 199270 699014 199322 699066
rect 199334 699014 199386 699066
rect 234822 699014 234874 699066
rect 234886 699014 234938 699066
rect 234950 699014 235002 699066
rect 235014 699014 235066 699066
rect 235078 699014 235130 699066
rect 235142 699014 235194 699066
rect 235206 699014 235258 699066
rect 235270 699014 235322 699066
rect 235334 699014 235386 699066
rect 270822 699014 270874 699066
rect 270886 699014 270938 699066
rect 270950 699014 271002 699066
rect 271014 699014 271066 699066
rect 271078 699014 271130 699066
rect 271142 699014 271194 699066
rect 271206 699014 271258 699066
rect 271270 699014 271322 699066
rect 271334 699014 271386 699066
rect 306822 699014 306874 699066
rect 306886 699014 306938 699066
rect 306950 699014 307002 699066
rect 307014 699014 307066 699066
rect 307078 699014 307130 699066
rect 307142 699014 307194 699066
rect 307206 699014 307258 699066
rect 307270 699014 307322 699066
rect 307334 699014 307386 699066
rect 342822 699014 342874 699066
rect 342886 699014 342938 699066
rect 342950 699014 343002 699066
rect 343014 699014 343066 699066
rect 343078 699014 343130 699066
rect 343142 699014 343194 699066
rect 343206 699014 343258 699066
rect 343270 699014 343322 699066
rect 343334 699014 343386 699066
rect 378822 699014 378874 699066
rect 378886 699014 378938 699066
rect 378950 699014 379002 699066
rect 379014 699014 379066 699066
rect 379078 699014 379130 699066
rect 379142 699014 379194 699066
rect 379206 699014 379258 699066
rect 379270 699014 379322 699066
rect 379334 699014 379386 699066
rect 414822 699014 414874 699066
rect 414886 699014 414938 699066
rect 414950 699014 415002 699066
rect 415014 699014 415066 699066
rect 415078 699014 415130 699066
rect 415142 699014 415194 699066
rect 415206 699014 415258 699066
rect 415270 699014 415322 699066
rect 415334 699014 415386 699066
rect 450822 699014 450874 699066
rect 450886 699014 450938 699066
rect 450950 699014 451002 699066
rect 451014 699014 451066 699066
rect 451078 699014 451130 699066
rect 451142 699014 451194 699066
rect 451206 699014 451258 699066
rect 451270 699014 451322 699066
rect 451334 699014 451386 699066
rect 486822 699014 486874 699066
rect 486886 699014 486938 699066
rect 486950 699014 487002 699066
rect 487014 699014 487066 699066
rect 487078 699014 487130 699066
rect 487142 699014 487194 699066
rect 487206 699014 487258 699066
rect 487270 699014 487322 699066
rect 487334 699014 487386 699066
rect 522822 699014 522874 699066
rect 522886 699014 522938 699066
rect 522950 699014 523002 699066
rect 523014 699014 523066 699066
rect 523078 699014 523130 699066
rect 523142 699014 523194 699066
rect 523206 699014 523258 699066
rect 523270 699014 523322 699066
rect 523334 699014 523386 699066
rect 558822 699014 558874 699066
rect 558886 699014 558938 699066
rect 558950 699014 559002 699066
rect 559014 699014 559066 699066
rect 559078 699014 559130 699066
rect 559142 699014 559194 699066
rect 559206 699014 559258 699066
rect 559270 699014 559322 699066
rect 559334 699014 559386 699066
rect 119160 698912 119212 698964
rect 244096 698912 244148 698964
rect 244188 698912 244240 698964
rect 244280 698912 244332 698964
rect 244372 698912 244424 698964
rect 253756 698912 253808 698964
rect 253848 698912 253900 698964
rect 282920 698912 282972 698964
rect 321560 698912 321612 698964
rect 321652 698912 321704 698964
rect 344928 698912 344980 698964
rect 579160 698912 579212 698964
rect 57612 698844 57664 698896
rect 107568 698844 107620 698896
rect 114376 698844 114428 698896
rect 577780 698844 577832 698896
rect 5264 698776 5316 698828
rect 474188 698776 474240 698828
rect 33968 698708 34020 698760
rect 89720 698708 89772 698760
rect 104992 698708 105044 698760
rect 579068 698708 579120 698760
rect 90732 698640 90784 698692
rect 578976 698640 579028 698692
rect 5356 698572 5408 698624
rect 502524 698572 502576 698624
rect 36822 698470 36874 698522
rect 36886 698470 36938 698522
rect 36950 698470 37002 698522
rect 37014 698470 37066 698522
rect 37078 698470 37130 698522
rect 37142 698470 37194 698522
rect 37206 698470 37258 698522
rect 37270 698470 37322 698522
rect 37334 698470 37386 698522
rect 72822 698470 72874 698522
rect 72886 698470 72938 698522
rect 72950 698470 73002 698522
rect 73014 698470 73066 698522
rect 73078 698470 73130 698522
rect 73142 698470 73194 698522
rect 73206 698470 73258 698522
rect 73270 698470 73322 698522
rect 73334 698470 73386 698522
rect 108822 698470 108874 698522
rect 108886 698470 108938 698522
rect 108950 698470 109002 698522
rect 109014 698470 109066 698522
rect 109078 698470 109130 698522
rect 109142 698470 109194 698522
rect 109206 698470 109258 698522
rect 109270 698470 109322 698522
rect 109334 698470 109386 698522
rect 144822 698470 144874 698522
rect 144886 698470 144938 698522
rect 144950 698470 145002 698522
rect 145014 698470 145066 698522
rect 145078 698470 145130 698522
rect 145142 698470 145194 698522
rect 145206 698470 145258 698522
rect 145270 698470 145322 698522
rect 145334 698470 145386 698522
rect 180822 698470 180874 698522
rect 180886 698470 180938 698522
rect 180950 698470 181002 698522
rect 181014 698470 181066 698522
rect 181078 698470 181130 698522
rect 181142 698470 181194 698522
rect 181206 698470 181258 698522
rect 181270 698470 181322 698522
rect 181334 698470 181386 698522
rect 216822 698470 216874 698522
rect 216886 698470 216938 698522
rect 216950 698470 217002 698522
rect 217014 698470 217066 698522
rect 217078 698470 217130 698522
rect 217142 698470 217194 698522
rect 217206 698470 217258 698522
rect 217270 698470 217322 698522
rect 217334 698470 217386 698522
rect 252822 698470 252874 698522
rect 252886 698470 252938 698522
rect 252950 698470 253002 698522
rect 253014 698470 253066 698522
rect 253078 698470 253130 698522
rect 253142 698470 253194 698522
rect 253206 698470 253258 698522
rect 253270 698470 253322 698522
rect 253334 698470 253386 698522
rect 288822 698470 288874 698522
rect 288886 698470 288938 698522
rect 288950 698470 289002 698522
rect 289014 698470 289066 698522
rect 289078 698470 289130 698522
rect 289142 698470 289194 698522
rect 289206 698470 289258 698522
rect 289270 698470 289322 698522
rect 289334 698470 289386 698522
rect 324822 698470 324874 698522
rect 324886 698470 324938 698522
rect 324950 698470 325002 698522
rect 325014 698470 325066 698522
rect 325078 698470 325130 698522
rect 325142 698470 325194 698522
rect 325206 698470 325258 698522
rect 325270 698470 325322 698522
rect 325334 698470 325386 698522
rect 360822 698470 360874 698522
rect 360886 698470 360938 698522
rect 360950 698470 361002 698522
rect 361014 698470 361066 698522
rect 361078 698470 361130 698522
rect 361142 698470 361194 698522
rect 361206 698470 361258 698522
rect 361270 698470 361322 698522
rect 361334 698470 361386 698522
rect 396822 698470 396874 698522
rect 396886 698470 396938 698522
rect 396950 698470 397002 698522
rect 397014 698470 397066 698522
rect 397078 698470 397130 698522
rect 397142 698470 397194 698522
rect 397206 698470 397258 698522
rect 397270 698470 397322 698522
rect 397334 698470 397386 698522
rect 432822 698470 432874 698522
rect 432886 698470 432938 698522
rect 432950 698470 433002 698522
rect 433014 698470 433066 698522
rect 433078 698470 433130 698522
rect 433142 698470 433194 698522
rect 433206 698470 433258 698522
rect 433270 698470 433322 698522
rect 433334 698470 433386 698522
rect 468822 698470 468874 698522
rect 468886 698470 468938 698522
rect 468950 698470 469002 698522
rect 469014 698470 469066 698522
rect 469078 698470 469130 698522
rect 469142 698470 469194 698522
rect 469206 698470 469258 698522
rect 469270 698470 469322 698522
rect 469334 698470 469386 698522
rect 504822 698470 504874 698522
rect 504886 698470 504938 698522
rect 504950 698470 505002 698522
rect 505014 698470 505066 698522
rect 505078 698470 505130 698522
rect 505142 698470 505194 698522
rect 505206 698470 505258 698522
rect 505270 698470 505322 698522
rect 505334 698470 505386 698522
rect 540822 698470 540874 698522
rect 540886 698470 540938 698522
rect 540950 698470 541002 698522
rect 541014 698470 541066 698522
rect 541078 698470 541130 698522
rect 541142 698470 541194 698522
rect 541206 698470 541258 698522
rect 541270 698470 541322 698522
rect 541334 698470 541386 698522
rect 576822 698470 576874 698522
rect 576886 698470 576938 698522
rect 576950 698470 577002 698522
rect 577014 698470 577066 698522
rect 577078 698470 577130 698522
rect 577142 698470 577194 698522
rect 577206 698470 577258 698522
rect 577270 698470 577322 698522
rect 577334 698470 577386 698522
rect 76564 698368 76616 698420
rect 218060 698368 218112 698420
rect 218428 698368 218480 698420
rect 578884 698368 578936 698420
rect 62304 698300 62356 698352
rect 577596 698300 577648 698352
rect 5816 698232 5868 698284
rect 218060 698232 218112 698284
rect 218428 698232 218480 698284
rect 5908 698164 5960 698216
rect 215116 698207 215168 698216
rect 215116 698173 215125 698207
rect 215125 698173 215159 698207
rect 215159 698173 215168 698207
rect 215116 698164 215168 698173
rect 218152 698164 218204 698216
rect 218336 698164 218388 698216
rect 226340 698164 226392 698216
rect 235908 698164 235960 698216
rect 237380 698164 237432 698216
rect 237564 698164 237616 698216
rect 253848 698164 253900 698216
rect 254032 698164 254084 698216
rect 350448 698164 350500 698216
rect 350724 698232 350776 698284
rect 365260 698232 365312 698284
rect 393964 698232 394016 698284
rect 351092 698164 351144 698216
rect 580540 698164 580592 698216
rect 193312 698139 193364 698148
rect 193312 698105 193321 698139
rect 193321 698105 193355 698139
rect 193355 698105 193364 698139
rect 193312 698096 193364 698105
rect 202788 698096 202840 698148
rect 208952 698096 209004 698148
rect 209044 698096 209096 698148
rect 576032 698096 576084 698148
rect 213828 698028 213880 698080
rect 579620 698028 579672 698080
rect 6092 697960 6144 698012
rect 379520 697960 379572 698012
rect 194876 697892 194928 697944
rect 574652 697892 574704 697944
rect 6092 697824 6144 697876
rect 393688 697824 393740 697876
rect 393964 697824 394016 697876
rect 580632 697824 580684 697876
rect 7472 697756 7524 697808
rect 398380 697756 398432 697808
rect 180708 697688 180760 697740
rect 575388 697688 575440 697740
rect 6828 697620 6880 697672
rect 407856 697620 407908 697672
rect 166448 697552 166500 697604
rect 575296 697552 575348 697604
rect 6736 697484 6788 697536
rect 422116 697484 422168 697536
rect 152280 697416 152332 697468
rect 575204 697416 575256 697468
rect 6552 697348 6604 697400
rect 436284 697348 436336 697400
rect 6368 697280 6420 697332
rect 455236 697280 455288 697332
rect 6276 697212 6328 697264
rect 464712 697212 464764 697264
rect 7932 697144 7984 697196
rect 493048 697144 493100 697196
rect 7564 697076 7616 697128
rect 535644 697076 535696 697128
rect 38660 697008 38712 697060
rect 574928 697008 574980 697060
rect 24492 696940 24544 696992
rect 574836 696940 574888 696992
rect 232964 696872 233016 696924
rect 233056 696872 233108 696924
rect 248328 696872 248380 696924
rect 248420 696872 248472 696924
rect 284484 696872 284536 696924
rect 289728 696804 289780 696856
rect 309140 696804 309192 696856
rect 4068 696668 4120 696720
rect 5448 696600 5500 696652
rect 160100 696736 160152 696788
rect 160192 696736 160244 696788
rect 234528 696736 234580 696788
rect 244280 696736 244332 696788
rect 299480 696736 299532 696788
rect 309048 696736 309100 696788
rect 321560 696736 321612 696788
rect 328460 696736 328512 696788
rect 342628 696736 342680 696788
rect 360200 696872 360252 696924
rect 388996 696736 389048 696788
rect 218520 696668 218572 696720
rect 578700 696668 578752 696720
rect 146944 696600 146996 696652
rect 580724 696600 580776 696652
rect 142712 696532 142764 696584
rect 580356 696532 580408 696584
rect 3148 696464 3200 696516
rect 374736 696464 374788 696516
rect 403348 696464 403400 696516
rect 580816 696464 580868 696516
rect 3884 696192 3936 696244
rect 165528 696396 165580 696448
rect 165712 696396 165764 696448
rect 204352 696396 204404 696448
rect 578792 696396 578844 696448
rect 224960 696328 225012 696380
rect 234528 696328 234580 696380
rect 244280 696328 244332 696380
rect 253848 696328 253900 696380
rect 263600 696328 263652 696380
rect 273168 696328 273220 696380
rect 282920 696328 282972 696380
rect 292488 696328 292540 696380
rect 190184 696260 190236 696312
rect 81256 696235 81308 696244
rect 81256 696201 81265 696235
rect 81265 696201 81299 696235
rect 81299 696201 81308 696235
rect 81256 696192 81308 696201
rect 107568 696192 107620 696244
rect 580448 696192 580500 696244
rect 3332 696124 3384 696176
rect 403164 696124 403216 696176
rect 579528 696124 579580 696176
rect 8208 696056 8260 696108
rect 412640 696056 412692 696108
rect 425152 696056 425204 696108
rect 426900 696056 426952 696108
rect 5172 695988 5224 696040
rect 431316 695988 431368 696040
rect 6460 695920 6512 695972
rect 450084 695920 450136 695972
rect 3792 695852 3844 695904
rect 469220 695852 469272 695904
rect 8024 695784 8076 695836
rect 478788 695784 478840 695836
rect 485780 695784 485832 695836
rect 492588 695784 492640 695836
rect 4896 695648 4948 695700
rect 487988 695716 488040 695768
rect 562324 695716 562376 695768
rect 567108 695716 567160 695768
rect 7748 695648 7800 695700
rect 506940 695648 506992 695700
rect 540980 695648 541032 695700
rect 543832 695648 543884 695700
rect 53288 695580 53340 695632
rect 575020 695580 575072 695632
rect 3516 695512 3568 695564
rect 530676 695512 530728 695564
rect 7288 695444 7340 695496
rect 355508 695444 355560 695496
rect 375380 695444 375432 695496
rect 384948 695444 385000 695496
rect 7380 695376 7432 695428
rect 369952 695376 370004 695428
rect 3240 695308 3292 695360
rect 383844 695308 383896 695360
rect 440700 695351 440752 695360
rect 440700 695317 440709 695351
rect 440709 695317 440743 695351
rect 440743 695317 440752 695351
rect 440700 695308 440752 695317
rect 483388 695351 483440 695360
rect 483388 695317 483397 695351
rect 483397 695317 483431 695351
rect 483431 695317 483440 695351
rect 483388 695308 483440 695317
rect 497556 695351 497608 695360
rect 497556 695317 497565 695351
rect 497565 695317 497599 695351
rect 497599 695317 497608 695351
rect 497556 695308 497608 695317
rect 511908 695351 511960 695360
rect 511908 695317 511917 695351
rect 511917 695317 511951 695351
rect 511951 695317 511960 695351
rect 511908 695308 511960 695317
rect 29552 695283 29604 695292
rect 29552 695249 29561 695283
rect 29561 695249 29595 695283
rect 29595 695249 29604 695283
rect 29552 695240 29604 695249
rect 43720 695283 43772 695292
rect 43720 695249 43729 695283
rect 43729 695249 43763 695283
rect 43763 695249 43772 695283
rect 43720 695240 43772 695249
rect 67456 695283 67508 695292
rect 67456 695249 67465 695283
rect 67465 695249 67499 695283
rect 67499 695249 67508 695283
rect 67456 695240 67508 695249
rect 86408 695283 86460 695292
rect 86408 695249 86417 695283
rect 86417 695249 86451 695283
rect 86451 695249 86460 695283
rect 86408 695240 86460 695249
rect 95792 695283 95844 695292
rect 95792 695249 95801 695283
rect 95801 695249 95835 695283
rect 95835 695249 95844 695283
rect 95792 695240 95844 695249
rect 109960 695283 110012 695292
rect 109960 695249 109969 695283
rect 109969 695249 110003 695283
rect 110003 695249 110012 695283
rect 109960 695240 110012 695249
rect 124128 695283 124180 695292
rect 124128 695249 124137 695283
rect 124137 695249 124171 695283
rect 124171 695249 124180 695283
rect 124128 695240 124180 695249
rect 128912 695283 128964 695292
rect 128912 695249 128921 695283
rect 128921 695249 128955 695283
rect 128955 695249 128964 695283
rect 128912 695240 128964 695249
rect 138480 695283 138532 695292
rect 138480 695249 138489 695283
rect 138489 695249 138523 695283
rect 138523 695249 138532 695283
rect 138480 695240 138532 695249
rect 171600 695240 171652 695292
rect 185768 695240 185820 695292
rect 199936 695240 199988 695292
rect 577412 695240 577464 695292
rect 578148 695308 578200 695360
rect 578056 695104 578108 695156
rect 3976 695036 4028 695088
rect 8116 695036 8168 695088
rect 576768 694968 576820 695020
rect 577872 694900 577924 694952
rect 576676 694832 576728 694884
rect 576584 694764 576636 694816
rect 569316 694696 569368 694748
rect 577504 694696 577556 694748
rect 3700 694560 3752 694612
rect 576492 694628 576544 694680
rect 7840 694560 7892 694612
rect 577688 694492 577740 694544
rect 576400 694424 576452 694476
rect 575112 694356 575164 694408
rect 3608 694288 3660 694340
rect 576308 694220 576360 694272
rect 576216 694152 576268 694204
rect 578700 687148 578752 687200
rect 580908 687148 580960 687200
rect 2964 682524 3016 682576
rect 5816 682524 5868 682576
rect 576032 674772 576084 674824
rect 579804 674772 579856 674824
rect 2780 668176 2832 668228
rect 5448 668176 5500 668228
rect 3056 653964 3108 654016
rect 7288 653964 7340 654016
rect 577412 651312 577464 651364
rect 579620 651312 579672 651364
rect 578792 640160 578844 640212
rect 580908 640160 580960 640212
rect 575480 627852 575532 627904
rect 579804 627852 579856 627904
rect 2964 624860 3016 624912
rect 5908 624860 5960 624912
rect 578148 604256 578200 604308
rect 579620 604256 579672 604308
rect 3148 596028 3200 596080
rect 7380 596028 7432 596080
rect 575388 580864 575440 580916
rect 580172 580864 580224 580916
rect 3056 567604 3108 567656
rect 6000 567604 6052 567656
rect 578056 557336 578108 557388
rect 579620 557336 579672 557388
rect 3884 539384 3936 539436
rect 5356 539384 5408 539436
rect 575296 534012 575348 534064
rect 579804 534012 579856 534064
rect 577964 510552 578016 510604
rect 580080 510552 580132 510604
rect 3056 510348 3108 510400
rect 6092 510348 6144 510400
rect 575204 487092 575256 487144
rect 580172 487092 580224 487144
rect 3332 481108 3384 481160
rect 7472 481108 7524 481160
rect 3332 452412 3384 452464
rect 6828 452412 6880 452464
rect 576768 440172 576820 440224
rect 579988 440172 580040 440224
rect 3332 438880 3384 438932
rect 5264 438880 5316 438932
rect 2872 423852 2924 423904
rect 8208 423852 8260 423904
rect 577872 416576 577924 416628
rect 579620 416576 579672 416628
rect 3240 395700 3292 395752
rect 6736 395700 6788 395752
rect 576676 393184 576728 393236
rect 579620 393184 579672 393236
rect 2780 380604 2832 380656
rect 5172 380604 5224 380656
rect 577780 369792 577832 369844
rect 580724 369792 580776 369844
rect 3240 367004 3292 367056
rect 6644 367004 6696 367056
rect 576584 346332 576636 346384
rect 580172 346332 580224 346384
rect 3240 337628 3292 337680
rect 6552 337628 6604 337680
rect 3240 308864 3292 308916
rect 8116 308864 8168 308916
rect 576492 299412 576544 299464
rect 580172 299412 580224 299464
rect 3240 294720 3292 294772
rect 6460 294720 6512 294772
rect 2780 280032 2832 280084
rect 5080 280032 5132 280084
rect 577688 275952 577740 276004
rect 579620 275952 579672 276004
rect 2964 266296 3016 266348
rect 6368 266296 6420 266348
rect 3240 252492 3292 252544
rect 6276 252492 6328 252544
rect 576400 252492 576452 252544
rect 580172 252492 580224 252544
rect 3332 208156 3384 208208
rect 8024 208156 8076 208208
rect 575112 205504 575164 205556
rect 580172 205504 580224 205556
rect 2780 194420 2832 194472
rect 4896 194420 4948 194472
rect 577596 170620 577648 170672
rect 580632 170620 580684 170672
rect 3332 165044 3384 165096
rect 7932 165044 7984 165096
rect 575020 158652 575072 158704
rect 579620 158652 579672 158704
rect 3332 136348 3384 136400
rect 7840 136348 7892 136400
rect 576308 135192 576360 135244
rect 580172 135192 580224 135244
rect 3332 122136 3384 122188
rect 7748 122136 7800 122188
rect 574928 111732 574980 111784
rect 580172 111732 580224 111784
rect 2780 107992 2832 108044
rect 4988 107992 5040 108044
rect 576216 88272 576268 88324
rect 579896 88272 579948 88324
rect 3056 79840 3108 79892
rect 7656 79840 7708 79892
rect 574928 64812 574980 64864
rect 579804 64812 579856 64864
rect 576124 41216 576176 41268
rect 580172 41216 580224 41268
rect 3424 35776 3476 35828
rect 7564 35776 7616 35828
rect 577504 30268 577556 30320
rect 579620 30268 579672 30320
rect 2780 21836 2832 21888
rect 4804 21836 4856 21888
rect 575020 17824 575072 17876
rect 580172 17824 580224 17876
rect 3148 7148 3200 7200
rect 6184 7148 6236 7200
rect 378140 6808 378192 6860
rect 388260 6808 388312 6860
rect 399668 6808 399720 6860
rect 408500 6808 408552 6860
rect 423496 6808 423548 6860
rect 433892 6808 433944 6860
rect 451832 6808 451884 6860
rect 463332 6808 463384 6860
rect 473360 6808 473412 6860
rect 484400 6808 484452 6860
rect 485872 6808 485924 6860
rect 496820 6808 496872 6860
rect 499488 6808 499540 6860
rect 510436 6808 510488 6860
rect 514208 6808 514260 6860
rect 524512 6808 524564 6860
rect 373632 6740 373684 6792
rect 383568 6740 383620 6792
rect 383844 6740 383896 6792
rect 394240 6740 394292 6792
rect 400772 6740 400824 6792
rect 412088 6740 412140 6792
rect 415584 6740 415636 6792
rect 426532 6740 426584 6792
rect 426900 6740 426952 6792
rect 437480 6740 437532 6792
rect 441620 6740 441672 6792
rect 453120 6740 453172 6792
rect 462044 6740 462096 6792
rect 472900 6740 472952 6792
rect 479064 6740 479116 6792
rect 491116 6740 491168 6792
rect 498292 6740 498344 6792
rect 510528 6740 510580 6792
rect 515312 6740 515364 6792
rect 525800 6740 525852 6792
rect 371332 6672 371384 6724
rect 381176 6672 381228 6724
rect 384948 6672 385000 6724
rect 331680 6604 331732 6656
rect 333980 6604 334032 6656
rect 377036 6604 377088 6656
rect 387064 6604 387116 6656
rect 390560 6672 390612 6724
rect 401324 6672 401376 6724
rect 403072 6672 403124 6724
rect 414480 6672 414532 6724
rect 394056 6604 394108 6656
rect 396264 6604 396316 6656
rect 407304 6604 407356 6656
rect 419172 6672 419224 6724
rect 434812 6672 434864 6724
rect 445852 6672 445904 6724
rect 449532 6672 449584 6724
rect 459560 6672 459612 6724
rect 460940 6672 460992 6724
rect 472532 6672 472584 6724
rect 476764 6672 476816 6724
rect 487436 6672 487488 6724
rect 493784 6672 493836 6724
rect 503904 6672 503956 6724
rect 505100 6672 505152 6724
rect 521476 6672 521528 6724
rect 523224 6672 523276 6724
rect 540520 6672 540572 6724
rect 418988 6604 419040 6656
rect 429200 6604 429252 6656
rect 431408 6604 431460 6656
rect 442356 6604 442408 6656
rect 446128 6604 446180 6656
rect 456800 6604 456852 6656
rect 464252 6604 464304 6656
rect 474740 6604 474792 6656
rect 477868 6604 477920 6656
rect 488540 6604 488592 6656
rect 506204 6604 506256 6656
rect 520832 6604 520884 6656
rect 524420 6604 524472 6656
rect 536748 6604 536800 6656
rect 360016 6536 360068 6588
rect 369216 6536 369268 6588
rect 370228 6536 370280 6588
rect 379980 6536 380032 6588
rect 401968 6536 402020 6588
rect 413284 6536 413336 6588
rect 416688 6536 416740 6588
rect 426440 6536 426492 6588
rect 426532 6536 426584 6588
rect 427544 6536 427596 6588
rect 430304 6536 430356 6588
rect 439044 6536 439096 6588
rect 442724 6536 442776 6588
rect 453672 6536 453724 6588
rect 454132 6536 454184 6588
rect 464436 6536 464488 6588
rect 467656 6536 467708 6588
rect 477592 6536 477644 6588
rect 482468 6536 482520 6588
rect 497740 6536 497792 6588
rect 502800 6536 502852 6588
rect 519084 6536 519136 6588
rect 521016 6536 521068 6588
rect 535920 6536 535972 6588
rect 70676 6468 70728 6520
rect 75460 6468 75512 6520
rect 356612 6468 356664 6520
rect 365720 6468 365772 6520
rect 369032 6468 369084 6520
rect 378692 6468 378744 6520
rect 382648 6468 382700 6520
rect 392768 6468 392820 6520
rect 392860 6468 392912 6520
rect 403716 6468 403768 6520
rect 407580 6468 407632 6520
rect 362224 6400 362276 6452
rect 371608 6400 371660 6452
rect 374736 6400 374788 6452
rect 384672 6400 384724 6452
rect 387248 6400 387300 6452
rect 397828 6400 397880 6452
rect 398564 6400 398616 6452
rect 409696 6400 409748 6452
rect 412180 6468 412232 6520
rect 423588 6468 423640 6520
rect 424600 6468 424652 6520
rect 434536 6468 434588 6520
rect 437112 6468 437164 6520
rect 447140 6468 447192 6520
rect 457536 6468 457588 6520
rect 467840 6468 467892 6520
rect 472256 6468 472308 6520
rect 483296 6468 483348 6520
rect 484676 6468 484728 6520
rect 500132 6468 500184 6520
rect 503996 6468 504048 6520
rect 514760 6468 514812 6520
rect 517612 6468 517664 6520
rect 534540 6468 534592 6520
rect 417792 6400 417844 6452
rect 427820 6400 427872 6452
rect 435916 6400 435968 6452
rect 445760 6400 445812 6452
rect 448428 6400 448480 6452
rect 458180 6400 458232 6452
rect 466552 6400 466604 6452
rect 477500 6400 477552 6452
rect 481272 6400 481324 6452
rect 496544 6400 496596 6452
rect 497188 6400 497240 6452
rect 513196 6400 513248 6452
rect 93308 6332 93360 6384
rect 96988 6332 97040 6384
rect 272708 6332 272760 6384
rect 275100 6332 275152 6384
rect 284024 6332 284076 6384
rect 285680 6332 285732 6384
rect 319168 6332 319220 6384
rect 322480 6332 322532 6384
rect 328276 6332 328328 6384
rect 330576 6332 330628 6384
rect 340696 6332 340748 6384
rect 342720 6332 342772 6384
rect 347504 6332 347556 6384
rect 356152 6332 356204 6384
rect 361120 6332 361172 6384
rect 370412 6332 370464 6384
rect 379244 6332 379296 6384
rect 389088 6332 389140 6384
rect 391756 6332 391808 6384
rect 402520 6332 402572 6384
rect 406476 6332 406528 6384
rect 417976 6332 418028 6384
rect 421196 6332 421248 6384
rect 432696 6332 432748 6384
rect 438216 6332 438268 6384
rect 448612 6332 448664 6384
rect 450728 6332 450780 6384
rect 462228 6332 462280 6384
rect 468852 6332 468904 6384
rect 478972 6332 479024 6384
rect 483572 6332 483624 6384
rect 491484 6332 491536 6384
rect 507216 6332 507268 6384
rect 507400 6332 507452 6384
rect 523868 6332 523920 6384
rect 353208 6264 353260 6316
rect 362132 6264 362184 6316
rect 364524 6264 364576 6316
rect 367468 6264 367520 6316
rect 367928 6264 367980 6316
rect 377588 6264 377640 6316
rect 386052 6264 386104 6316
rect 396632 6264 396684 6316
rect 397368 6264 397420 6316
rect 408408 6264 408460 6316
rect 413192 6264 413244 6316
rect 424968 6264 425020 6316
rect 429108 6264 429160 6316
rect 438860 6264 438912 6316
rect 443920 6264 443972 6316
rect 454132 6264 454184 6316
rect 458640 6264 458692 6316
rect 469496 6264 469548 6316
rect 480168 6264 480220 6316
rect 490748 6264 490800 6316
rect 494888 6264 494940 6316
rect 510804 6264 510856 6316
rect 516416 6264 516468 6316
rect 533344 6264 533396 6316
rect 83832 6196 83884 6248
rect 87880 6196 87932 6248
rect 264796 6196 264848 6248
rect 266360 6196 266412 6248
rect 273812 6196 273864 6248
rect 276020 6196 276072 6248
rect 337292 6196 337344 6248
rect 339684 6196 339736 6248
rect 354312 6196 354364 6248
rect 363328 6196 363380 6248
rect 363420 6196 363472 6248
rect 372804 6196 372856 6248
rect 375840 6196 375892 6248
rect 385868 6196 385920 6248
rect 388352 6196 388404 6248
rect 399024 6196 399076 6248
rect 404176 6196 404228 6248
rect 414112 6196 414164 6248
rect 420092 6196 420144 6248
rect 430580 6196 430632 6248
rect 432512 6196 432564 6248
rect 443552 6196 443604 6248
rect 447324 6196 447376 6248
rect 458272 6196 458324 6248
rect 463148 6196 463200 6248
rect 474096 6196 474148 6248
rect 475660 6196 475712 6248
rect 484676 6196 484728 6248
rect 486976 6196 487028 6248
rect 502432 6196 502484 6248
rect 508504 6196 508556 6248
rect 525064 6196 525116 6248
rect 530032 6196 530084 6248
rect 541440 6196 541492 6248
rect 5540 6128 5592 6180
rect 10784 6128 10836 6180
rect 63592 6128 63644 6180
rect 68652 6128 68704 6180
rect 87328 6128 87380 6180
rect 91284 6128 91336 6180
rect 199016 6128 199068 6180
rect 200396 6128 200448 6180
rect 235264 6128 235316 6180
rect 238392 6128 238444 6180
rect 342996 6128 343048 6180
rect 345940 6128 345992 6180
rect 355416 6128 355468 6180
rect 364524 6128 364576 6180
rect 372436 6128 372488 6180
rect 382372 6128 382424 6180
rect 389456 6128 389508 6180
rect 400220 6128 400272 6180
rect 405372 6128 405424 6180
rect 416688 6128 416740 6180
rect 422392 6128 422444 6180
rect 245476 6060 245528 6112
rect 247040 6060 247092 6112
rect 254584 6060 254636 6112
rect 256700 6060 256752 6112
rect 290832 6060 290884 6112
rect 292580 6060 292632 6112
rect 293132 6060 293184 6112
rect 295432 6060 295484 6112
rect 302148 6060 302200 6112
rect 304264 6060 304316 6112
rect 314660 6060 314712 6112
rect 318248 6060 318300 6112
rect 332784 6060 332836 6112
rect 336280 6060 336332 6112
rect 393964 6060 394016 6112
rect 403808 6060 403860 6112
rect 414388 6060 414440 6112
rect 424324 6060 424376 6112
rect 428004 6128 428056 6180
rect 438952 6128 439004 6180
rect 452936 6128 452988 6180
rect 463700 6128 463752 6180
rect 474464 6128 474516 6180
rect 489184 6128 489236 6180
rect 489276 6128 489328 6180
rect 500592 6128 500644 6180
rect 501696 6128 501748 6180
rect 517888 6128 517940 6180
rect 522120 6128 522172 6180
rect 539324 6128 539376 6180
rect 434628 6060 434680 6112
rect 439320 6060 439372 6112
rect 448520 6060 448572 6112
rect 455236 6060 455288 6112
rect 464252 6060 464304 6112
rect 465448 6060 465500 6112
rect 476120 6060 476172 6112
rect 494152 6060 494204 6112
rect 496084 6060 496136 6112
rect 506480 6060 506532 6112
rect 509608 6060 509660 6112
rect 521200 6060 521252 6112
rect 549352 6060 549404 6112
rect 550548 6060 550600 6112
rect 18822 5958 18874 6010
rect 18886 5958 18938 6010
rect 18950 5958 19002 6010
rect 19014 5958 19066 6010
rect 19078 5958 19130 6010
rect 19142 5958 19194 6010
rect 19206 5958 19258 6010
rect 19270 5958 19322 6010
rect 19334 5958 19386 6010
rect 54822 5958 54874 6010
rect 54886 5958 54938 6010
rect 54950 5958 55002 6010
rect 55014 5958 55066 6010
rect 55078 5958 55130 6010
rect 55142 5958 55194 6010
rect 55206 5958 55258 6010
rect 55270 5958 55322 6010
rect 55334 5958 55386 6010
rect 90822 5958 90874 6010
rect 90886 5958 90938 6010
rect 90950 5958 91002 6010
rect 91014 5958 91066 6010
rect 91078 5958 91130 6010
rect 91142 5958 91194 6010
rect 91206 5958 91258 6010
rect 91270 5958 91322 6010
rect 91334 5958 91386 6010
rect 126822 5958 126874 6010
rect 126886 5958 126938 6010
rect 126950 5958 127002 6010
rect 127014 5958 127066 6010
rect 127078 5958 127130 6010
rect 127142 5958 127194 6010
rect 127206 5958 127258 6010
rect 127270 5958 127322 6010
rect 127334 5958 127386 6010
rect 162822 5958 162874 6010
rect 162886 5958 162938 6010
rect 162950 5958 163002 6010
rect 163014 5958 163066 6010
rect 163078 5958 163130 6010
rect 163142 5958 163194 6010
rect 163206 5958 163258 6010
rect 163270 5958 163322 6010
rect 163334 5958 163386 6010
rect 198822 5958 198874 6010
rect 198886 5958 198938 6010
rect 198950 5958 199002 6010
rect 199014 5958 199066 6010
rect 199078 5958 199130 6010
rect 199142 5958 199194 6010
rect 199206 5958 199258 6010
rect 199270 5958 199322 6010
rect 199334 5958 199386 6010
rect 234822 5958 234874 6010
rect 234886 5958 234938 6010
rect 234950 5958 235002 6010
rect 235014 5958 235066 6010
rect 235078 5958 235130 6010
rect 235142 5958 235194 6010
rect 235206 5958 235258 6010
rect 235270 5958 235322 6010
rect 235334 5958 235386 6010
rect 270822 5958 270874 6010
rect 270886 5958 270938 6010
rect 270950 5958 271002 6010
rect 271014 5958 271066 6010
rect 271078 5958 271130 6010
rect 271142 5958 271194 6010
rect 271206 5958 271258 6010
rect 271270 5958 271322 6010
rect 271334 5958 271386 6010
rect 306822 5958 306874 6010
rect 306886 5958 306938 6010
rect 306950 5958 307002 6010
rect 307014 5958 307066 6010
rect 307078 5958 307130 6010
rect 307142 5958 307194 6010
rect 307206 5958 307258 6010
rect 307270 5958 307322 6010
rect 307334 5958 307386 6010
rect 342822 5958 342874 6010
rect 342886 5958 342938 6010
rect 342950 5958 343002 6010
rect 343014 5958 343066 6010
rect 343078 5958 343130 6010
rect 343142 5958 343194 6010
rect 343206 5958 343258 6010
rect 343270 5958 343322 6010
rect 343334 5958 343386 6010
rect 378822 5958 378874 6010
rect 378886 5958 378938 6010
rect 378950 5958 379002 6010
rect 379014 5958 379066 6010
rect 379078 5958 379130 6010
rect 379142 5958 379194 6010
rect 379206 5958 379258 6010
rect 379270 5958 379322 6010
rect 379334 5958 379386 6010
rect 414822 5958 414874 6010
rect 414886 5958 414938 6010
rect 414950 5958 415002 6010
rect 415014 5958 415066 6010
rect 415078 5958 415130 6010
rect 415142 5958 415194 6010
rect 415206 5958 415258 6010
rect 415270 5958 415322 6010
rect 415334 5958 415386 6010
rect 450822 5958 450874 6010
rect 450886 5958 450938 6010
rect 450950 5958 451002 6010
rect 451014 5958 451066 6010
rect 451078 5958 451130 6010
rect 451142 5958 451194 6010
rect 451206 5958 451258 6010
rect 451270 5958 451322 6010
rect 451334 5958 451386 6010
rect 486822 5958 486874 6010
rect 486886 5958 486938 6010
rect 486950 5958 487002 6010
rect 487014 5958 487066 6010
rect 487078 5958 487130 6010
rect 487142 5958 487194 6010
rect 487206 5958 487258 6010
rect 487270 5958 487322 6010
rect 487334 5958 487386 6010
rect 522822 5958 522874 6010
rect 522886 5958 522938 6010
rect 522950 5958 523002 6010
rect 523014 5958 523066 6010
rect 523078 5958 523130 6010
rect 523142 5958 523194 6010
rect 523206 5958 523258 6010
rect 523270 5958 523322 6010
rect 523334 5958 523386 6010
rect 558822 5958 558874 6010
rect 558886 5958 558938 6010
rect 558950 5958 559002 6010
rect 559014 5958 559066 6010
rect 559078 5958 559130 6010
rect 559142 5958 559194 6010
rect 559206 5958 559258 6010
rect 559270 5958 559322 6010
rect 559334 5958 559386 6010
rect 267004 5856 267056 5908
rect 269672 5856 269724 5908
rect 315764 5856 315816 5908
rect 318708 5856 318760 5908
rect 322572 5856 322624 5908
rect 324320 5856 324372 5908
rect 324872 5856 324924 5908
rect 328276 5856 328328 5908
rect 335084 5856 335136 5908
rect 337384 5856 337436 5908
rect 408776 5856 408828 5908
rect 418160 5856 418212 5908
rect 445024 5856 445076 5908
rect 454684 5856 454736 5908
rect 459744 5856 459796 5908
rect 469404 5856 469456 5908
rect 492680 5856 492732 5908
rect 503996 5856 504048 5908
rect 510712 5856 510764 5908
rect 522396 5856 522448 5908
rect 94504 5788 94556 5840
rect 98092 5788 98144 5840
rect 238668 5788 238720 5840
rect 240140 5788 240192 5840
rect 257988 5788 258040 5840
rect 260104 5788 260156 5840
rect 265900 5788 265952 5840
rect 269028 5788 269080 5840
rect 282920 5788 282972 5840
rect 285772 5788 285824 5840
rect 286324 5788 286376 5840
rect 289452 5788 289504 5840
rect 295340 5788 295392 5840
rect 298928 5788 298980 5840
rect 301044 5788 301096 5840
rect 303712 5788 303764 5840
rect 304448 5788 304500 5840
rect 307668 5788 307720 5840
rect 321468 5788 321520 5840
rect 323584 5788 323636 5840
rect 330484 5788 330536 5840
rect 332968 5788 333020 5840
rect 344100 5788 344152 5840
rect 347412 5788 347464 5840
rect 348700 5788 348752 5840
rect 351736 5788 351788 5840
rect 380440 5788 380492 5840
rect 382280 5788 382332 5840
rect 433708 5788 433760 5840
rect 444380 5788 444432 5840
rect 469956 5788 470008 5840
rect 478880 5788 478932 5840
rect 500500 5788 500552 5840
rect 511908 5788 511960 5840
rect 513012 5788 513064 5840
rect 529848 5788 529900 5840
rect 23848 5720 23900 5772
rect 25504 5720 25556 5772
rect 79048 5720 79100 5772
rect 83372 5720 83424 5772
rect 84936 5720 84988 5772
rect 88984 5720 89036 5772
rect 89720 5720 89772 5772
rect 93584 5720 93636 5772
rect 96896 5720 96948 5772
rect 100392 5720 100444 5772
rect 105176 5720 105228 5772
rect 108304 5720 108356 5772
rect 118240 5720 118292 5772
rect 120816 5720 120868 5772
rect 226248 5720 226300 5772
rect 228916 5720 228968 5772
rect 234160 5720 234212 5772
rect 237196 5720 237248 5772
rect 243176 5720 243228 5772
rect 246764 5720 246816 5772
rect 247776 5720 247828 5772
rect 251088 5720 251140 5772
rect 252284 5720 252336 5772
rect 254216 5720 254268 5772
rect 277216 5720 277268 5772
rect 279792 5720 279844 5772
rect 280620 5720 280672 5772
rect 283196 5720 283248 5772
rect 289728 5720 289780 5772
rect 292488 5720 292540 5772
rect 308956 5720 309008 5772
rect 311808 5720 311860 5772
rect 323676 5720 323728 5772
rect 326988 5720 327040 5772
rect 410984 5720 411036 5772
rect 413928 5720 413980 5772
rect 490380 5720 490432 5772
rect 506020 5720 506072 5772
rect 15200 5652 15252 5704
rect 17592 5652 17644 5704
rect 18604 5652 18656 5704
rect 20996 5652 21048 5704
rect 23112 5652 23164 5704
rect 24400 5652 24452 5704
rect 26240 5652 26292 5704
rect 28908 5652 28960 5704
rect 75460 5652 75512 5704
rect 79968 5652 80020 5704
rect 80244 5652 80296 5704
rect 84476 5652 84528 5704
rect 88524 5652 88576 5704
rect 92388 5652 92440 5704
rect 95700 5652 95752 5704
rect 99196 5652 99248 5704
rect 100484 5652 100536 5704
rect 103796 5652 103848 5704
rect 103980 5652 104032 5704
rect 107200 5652 107252 5704
rect 107568 5652 107620 5704
rect 110604 5652 110656 5704
rect 111156 5652 111208 5704
rect 114008 5652 114060 5704
rect 114744 5652 114796 5704
rect 117412 5652 117464 5704
rect 120632 5652 120684 5704
rect 123024 5652 123076 5704
rect 132592 5652 132644 5704
rect 134340 5652 134392 5704
rect 143264 5652 143316 5704
rect 144552 5652 144604 5704
rect 145656 5652 145708 5704
rect 146852 5652 146904 5704
rect 195612 5652 195664 5704
rect 196808 5652 196860 5704
rect 206928 5652 206980 5704
rect 208676 5652 208728 5704
rect 214840 5652 214892 5704
rect 216680 5652 216732 5704
rect 220544 5652 220596 5704
rect 222936 5652 222988 5704
rect 223948 5652 224000 5704
rect 226524 5652 226576 5704
rect 228456 5652 228508 5704
rect 231308 5652 231360 5704
rect 231860 5652 231912 5704
rect 234712 5652 234764 5704
rect 242072 5652 242124 5704
rect 245568 5652 245620 5704
rect 249984 5652 250036 5704
rect 253848 5652 253900 5704
rect 260196 5652 260248 5704
rect 262404 5652 262456 5704
rect 262496 5652 262548 5704
rect 264980 5652 265032 5704
rect 270408 5652 270460 5704
rect 272984 5652 273036 5704
rect 276112 5652 276164 5704
rect 279332 5652 279384 5704
rect 281724 5652 281776 5704
rect 284392 5652 284444 5704
rect 291936 5652 291988 5704
rect 294328 5652 294380 5704
rect 296536 5652 296588 5704
rect 299204 5652 299256 5704
rect 299940 5652 299992 5704
rect 303068 5652 303120 5704
rect 303344 5652 303396 5704
rect 305000 5652 305052 5704
rect 305552 5652 305604 5704
rect 308220 5652 308272 5704
rect 310152 5652 310204 5704
rect 313096 5652 313148 5704
rect 318064 5652 318116 5704
rect 321468 5652 321520 5704
rect 329380 5652 329432 5704
rect 332416 5652 332468 5704
rect 338488 5652 338540 5704
rect 341800 5652 341852 5704
rect 341892 5652 341944 5704
rect 343640 5652 343692 5704
rect 349804 5652 349856 5704
rect 352288 5652 352340 5704
rect 357716 5652 357768 5704
rect 360752 5652 360804 5704
rect 381544 5652 381596 5704
rect 384948 5652 385000 5704
rect 409880 5652 409932 5704
rect 413376 5652 413428 5704
rect 440516 5652 440568 5704
rect 444288 5652 444340 5704
rect 13820 5584 13872 5636
rect 16488 5584 16540 5636
rect 18052 5584 18104 5636
rect 19892 5584 19944 5636
rect 20720 5584 20772 5636
rect 23296 5584 23348 5636
rect 27712 5584 27764 5636
rect 30104 5584 30156 5636
rect 34520 5584 34572 5636
rect 36912 5584 36964 5636
rect 37464 5584 37516 5636
rect 39120 5584 39172 5636
rect 69480 5584 69532 5636
rect 74264 5584 74316 5636
rect 77852 5584 77904 5636
rect 82268 5584 82320 5636
rect 82636 5584 82688 5636
rect 86776 5584 86828 5636
rect 90732 5584 90784 5636
rect 94688 5584 94740 5636
rect 98092 5584 98144 5636
rect 101496 5584 101548 5636
rect 101588 5584 101640 5636
rect 104900 5584 104952 5636
rect 106372 5584 106424 5636
rect 109408 5584 109460 5636
rect 109960 5584 110012 5636
rect 112812 5584 112864 5636
rect 113548 5584 113600 5636
rect 116216 5584 116268 5636
rect 117136 5584 117188 5636
rect 119620 5584 119672 5636
rect 121828 5584 121880 5636
rect 124128 5584 124180 5636
rect 124220 5584 124272 5636
rect 126428 5584 126480 5636
rect 126612 5584 126664 5636
rect 128728 5584 128780 5636
rect 129004 5584 129056 5636
rect 130936 5584 130988 5636
rect 131396 5584 131448 5636
rect 133236 5584 133288 5636
rect 134892 5584 134944 5636
rect 136640 5584 136692 5636
rect 137284 5584 137336 5636
rect 138940 5584 138992 5636
rect 139676 5584 139728 5636
rect 141148 5584 141200 5636
rect 142068 5584 142120 5636
rect 143448 5584 143500 5636
rect 197912 5584 197964 5636
rect 198740 5584 198792 5636
rect 201224 5584 201276 5636
rect 202696 5584 202748 5636
rect 203524 5584 203576 5636
rect 205088 5584 205140 5636
rect 205824 5584 205876 5636
rect 207480 5584 207532 5636
rect 209228 5584 209280 5636
rect 211068 5584 211120 5636
rect 211436 5584 211488 5636
rect 213460 5584 213512 5636
rect 213736 5584 213788 5636
rect 215852 5584 215904 5636
rect 217140 5584 217192 5636
rect 219348 5584 219400 5636
rect 219440 5584 219492 5636
rect 221740 5584 221792 5636
rect 222844 5584 222896 5636
rect 225328 5584 225380 5636
rect 227352 5584 227404 5636
rect 230112 5584 230164 5636
rect 230756 5584 230808 5636
rect 233700 5584 233752 5636
rect 236368 5584 236420 5636
rect 239588 5584 239640 5636
rect 239772 5584 239824 5636
rect 242808 5584 242860 5636
rect 244372 5584 244424 5636
rect 247960 5584 248012 5636
rect 248880 5584 248932 5636
rect 252468 5584 252520 5636
rect 253388 5584 253440 5636
rect 255412 5584 255464 5636
rect 256792 5584 256844 5636
rect 260748 5584 260800 5636
rect 261392 5584 261444 5636
rect 263692 5584 263744 5636
rect 269304 5584 269356 5636
rect 271880 5584 271932 5636
rect 278320 5584 278372 5636
rect 280896 5584 280948 5636
rect 287428 5584 287480 5636
rect 290188 5584 290240 5636
rect 297640 5584 297692 5636
rect 300676 5584 300728 5636
rect 307852 5584 307904 5636
rect 311164 5584 311216 5636
rect 312360 5584 312412 5636
rect 314660 5584 314712 5636
rect 316868 5584 316920 5636
rect 320088 5584 320140 5636
rect 327080 5584 327132 5636
rect 330852 5584 330904 5636
rect 333888 5584 333940 5636
rect 336648 5584 336700 5636
rect 345296 5584 345348 5636
rect 348976 5584 349028 5636
rect 350908 5584 350960 5636
rect 353300 5584 353352 5636
rect 365628 5584 365680 5636
rect 367100 5584 367152 5636
rect 488080 5584 488132 5636
rect 491208 5584 491260 5636
rect 11060 5516 11112 5568
rect 14188 5516 14240 5568
rect 16948 5516 17000 5568
rect 18696 5516 18748 5568
rect 19432 5516 19484 5568
rect 22100 5516 22152 5568
rect 29000 5516 29052 5568
rect 31208 5516 31260 5568
rect 31760 5516 31812 5568
rect 33140 5516 33192 5568
rect 36452 5516 36504 5568
rect 38016 5516 38068 5568
rect 42800 5516 42852 5568
rect 44824 5516 44876 5568
rect 55404 5516 55456 5568
rect 60648 5516 60700 5568
rect 62396 5516 62448 5568
rect 67456 5516 67508 5568
rect 71872 5516 71924 5568
rect 76564 5516 76616 5568
rect 76656 5516 76708 5568
rect 81072 5516 81124 5568
rect 81440 5516 81492 5568
rect 85580 5516 85632 5568
rect 86132 5516 86184 5568
rect 90180 5516 90232 5568
rect 92112 5516 92164 5568
rect 95792 5516 95844 5568
rect 99288 5516 99340 5568
rect 102600 5516 102652 5568
rect 102784 5516 102836 5568
rect 106004 5516 106056 5568
rect 108672 5516 108724 5568
rect 111708 5516 111760 5568
rect 112352 5516 112404 5568
rect 115112 5516 115164 5568
rect 115940 5516 115992 5568
rect 118516 5516 118568 5568
rect 119436 5516 119488 5568
rect 121920 5516 121972 5568
rect 123024 5516 123076 5568
rect 125324 5516 125376 5568
rect 125416 5516 125468 5568
rect 127532 5516 127584 5568
rect 127808 5516 127860 5568
rect 129832 5516 129884 5568
rect 130200 5516 130252 5568
rect 132132 5516 132184 5568
rect 133788 5516 133840 5568
rect 135536 5516 135588 5568
rect 136088 5516 136140 5568
rect 137744 5516 137796 5568
rect 138480 5516 138532 5568
rect 140044 5516 140096 5568
rect 140872 5516 140924 5568
rect 142344 5516 142396 5568
rect 144460 5516 144512 5568
rect 145748 5516 145800 5568
rect 146852 5516 146904 5568
rect 147956 5516 148008 5568
rect 148048 5516 148100 5568
rect 149152 5516 149204 5568
rect 151544 5516 151596 5568
rect 152556 5516 152608 5568
rect 152740 5516 152792 5568
rect 153660 5516 153712 5568
rect 153936 5516 153988 5568
rect 154764 5516 154816 5568
rect 155132 5516 155184 5568
rect 155960 5516 156012 5568
rect 181996 5516 182048 5568
rect 182548 5516 182600 5568
rect 183100 5516 183152 5568
rect 183744 5516 183796 5568
rect 188804 5516 188856 5568
rect 189632 5516 189684 5568
rect 189908 5516 189960 5568
rect 190828 5516 190880 5568
rect 191104 5516 191156 5568
rect 192024 5516 192076 5568
rect 192208 5516 192260 5568
rect 193220 5516 193272 5568
rect 194508 5516 194560 5568
rect 195612 5516 195664 5568
rect 196716 5516 196768 5568
rect 198004 5516 198056 5568
rect 200120 5516 200172 5568
rect 201500 5516 201552 5568
rect 202420 5516 202472 5568
rect 203892 5516 203944 5568
rect 204628 5516 204680 5568
rect 206284 5516 206336 5568
rect 208032 5516 208084 5568
rect 209872 5516 209924 5568
rect 210332 5516 210384 5568
rect 212264 5516 212316 5568
rect 212632 5516 212684 5568
rect 214656 5516 214708 5568
rect 216036 5516 216088 5568
rect 218152 5516 218204 5568
rect 218244 5516 218296 5568
rect 220544 5516 220596 5568
rect 221648 5516 221700 5568
rect 224132 5516 224184 5568
rect 225052 5516 225104 5568
rect 227720 5516 227772 5568
rect 229652 5516 229704 5568
rect 232504 5516 232556 5568
rect 233056 5516 233108 5568
rect 235908 5516 235960 5568
rect 237564 5516 237616 5568
rect 240784 5516 240836 5568
rect 240968 5516 241020 5568
rect 244188 5516 244240 5568
rect 246580 5516 246632 5568
rect 249248 5516 249300 5568
rect 251180 5516 251232 5568
rect 255044 5516 255096 5568
rect 255688 5516 255740 5568
rect 259000 5516 259052 5568
rect 259092 5516 259144 5568
rect 261208 5516 261260 5568
rect 263600 5516 263652 5568
rect 266452 5516 266504 5568
rect 268200 5516 268252 5568
rect 270500 5516 270552 5568
rect 271604 5516 271656 5568
rect 273996 5516 274048 5568
rect 274916 5516 274968 5568
rect 278412 5516 278464 5568
rect 279516 5516 279568 5568
rect 282092 5516 282144 5568
rect 285128 5516 285180 5568
rect 288256 5516 288308 5568
rect 288532 5516 288584 5568
rect 291384 5516 291436 5568
rect 294236 5516 294288 5568
rect 297824 5516 297876 5568
rect 298744 5516 298796 5568
rect 301780 5516 301832 5568
rect 306748 5516 306800 5568
rect 309968 5516 310020 5568
rect 311256 5516 311308 5568
rect 313372 5516 313424 5568
rect 313464 5516 313516 5568
rect 317236 5516 317288 5568
rect 320272 5516 320324 5568
rect 323032 5516 323084 5568
rect 325976 5516 326028 5568
rect 329748 5516 329800 5568
rect 336188 5516 336240 5568
rect 339408 5516 339460 5568
rect 339592 5516 339644 5568
rect 342260 5516 342312 5568
rect 346400 5516 346452 5568
rect 350356 5516 350408 5568
rect 352012 5516 352064 5568
rect 355508 5516 355560 5568
rect 358820 5516 358872 5568
rect 361580 5516 361632 5568
rect 366824 5516 366876 5568
rect 368480 5516 368532 5568
rect 395160 5516 395212 5568
rect 398656 5516 398708 5568
rect 425704 5516 425756 5568
rect 428832 5516 428884 5568
rect 456340 5516 456392 5568
rect 458640 5516 458692 5568
rect 471060 5516 471112 5568
rect 474648 5516 474700 5568
rect 36822 5414 36874 5466
rect 36886 5414 36938 5466
rect 36950 5414 37002 5466
rect 37014 5414 37066 5466
rect 37078 5414 37130 5466
rect 37142 5414 37194 5466
rect 37206 5414 37258 5466
rect 37270 5414 37322 5466
rect 37334 5414 37386 5466
rect 72822 5414 72874 5466
rect 72886 5414 72938 5466
rect 72950 5414 73002 5466
rect 73014 5414 73066 5466
rect 73078 5414 73130 5466
rect 73142 5414 73194 5466
rect 73206 5414 73258 5466
rect 73270 5414 73322 5466
rect 73334 5414 73386 5466
rect 108822 5414 108874 5466
rect 108886 5414 108938 5466
rect 108950 5414 109002 5466
rect 109014 5414 109066 5466
rect 109078 5414 109130 5466
rect 109142 5414 109194 5466
rect 109206 5414 109258 5466
rect 109270 5414 109322 5466
rect 109334 5414 109386 5466
rect 144822 5414 144874 5466
rect 144886 5414 144938 5466
rect 144950 5414 145002 5466
rect 145014 5414 145066 5466
rect 145078 5414 145130 5466
rect 145142 5414 145194 5466
rect 145206 5414 145258 5466
rect 145270 5414 145322 5466
rect 145334 5414 145386 5466
rect 180822 5414 180874 5466
rect 180886 5414 180938 5466
rect 180950 5414 181002 5466
rect 181014 5414 181066 5466
rect 181078 5414 181130 5466
rect 181142 5414 181194 5466
rect 181206 5414 181258 5466
rect 181270 5414 181322 5466
rect 181334 5414 181386 5466
rect 216822 5414 216874 5466
rect 216886 5414 216938 5466
rect 216950 5414 217002 5466
rect 217014 5414 217066 5466
rect 217078 5414 217130 5466
rect 217142 5414 217194 5466
rect 217206 5414 217258 5466
rect 217270 5414 217322 5466
rect 217334 5414 217386 5466
rect 252822 5414 252874 5466
rect 252886 5414 252938 5466
rect 252950 5414 253002 5466
rect 253014 5414 253066 5466
rect 253078 5414 253130 5466
rect 253142 5414 253194 5466
rect 253206 5414 253258 5466
rect 253270 5414 253322 5466
rect 253334 5414 253386 5466
rect 288822 5414 288874 5466
rect 288886 5414 288938 5466
rect 288950 5414 289002 5466
rect 289014 5414 289066 5466
rect 289078 5414 289130 5466
rect 289142 5414 289194 5466
rect 289206 5414 289258 5466
rect 289270 5414 289322 5466
rect 289334 5414 289386 5466
rect 324822 5414 324874 5466
rect 324886 5414 324938 5466
rect 324950 5414 325002 5466
rect 325014 5414 325066 5466
rect 325078 5414 325130 5466
rect 325142 5414 325194 5466
rect 325206 5414 325258 5466
rect 325270 5414 325322 5466
rect 325334 5414 325386 5466
rect 360822 5414 360874 5466
rect 360886 5414 360938 5466
rect 360950 5414 361002 5466
rect 361014 5414 361066 5466
rect 361078 5414 361130 5466
rect 361142 5414 361194 5466
rect 361206 5414 361258 5466
rect 361270 5414 361322 5466
rect 361334 5414 361386 5466
rect 396822 5414 396874 5466
rect 396886 5414 396938 5466
rect 396950 5414 397002 5466
rect 397014 5414 397066 5466
rect 397078 5414 397130 5466
rect 397142 5414 397194 5466
rect 397206 5414 397258 5466
rect 397270 5414 397322 5466
rect 397334 5414 397386 5466
rect 432822 5414 432874 5466
rect 432886 5414 432938 5466
rect 432950 5414 433002 5466
rect 433014 5414 433066 5466
rect 433078 5414 433130 5466
rect 433142 5414 433194 5466
rect 433206 5414 433258 5466
rect 433270 5414 433322 5466
rect 433334 5414 433386 5466
rect 468822 5414 468874 5466
rect 468886 5414 468938 5466
rect 468950 5414 469002 5466
rect 469014 5414 469066 5466
rect 469078 5414 469130 5466
rect 469142 5414 469194 5466
rect 469206 5414 469258 5466
rect 469270 5414 469322 5466
rect 469334 5414 469386 5466
rect 504822 5414 504874 5466
rect 504886 5414 504938 5466
rect 504950 5414 505002 5466
rect 505014 5414 505066 5466
rect 505078 5414 505130 5466
rect 505142 5414 505194 5466
rect 505206 5414 505258 5466
rect 505270 5414 505322 5466
rect 505334 5414 505386 5466
rect 540822 5414 540874 5466
rect 540886 5414 540938 5466
rect 540950 5414 541002 5466
rect 541014 5414 541066 5466
rect 541078 5414 541130 5466
rect 541142 5414 541194 5466
rect 541206 5414 541258 5466
rect 541270 5414 541322 5466
rect 541334 5414 541386 5466
rect 576822 5414 576874 5466
rect 576886 5414 576938 5466
rect 576950 5414 577002 5466
rect 577014 5414 577066 5466
rect 577078 5414 577130 5466
rect 577142 5414 577194 5466
rect 577206 5414 577258 5466
rect 577270 5414 577322 5466
rect 577334 5414 577386 5466
rect 18822 4870 18874 4922
rect 18886 4870 18938 4922
rect 18950 4870 19002 4922
rect 19014 4870 19066 4922
rect 19078 4870 19130 4922
rect 19142 4870 19194 4922
rect 19206 4870 19258 4922
rect 19270 4870 19322 4922
rect 19334 4870 19386 4922
rect 54822 4870 54874 4922
rect 54886 4870 54938 4922
rect 54950 4870 55002 4922
rect 55014 4870 55066 4922
rect 55078 4870 55130 4922
rect 55142 4870 55194 4922
rect 55206 4870 55258 4922
rect 55270 4870 55322 4922
rect 55334 4870 55386 4922
rect 90822 4870 90874 4922
rect 90886 4870 90938 4922
rect 90950 4870 91002 4922
rect 91014 4870 91066 4922
rect 91078 4870 91130 4922
rect 91142 4870 91194 4922
rect 91206 4870 91258 4922
rect 91270 4870 91322 4922
rect 91334 4870 91386 4922
rect 126822 4870 126874 4922
rect 126886 4870 126938 4922
rect 126950 4870 127002 4922
rect 127014 4870 127066 4922
rect 127078 4870 127130 4922
rect 127142 4870 127194 4922
rect 127206 4870 127258 4922
rect 127270 4870 127322 4922
rect 127334 4870 127386 4922
rect 162822 4870 162874 4922
rect 162886 4870 162938 4922
rect 162950 4870 163002 4922
rect 163014 4870 163066 4922
rect 163078 4870 163130 4922
rect 163142 4870 163194 4922
rect 163206 4870 163258 4922
rect 163270 4870 163322 4922
rect 163334 4870 163386 4922
rect 198822 4870 198874 4922
rect 198886 4870 198938 4922
rect 198950 4870 199002 4922
rect 199014 4870 199066 4922
rect 199078 4870 199130 4922
rect 199142 4870 199194 4922
rect 199206 4870 199258 4922
rect 199270 4870 199322 4922
rect 199334 4870 199386 4922
rect 234822 4870 234874 4922
rect 234886 4870 234938 4922
rect 234950 4870 235002 4922
rect 235014 4870 235066 4922
rect 235078 4870 235130 4922
rect 235142 4870 235194 4922
rect 235206 4870 235258 4922
rect 235270 4870 235322 4922
rect 235334 4870 235386 4922
rect 270822 4870 270874 4922
rect 270886 4870 270938 4922
rect 270950 4870 271002 4922
rect 271014 4870 271066 4922
rect 271078 4870 271130 4922
rect 271142 4870 271194 4922
rect 271206 4870 271258 4922
rect 271270 4870 271322 4922
rect 271334 4870 271386 4922
rect 306822 4870 306874 4922
rect 306886 4870 306938 4922
rect 306950 4870 307002 4922
rect 307014 4870 307066 4922
rect 307078 4870 307130 4922
rect 307142 4870 307194 4922
rect 307206 4870 307258 4922
rect 307270 4870 307322 4922
rect 307334 4870 307386 4922
rect 342822 4870 342874 4922
rect 342886 4870 342938 4922
rect 342950 4870 343002 4922
rect 343014 4870 343066 4922
rect 343078 4870 343130 4922
rect 343142 4870 343194 4922
rect 343206 4870 343258 4922
rect 343270 4870 343322 4922
rect 343334 4870 343386 4922
rect 378822 4870 378874 4922
rect 378886 4870 378938 4922
rect 378950 4870 379002 4922
rect 379014 4870 379066 4922
rect 379078 4870 379130 4922
rect 379142 4870 379194 4922
rect 379206 4870 379258 4922
rect 379270 4870 379322 4922
rect 379334 4870 379386 4922
rect 414822 4870 414874 4922
rect 414886 4870 414938 4922
rect 414950 4870 415002 4922
rect 415014 4870 415066 4922
rect 415078 4870 415130 4922
rect 415142 4870 415194 4922
rect 415206 4870 415258 4922
rect 415270 4870 415322 4922
rect 415334 4870 415386 4922
rect 450822 4870 450874 4922
rect 450886 4870 450938 4922
rect 450950 4870 451002 4922
rect 451014 4870 451066 4922
rect 451078 4870 451130 4922
rect 451142 4870 451194 4922
rect 451206 4870 451258 4922
rect 451270 4870 451322 4922
rect 451334 4870 451386 4922
rect 486822 4870 486874 4922
rect 486886 4870 486938 4922
rect 486950 4870 487002 4922
rect 487014 4870 487066 4922
rect 487078 4870 487130 4922
rect 487142 4870 487194 4922
rect 487206 4870 487258 4922
rect 487270 4870 487322 4922
rect 487334 4870 487386 4922
rect 522822 4870 522874 4922
rect 522886 4870 522938 4922
rect 522950 4870 523002 4922
rect 523014 4870 523066 4922
rect 523078 4870 523130 4922
rect 523142 4870 523194 4922
rect 523206 4870 523258 4922
rect 523270 4870 523322 4922
rect 523334 4870 523386 4922
rect 558822 4870 558874 4922
rect 558886 4870 558938 4922
rect 558950 4870 559002 4922
rect 559014 4870 559066 4922
rect 559078 4870 559130 4922
rect 559142 4870 559194 4922
rect 559206 4870 559258 4922
rect 559270 4870 559322 4922
rect 559334 4870 559386 4922
rect 36822 4326 36874 4378
rect 36886 4326 36938 4378
rect 36950 4326 37002 4378
rect 37014 4326 37066 4378
rect 37078 4326 37130 4378
rect 37142 4326 37194 4378
rect 37206 4326 37258 4378
rect 37270 4326 37322 4378
rect 37334 4326 37386 4378
rect 72822 4326 72874 4378
rect 72886 4326 72938 4378
rect 72950 4326 73002 4378
rect 73014 4326 73066 4378
rect 73078 4326 73130 4378
rect 73142 4326 73194 4378
rect 73206 4326 73258 4378
rect 73270 4326 73322 4378
rect 73334 4326 73386 4378
rect 108822 4326 108874 4378
rect 108886 4326 108938 4378
rect 108950 4326 109002 4378
rect 109014 4326 109066 4378
rect 109078 4326 109130 4378
rect 109142 4326 109194 4378
rect 109206 4326 109258 4378
rect 109270 4326 109322 4378
rect 109334 4326 109386 4378
rect 144822 4326 144874 4378
rect 144886 4326 144938 4378
rect 144950 4326 145002 4378
rect 145014 4326 145066 4378
rect 145078 4326 145130 4378
rect 145142 4326 145194 4378
rect 145206 4326 145258 4378
rect 145270 4326 145322 4378
rect 145334 4326 145386 4378
rect 180822 4326 180874 4378
rect 180886 4326 180938 4378
rect 180950 4326 181002 4378
rect 181014 4326 181066 4378
rect 181078 4326 181130 4378
rect 181142 4326 181194 4378
rect 181206 4326 181258 4378
rect 181270 4326 181322 4378
rect 181334 4326 181386 4378
rect 216822 4326 216874 4378
rect 216886 4326 216938 4378
rect 216950 4326 217002 4378
rect 217014 4326 217066 4378
rect 217078 4326 217130 4378
rect 217142 4326 217194 4378
rect 217206 4326 217258 4378
rect 217270 4326 217322 4378
rect 217334 4326 217386 4378
rect 252822 4326 252874 4378
rect 252886 4326 252938 4378
rect 252950 4326 253002 4378
rect 253014 4326 253066 4378
rect 253078 4326 253130 4378
rect 253142 4326 253194 4378
rect 253206 4326 253258 4378
rect 253270 4326 253322 4378
rect 253334 4326 253386 4378
rect 288822 4326 288874 4378
rect 288886 4326 288938 4378
rect 288950 4326 289002 4378
rect 289014 4326 289066 4378
rect 289078 4326 289130 4378
rect 289142 4326 289194 4378
rect 289206 4326 289258 4378
rect 289270 4326 289322 4378
rect 289334 4326 289386 4378
rect 324822 4326 324874 4378
rect 324886 4326 324938 4378
rect 324950 4326 325002 4378
rect 325014 4326 325066 4378
rect 325078 4326 325130 4378
rect 325142 4326 325194 4378
rect 325206 4326 325258 4378
rect 325270 4326 325322 4378
rect 325334 4326 325386 4378
rect 360822 4326 360874 4378
rect 360886 4326 360938 4378
rect 360950 4326 361002 4378
rect 361014 4326 361066 4378
rect 361078 4326 361130 4378
rect 361142 4326 361194 4378
rect 361206 4326 361258 4378
rect 361270 4326 361322 4378
rect 361334 4326 361386 4378
rect 396822 4326 396874 4378
rect 396886 4326 396938 4378
rect 396950 4326 397002 4378
rect 397014 4326 397066 4378
rect 397078 4326 397130 4378
rect 397142 4326 397194 4378
rect 397206 4326 397258 4378
rect 397270 4326 397322 4378
rect 397334 4326 397386 4378
rect 432822 4326 432874 4378
rect 432886 4326 432938 4378
rect 432950 4326 433002 4378
rect 433014 4326 433066 4378
rect 433078 4326 433130 4378
rect 433142 4326 433194 4378
rect 433206 4326 433258 4378
rect 433270 4326 433322 4378
rect 433334 4326 433386 4378
rect 468822 4326 468874 4378
rect 468886 4326 468938 4378
rect 468950 4326 469002 4378
rect 469014 4326 469066 4378
rect 469078 4326 469130 4378
rect 469142 4326 469194 4378
rect 469206 4326 469258 4378
rect 469270 4326 469322 4378
rect 469334 4326 469386 4378
rect 504822 4326 504874 4378
rect 504886 4326 504938 4378
rect 504950 4326 505002 4378
rect 505014 4326 505066 4378
rect 505078 4326 505130 4378
rect 505142 4326 505194 4378
rect 505206 4326 505258 4378
rect 505270 4326 505322 4378
rect 505334 4326 505386 4378
rect 540822 4326 540874 4378
rect 540886 4326 540938 4378
rect 540950 4326 541002 4378
rect 541014 4326 541066 4378
rect 541078 4326 541130 4378
rect 541142 4326 541194 4378
rect 541206 4326 541258 4378
rect 541270 4326 541322 4378
rect 541334 4326 541386 4378
rect 576822 4326 576874 4378
rect 576886 4326 576938 4378
rect 576950 4326 577002 4378
rect 577014 4326 577066 4378
rect 577078 4326 577130 4378
rect 577142 4326 577194 4378
rect 577206 4326 577258 4378
rect 577270 4326 577322 4378
rect 577334 4326 577386 4378
rect 20812 4088 20864 4140
rect 27528 4088 27580 4140
rect 42156 4088 42208 4140
rect 48228 4088 48280 4140
rect 61200 4088 61252 4140
rect 66352 4088 66404 4140
rect 279792 4088 279844 4140
rect 282460 4088 282512 4140
rect 285680 4088 285732 4140
rect 289544 4088 289596 4140
rect 295432 4088 295484 4140
rect 299112 4088 299164 4140
rect 303712 4088 303764 4140
rect 307484 4088 307536 4140
rect 313372 4088 313424 4140
rect 318064 4088 318116 4140
rect 322480 4088 322532 4140
rect 326436 4088 326488 4140
rect 351736 4088 351788 4140
rect 357348 4088 357400 4140
rect 408500 4088 408552 4140
rect 410892 4088 410944 4140
rect 434536 4088 434588 4140
rect 437020 4088 437072 4140
rect 448520 4088 448572 4140
rect 452476 4088 452528 4140
rect 453672 4088 453724 4140
rect 456064 4088 456116 4140
rect 459560 4088 459612 4140
rect 463240 4088 463292 4140
rect 472532 4088 472584 4140
rect 475108 4088 475160 4140
rect 477500 4088 477552 4140
rect 481088 4088 481140 4140
rect 484400 4088 484452 4140
rect 488172 4088 488224 4140
rect 535736 4088 535788 4140
rect 553584 4088 553636 4140
rect 553860 4088 553912 4140
rect 557264 4088 557316 4140
rect 576216 4088 576268 4140
rect 572 4020 624 4072
rect 8576 4020 8628 4072
rect 11244 4020 11296 4072
rect 16948 4020 17000 4072
rect 21916 4020 21968 4072
rect 26240 4020 26292 4072
rect 31484 4020 31536 4072
rect 36452 4020 36504 4072
rect 40960 4020 41012 4072
rect 46848 4020 46900 4072
rect 50528 4020 50580 4072
rect 56140 4020 56192 4072
rect 247040 4020 247092 4072
rect 249156 4020 249208 4072
rect 256700 4020 256752 4072
rect 258632 4020 258684 4072
rect 276020 4020 276072 4072
rect 278872 4020 278924 4072
rect 285772 4020 285824 4072
rect 288348 4020 288400 4072
rect 289452 4020 289504 4072
rect 291936 4020 291988 4072
rect 294328 4020 294380 4072
rect 297916 4020 297968 4072
rect 313096 4020 313148 4072
rect 316960 4020 317012 4072
rect 332416 4020 332468 4072
rect 337108 4020 337160 4072
rect 341800 4020 341852 4072
rect 346676 4020 346728 4072
rect 360752 4020 360804 4072
rect 366916 4020 366968 4072
rect 432696 4020 432748 4072
rect 433524 4020 433576 4072
rect 445760 4020 445812 4072
rect 448980 4020 449032 4072
rect 458180 4020 458232 4072
rect 462044 4020 462096 4072
rect 467840 4020 467892 4072
rect 471520 4020 471572 4072
rect 476120 4020 476172 4072
rect 479892 4020 479944 4072
rect 490748 4020 490800 4072
rect 495348 4020 495400 4072
rect 25504 3952 25556 4004
rect 31668 3952 31720 4004
rect 60004 3952 60056 4004
rect 65248 3952 65300 4004
rect 266452 3952 266504 4004
rect 268108 3952 268160 4004
rect 284392 3952 284444 4004
rect 287152 3952 287204 4004
rect 304264 3952 304316 4004
rect 308588 3952 308640 4004
rect 323032 3952 323084 4004
rect 327632 3952 327684 4004
rect 336280 3952 336332 4004
rect 340696 3952 340748 4004
rect 525800 3952 525852 4004
rect 532240 3952 532292 4004
rect 6460 3884 6512 3936
rect 11060 3884 11112 3936
rect 24308 3884 24360 3936
rect 29000 3884 29052 3936
rect 43352 3884 43404 3936
rect 49332 3884 49384 3936
rect 342720 3884 342772 3936
rect 349068 3884 349120 3936
rect 525524 3884 525576 3936
rect 541440 4020 541492 4072
rect 545948 4020 546000 4072
rect 560576 4020 560628 4072
rect 560668 4020 560720 4072
rect 579804 4020 579856 4072
rect 533436 3952 533488 4004
rect 551192 3952 551244 4004
rect 551560 3952 551612 4004
rect 570236 3952 570288 4004
rect 535920 3884 535972 3936
rect 538128 3884 538180 3936
rect 541624 3884 541676 3936
rect 558368 3884 558420 3936
rect 562968 3884 563020 3936
rect 582196 3884 582248 3936
rect 18822 3782 18874 3834
rect 18886 3782 18938 3834
rect 18950 3782 19002 3834
rect 19014 3782 19066 3834
rect 19078 3782 19130 3834
rect 19142 3782 19194 3834
rect 19206 3782 19258 3834
rect 19270 3782 19322 3834
rect 19334 3782 19386 3834
rect 54822 3782 54874 3834
rect 54886 3782 54938 3834
rect 54950 3782 55002 3834
rect 55014 3782 55066 3834
rect 55078 3782 55130 3834
rect 55142 3782 55194 3834
rect 55206 3782 55258 3834
rect 55270 3782 55322 3834
rect 55334 3782 55386 3834
rect 90822 3782 90874 3834
rect 90886 3782 90938 3834
rect 90950 3782 91002 3834
rect 91014 3782 91066 3834
rect 91078 3782 91130 3834
rect 91142 3782 91194 3834
rect 91206 3782 91258 3834
rect 91270 3782 91322 3834
rect 91334 3782 91386 3834
rect 126822 3782 126874 3834
rect 126886 3782 126938 3834
rect 126950 3782 127002 3834
rect 127014 3782 127066 3834
rect 127078 3782 127130 3834
rect 127142 3782 127194 3834
rect 127206 3782 127258 3834
rect 127270 3782 127322 3834
rect 127334 3782 127386 3834
rect 162822 3782 162874 3834
rect 162886 3782 162938 3834
rect 162950 3782 163002 3834
rect 163014 3782 163066 3834
rect 163078 3782 163130 3834
rect 163142 3782 163194 3834
rect 163206 3782 163258 3834
rect 163270 3782 163322 3834
rect 163334 3782 163386 3834
rect 198822 3782 198874 3834
rect 198886 3782 198938 3834
rect 198950 3782 199002 3834
rect 199014 3782 199066 3834
rect 199078 3782 199130 3834
rect 199142 3782 199194 3834
rect 199206 3782 199258 3834
rect 199270 3782 199322 3834
rect 199334 3782 199386 3834
rect 234822 3782 234874 3834
rect 234886 3782 234938 3834
rect 234950 3782 235002 3834
rect 235014 3782 235066 3834
rect 235078 3782 235130 3834
rect 235142 3782 235194 3834
rect 235206 3782 235258 3834
rect 235270 3782 235322 3834
rect 235334 3782 235386 3834
rect 270822 3782 270874 3834
rect 270886 3782 270938 3834
rect 270950 3782 271002 3834
rect 271014 3782 271066 3834
rect 271078 3782 271130 3834
rect 271142 3782 271194 3834
rect 271206 3782 271258 3834
rect 271270 3782 271322 3834
rect 271334 3782 271386 3834
rect 306822 3782 306874 3834
rect 306886 3782 306938 3834
rect 306950 3782 307002 3834
rect 307014 3782 307066 3834
rect 307078 3782 307130 3834
rect 307142 3782 307194 3834
rect 307206 3782 307258 3834
rect 307270 3782 307322 3834
rect 307334 3782 307386 3834
rect 342822 3782 342874 3834
rect 342886 3782 342938 3834
rect 342950 3782 343002 3834
rect 343014 3782 343066 3834
rect 343078 3782 343130 3834
rect 343142 3782 343194 3834
rect 343206 3782 343258 3834
rect 343270 3782 343322 3834
rect 343334 3782 343386 3834
rect 378822 3782 378874 3834
rect 378886 3782 378938 3834
rect 378950 3782 379002 3834
rect 379014 3782 379066 3834
rect 379078 3782 379130 3834
rect 379142 3782 379194 3834
rect 379206 3782 379258 3834
rect 379270 3782 379322 3834
rect 379334 3782 379386 3834
rect 414822 3782 414874 3834
rect 414886 3782 414938 3834
rect 414950 3782 415002 3834
rect 415014 3782 415066 3834
rect 415078 3782 415130 3834
rect 415142 3782 415194 3834
rect 415206 3782 415258 3834
rect 415270 3782 415322 3834
rect 415334 3782 415386 3834
rect 450822 3782 450874 3834
rect 450886 3782 450938 3834
rect 450950 3782 451002 3834
rect 451014 3782 451066 3834
rect 451078 3782 451130 3834
rect 451142 3782 451194 3834
rect 451206 3782 451258 3834
rect 451270 3782 451322 3834
rect 451334 3782 451386 3834
rect 486822 3782 486874 3834
rect 486886 3782 486938 3834
rect 486950 3782 487002 3834
rect 487014 3782 487066 3834
rect 487078 3782 487130 3834
rect 487142 3782 487194 3834
rect 487206 3782 487258 3834
rect 487270 3782 487322 3834
rect 487334 3782 487386 3834
rect 522822 3782 522874 3834
rect 522886 3782 522938 3834
rect 522950 3782 523002 3834
rect 523014 3782 523066 3834
rect 523078 3782 523130 3834
rect 523142 3782 523194 3834
rect 523206 3782 523258 3834
rect 523270 3782 523322 3834
rect 523334 3782 523386 3834
rect 558822 3782 558874 3834
rect 558886 3782 558938 3834
rect 558950 3782 559002 3834
rect 559014 3782 559066 3834
rect 559078 3782 559130 3834
rect 559142 3782 559194 3834
rect 559206 3782 559258 3834
rect 559270 3782 559322 3834
rect 559334 3782 559386 3834
rect 266360 3680 266412 3732
rect 269304 3680 269356 3732
rect 275100 3680 275152 3732
rect 277676 3680 277728 3732
rect 292580 3680 292632 3732
rect 296720 3680 296772 3732
rect 464436 3680 464488 3732
rect 467932 3680 467984 3732
rect 469496 3680 469548 3732
rect 472716 3680 472768 3732
rect 474096 3680 474148 3732
rect 477500 3680 477552 3732
rect 510436 3680 510488 3732
rect 515588 3680 515640 3732
rect 524512 3680 524564 3732
rect 531044 3680 531096 3732
rect 531228 3680 531280 3732
rect 548892 3680 548944 3732
rect 550456 3680 550508 3732
rect 552756 3680 552808 3732
rect 571432 3680 571484 3732
rect 29092 3612 29144 3664
rect 35716 3612 35768 3664
rect 45744 3612 45796 3664
rect 51632 3612 51684 3664
rect 64788 3612 64840 3664
rect 69756 3612 69808 3664
rect 332968 3612 333020 3664
rect 338304 3612 338356 3664
rect 342260 3612 342312 3664
rect 347872 3612 347924 3664
rect 413376 3612 413428 3664
rect 421564 3612 421616 3664
rect 472900 3612 472952 3664
rect 476304 3612 476356 3664
rect 478972 3612 479024 3664
rect 483480 3612 483532 3664
rect 518716 3612 518768 3664
rect 535736 3612 535788 3664
rect 538036 3612 538088 3664
rect 559472 3612 559524 3664
rect 559564 3612 559616 3664
rect 578608 3612 578660 3664
rect 5264 3544 5316 3596
rect 12256 3544 12308 3596
rect 16028 3544 16080 3596
rect 20720 3544 20772 3596
rect 34980 3544 35032 3596
rect 41328 3544 41380 3596
rect 44548 3544 44600 3596
rect 50436 3544 50488 3596
rect 52828 3544 52880 3596
rect 58440 3544 58492 3596
rect 74264 3544 74316 3596
rect 78864 3544 78916 3596
rect 292488 3544 292540 3596
rect 295524 3544 295576 3596
rect 305000 3544 305052 3596
rect 309784 3544 309836 3596
rect 311808 3544 311860 3596
rect 315764 3544 315816 3596
rect 324320 3544 324372 3596
rect 330024 3544 330076 3596
rect 333980 3544 334032 3596
rect 339500 3544 339552 3596
rect 352288 3544 352340 3596
rect 358544 3544 358596 3596
rect 367468 3544 367520 3596
rect 374000 3544 374052 3596
rect 433892 3544 433944 3596
rect 435824 3544 435876 3596
rect 456800 3544 456852 3596
rect 459652 3544 459704 3596
rect 463332 3544 463384 3596
rect 465632 3544 465684 3596
rect 488540 3544 488592 3596
rect 492956 3544 493008 3596
rect 496820 3544 496872 3596
rect 501236 3544 501288 3596
rect 510528 3544 510580 3596
rect 514392 3544 514444 3596
rect 519820 3544 519872 3596
rect 536932 3544 536984 3596
rect 7656 3476 7708 3528
rect 15016 3476 15068 3528
rect 17224 3476 17276 3528
rect 23112 3476 23164 3528
rect 26700 3476 26752 3528
rect 31760 3476 31812 3528
rect 33876 3476 33928 3528
rect 39948 3476 40000 3528
rect 51632 3476 51684 3528
rect 57244 3476 57296 3528
rect 57612 3476 57664 3528
rect 62948 3476 63000 3528
rect 65984 3476 66036 3528
rect 70860 3476 70912 3528
rect 72700 3476 72752 3528
rect 77668 3476 77720 3528
rect 149244 3476 149296 3528
rect 150256 3476 150308 3528
rect 150440 3476 150492 3528
rect 151360 3476 151412 3528
rect 156328 3476 156380 3528
rect 157064 3476 157116 3528
rect 187700 3476 187752 3528
rect 188436 3476 188488 3528
rect 193312 3476 193364 3528
rect 194416 3476 194468 3528
rect 255412 3476 255464 3528
rect 257436 3476 257488 3528
rect 262404 3476 262456 3528
rect 264612 3476 264664 3528
rect 264980 3476 265032 3528
rect 267004 3476 267056 3528
rect 282092 3476 282144 3528
rect 284760 3476 284812 3528
rect 290188 3476 290240 3528
rect 293132 3476 293184 3528
rect 300676 3476 300728 3528
rect 303804 3476 303856 3528
rect 311164 3476 311216 3528
rect 314568 3476 314620 3528
rect 323584 3476 323636 3528
rect 328828 3476 328880 3528
rect 329748 3476 329800 3528
rect 333612 3476 333664 3528
rect 339408 3476 339460 3528
rect 344284 3476 344336 3528
rect 353300 3476 353352 3528
rect 359740 3476 359792 3528
rect 474648 3476 474700 3528
rect 4068 3408 4120 3460
rect 11612 3408 11664 3460
rect 14832 3408 14884 3460
rect 19432 3408 19484 3460
rect 27896 3408 27948 3460
rect 34336 3408 34388 3460
rect 38568 3408 38620 3460
rect 42800 3408 42852 3460
rect 48136 3408 48188 3460
rect 53656 3408 53708 3460
rect 54024 3408 54076 3460
rect 59544 3408 59596 3460
rect 68284 3408 68336 3460
rect 73436 3408 73488 3460
rect 254216 3408 254268 3460
rect 256240 3408 256292 3460
rect 261208 3408 261260 3460
rect 263416 3408 263468 3460
rect 263692 3408 263744 3460
rect 265808 3408 265860 3460
rect 270500 3408 270552 3460
rect 272892 3408 272944 3460
rect 272984 3408 273036 3460
rect 275284 3408 275336 3460
rect 299204 3408 299256 3460
rect 302608 3408 302660 3460
rect 303068 3408 303120 3460
rect 306196 3408 306248 3460
rect 309968 3408 310020 3460
rect 313372 3408 313424 3460
rect 314660 3408 314712 3460
rect 319260 3408 319312 3460
rect 320088 3408 320140 3460
rect 324044 3408 324096 3460
rect 330852 3408 330904 3460
rect 334716 3408 334768 3460
rect 343640 3408 343692 3460
rect 350264 3408 350316 3460
rect 350356 3408 350408 3460
rect 354956 3408 355008 3460
rect 361580 3408 361632 3460
rect 368020 3408 368072 3460
rect 382280 3408 382332 3460
rect 390652 3408 390704 3460
rect 398656 3408 398708 3460
rect 406108 3408 406160 3460
rect 413928 3408 413980 3460
rect 422760 3408 422812 3460
rect 426440 3408 426492 3460
rect 428740 3408 428792 3460
rect 428832 3408 428884 3460
rect 438216 3408 438268 3460
rect 444288 3408 444340 3460
rect 453672 3408 453724 3460
rect 458640 3408 458692 3460
rect 8852 3340 8904 3392
rect 13820 3340 13872 3392
rect 18328 3340 18380 3392
rect 23848 3340 23900 3392
rect 36176 3340 36228 3392
rect 42524 3340 42576 3392
rect 58808 3340 58860 3392
rect 64052 3340 64104 3392
rect 280896 3340 280948 3392
rect 283656 3340 283708 3392
rect 291384 3340 291436 3392
rect 294328 3340 294380 3392
rect 301780 3340 301832 3392
rect 305000 3340 305052 3392
rect 321468 3340 321520 3392
rect 325424 3340 325476 3392
rect 348976 3340 349028 3392
rect 353760 3340 353812 3392
rect 368480 3340 368532 3392
rect 376392 3340 376444 3392
rect 394056 3340 394108 3392
rect 395436 3340 395488 3392
rect 429200 3340 429252 3392
rect 431132 3340 431184 3392
rect 437480 3340 437532 3392
rect 439412 3340 439464 3392
rect 442356 3340 442408 3392
rect 444196 3340 444248 3392
rect 445852 3340 445904 3392
rect 447784 3340 447836 3392
rect 453120 3340 453172 3392
rect 454868 3340 454920 3392
rect 462228 3408 462280 3460
rect 464436 3408 464488 3460
rect 469404 3408 469456 3460
rect 473912 3408 473964 3460
rect 474740 3408 474792 3460
rect 478696 3408 478748 3460
rect 478880 3476 478932 3528
rect 484584 3476 484636 3528
rect 506480 3476 506532 3528
rect 512000 3476 512052 3528
rect 527824 3476 527876 3528
rect 485780 3408 485832 3460
rect 491208 3408 491260 3460
rect 503628 3408 503680 3460
rect 511724 3408 511776 3460
rect 528652 3408 528704 3460
rect 534632 3408 534684 3460
rect 542544 3544 542596 3596
rect 547788 3544 547840 3596
rect 563152 3544 563204 3596
rect 564532 3544 564584 3596
rect 545304 3476 545356 3528
rect 546592 3476 546644 3528
rect 547052 3476 547104 3528
rect 569040 3476 569092 3528
rect 539140 3408 539192 3460
rect 544752 3408 544804 3460
rect 547604 3408 547656 3460
rect 470324 3340 470376 3392
rect 477592 3340 477644 3392
rect 482284 3340 482336 3392
rect 487436 3340 487488 3392
rect 491760 3340 491812 3392
rect 503904 3340 503956 3392
rect 509608 3340 509660 3392
rect 520832 3340 520884 3392
rect 522672 3340 522724 3392
rect 542912 3340 542964 3392
rect 543648 3340 543700 3392
rect 547788 3340 547840 3392
rect 558368 3340 558420 3392
rect 561680 3408 561732 3460
rect 561772 3408 561824 3460
rect 581000 3408 581052 3460
rect 561956 3340 562008 3392
rect 577412 3340 577464 3392
rect 36822 3238 36874 3290
rect 36886 3238 36938 3290
rect 36950 3238 37002 3290
rect 37014 3238 37066 3290
rect 37078 3238 37130 3290
rect 37142 3238 37194 3290
rect 37206 3238 37258 3290
rect 37270 3238 37322 3290
rect 37334 3238 37386 3290
rect 72822 3238 72874 3290
rect 72886 3238 72938 3290
rect 72950 3238 73002 3290
rect 73014 3238 73066 3290
rect 73078 3238 73130 3290
rect 73142 3238 73194 3290
rect 73206 3238 73258 3290
rect 73270 3238 73322 3290
rect 73334 3238 73386 3290
rect 108822 3238 108874 3290
rect 108886 3238 108938 3290
rect 108950 3238 109002 3290
rect 109014 3238 109066 3290
rect 109078 3238 109130 3290
rect 109142 3238 109194 3290
rect 109206 3238 109258 3290
rect 109270 3238 109322 3290
rect 109334 3238 109386 3290
rect 144822 3238 144874 3290
rect 144886 3238 144938 3290
rect 144950 3238 145002 3290
rect 145014 3238 145066 3290
rect 145078 3238 145130 3290
rect 145142 3238 145194 3290
rect 145206 3238 145258 3290
rect 145270 3238 145322 3290
rect 145334 3238 145386 3290
rect 180822 3238 180874 3290
rect 180886 3238 180938 3290
rect 180950 3238 181002 3290
rect 181014 3238 181066 3290
rect 181078 3238 181130 3290
rect 181142 3238 181194 3290
rect 181206 3238 181258 3290
rect 181270 3238 181322 3290
rect 181334 3238 181386 3290
rect 216822 3238 216874 3290
rect 216886 3238 216938 3290
rect 216950 3238 217002 3290
rect 217014 3238 217066 3290
rect 217078 3238 217130 3290
rect 217142 3238 217194 3290
rect 217206 3238 217258 3290
rect 217270 3238 217322 3290
rect 217334 3238 217386 3290
rect 252822 3238 252874 3290
rect 252886 3238 252938 3290
rect 252950 3238 253002 3290
rect 253014 3238 253066 3290
rect 253078 3238 253130 3290
rect 253142 3238 253194 3290
rect 253206 3238 253258 3290
rect 253270 3238 253322 3290
rect 253334 3238 253386 3290
rect 288822 3238 288874 3290
rect 288886 3238 288938 3290
rect 288950 3238 289002 3290
rect 289014 3238 289066 3290
rect 289078 3238 289130 3290
rect 289142 3238 289194 3290
rect 289206 3238 289258 3290
rect 289270 3238 289322 3290
rect 289334 3238 289386 3290
rect 324822 3238 324874 3290
rect 324886 3238 324938 3290
rect 324950 3238 325002 3290
rect 325014 3238 325066 3290
rect 325078 3238 325130 3290
rect 325142 3238 325194 3290
rect 325206 3238 325258 3290
rect 325270 3238 325322 3290
rect 325334 3238 325386 3290
rect 360822 3238 360874 3290
rect 360886 3238 360938 3290
rect 360950 3238 361002 3290
rect 361014 3238 361066 3290
rect 361078 3238 361130 3290
rect 361142 3238 361194 3290
rect 361206 3238 361258 3290
rect 361270 3238 361322 3290
rect 361334 3238 361386 3290
rect 396822 3238 396874 3290
rect 396886 3238 396938 3290
rect 396950 3238 397002 3290
rect 397014 3238 397066 3290
rect 397078 3238 397130 3290
rect 397142 3238 397194 3290
rect 397206 3238 397258 3290
rect 397270 3238 397322 3290
rect 397334 3238 397386 3290
rect 432822 3238 432874 3290
rect 432886 3238 432938 3290
rect 432950 3238 433002 3290
rect 433014 3238 433066 3290
rect 433078 3238 433130 3290
rect 433142 3238 433194 3290
rect 433206 3238 433258 3290
rect 433270 3238 433322 3290
rect 433334 3238 433386 3290
rect 468822 3238 468874 3290
rect 468886 3238 468938 3290
rect 468950 3238 469002 3290
rect 469014 3238 469066 3290
rect 469078 3238 469130 3290
rect 469142 3238 469194 3290
rect 469206 3238 469258 3290
rect 469270 3238 469322 3290
rect 469334 3238 469386 3290
rect 504822 3238 504874 3290
rect 504886 3238 504938 3290
rect 504950 3238 505002 3290
rect 505014 3238 505066 3290
rect 505078 3238 505130 3290
rect 505142 3238 505194 3290
rect 505206 3238 505258 3290
rect 505270 3238 505322 3290
rect 505334 3238 505386 3290
rect 540822 3238 540874 3290
rect 540886 3238 540938 3290
rect 540950 3238 541002 3290
rect 541014 3238 541066 3290
rect 541078 3238 541130 3290
rect 541142 3238 541194 3290
rect 541206 3238 541258 3290
rect 541270 3238 541322 3290
rect 541334 3238 541386 3290
rect 576822 3238 576874 3290
rect 576886 3238 576938 3290
rect 576950 3238 577002 3290
rect 577014 3238 577066 3290
rect 577078 3238 577130 3290
rect 577142 3238 577194 3290
rect 577206 3238 577258 3290
rect 577270 3238 577322 3290
rect 577334 3238 577386 3290
rect 13636 3136 13688 3188
rect 18604 3136 18656 3188
rect 23112 3136 23164 3188
rect 27712 3136 27764 3188
rect 49332 3136 49384 3188
rect 54668 3136 54720 3188
rect 56416 3136 56468 3188
rect 61844 3136 61896 3188
rect 67180 3136 67232 3188
rect 72056 3136 72108 3188
rect 273996 3136 274048 3188
rect 276480 3136 276532 3188
rect 283196 3136 283248 3188
rect 285956 3136 286008 3188
rect 307668 3136 307720 3188
rect 310980 3136 311032 3188
rect 317236 3136 317288 3188
rect 320456 3136 320508 3188
rect 326988 3136 327040 3188
rect 331220 3136 331272 3188
rect 336648 3136 336700 3188
rect 341892 3136 341944 3188
rect 345940 3136 345992 3188
rect 351368 3136 351420 3188
rect 367100 3136 367152 3188
rect 375196 3136 375248 3188
rect 414112 3136 414164 3188
rect 415676 3136 415728 3188
rect 418160 3136 418212 3188
rect 420368 3136 420420 3188
rect 427820 3136 427872 3188
rect 429936 3136 429988 3188
rect 430580 3136 430632 3188
rect 432328 3136 432380 3188
rect 438952 3136 439004 3188
rect 440608 3136 440660 3188
rect 443552 3136 443604 3188
rect 445392 3136 445444 3188
rect 448612 3136 448664 3188
rect 451464 3136 451516 3188
rect 454132 3136 454184 3188
rect 457260 3136 457312 3188
rect 458272 3136 458324 3188
rect 460848 3136 460900 3188
rect 483296 3136 483348 3188
rect 486700 3136 486752 3188
rect 514760 3136 514812 3188
rect 520280 3136 520332 3188
rect 540244 3136 540296 3188
rect 547696 3136 547748 3188
rect 2872 3068 2924 3120
rect 5540 3068 5592 3120
rect 32680 3068 32732 3120
rect 37464 3068 37516 3120
rect 46940 3068 46992 3120
rect 52736 3068 52788 3120
rect 318248 3068 318300 3120
rect 321652 3068 321704 3120
rect 330576 3068 330628 3120
rect 335912 3068 335964 3120
rect 339684 3068 339736 3120
rect 345480 3068 345532 3120
rect 424324 3068 424376 3120
rect 426348 3068 426400 3120
rect 438860 3068 438912 3120
rect 441804 3068 441856 3120
rect 447140 3068 447192 3120
rect 450176 3068 450228 3120
rect 454684 3068 454736 3120
rect 458456 3068 458508 3120
rect 463700 3068 463752 3120
rect 466828 3068 466880 3120
rect 484676 3068 484728 3120
rect 490564 3068 490616 3120
rect 500592 3068 500644 3120
rect 504732 3068 504784 3120
rect 526628 3068 526680 3120
rect 544108 3068 544160 3120
rect 557172 3136 557224 3188
rect 575020 3136 575072 3188
rect 555976 3068 556028 3120
rect 556160 3068 556212 3120
rect 12440 3000 12492 3052
rect 18052 3000 18104 3052
rect 269672 3000 269724 3052
rect 271696 3000 271748 3052
rect 271880 3000 271932 3052
rect 274088 3000 274140 3052
rect 279332 3000 279384 3052
rect 281264 3000 281316 3052
rect 298928 3000 298980 3052
rect 301412 3000 301464 3052
rect 318708 3000 318760 3052
rect 322848 3000 322900 3052
rect 328276 3000 328328 3052
rect 332416 3000 332468 3052
rect 347412 3000 347464 3052
rect 352564 3000 352616 3052
rect 403808 3000 403860 3052
rect 404912 3000 404964 3052
rect 439044 3000 439096 3052
rect 443000 3000 443052 3052
rect 444380 3000 444432 3052
rect 446588 3000 446640 3052
rect 464252 3000 464304 3052
rect 468668 3000 468720 3052
rect 494152 3000 494204 3052
rect 498936 3000 498988 3052
rect 503996 3000 504048 3052
rect 508412 3000 508464 3052
rect 521200 3000 521252 3052
rect 526260 3000 526312 3052
rect 536840 3000 536892 3052
rect 566740 3068 566792 3120
rect 573824 3068 573876 3120
rect 37464 2932 37516 2984
rect 43720 2932 43772 2984
rect 260104 2932 260156 2984
rect 262220 2932 262272 2984
rect 337384 2932 337436 2984
rect 342720 2932 342772 2984
rect 511908 2932 511960 2984
rect 516784 2932 516836 2984
rect 522396 2932 522448 2984
rect 527456 2932 527508 2984
rect 536748 2932 536800 2984
rect 541716 2932 541768 2984
rect 552388 2932 552440 2984
rect 1676 2864 1728 2916
rect 9588 2864 9640 2916
rect 10048 2864 10100 2916
rect 15200 2864 15252 2916
rect 240140 2864 240192 2916
rect 241980 2864 242032 2916
rect 249248 2864 249300 2916
rect 250352 2864 250404 2916
rect 259000 2864 259052 2916
rect 259828 2864 259880 2916
rect 269028 2864 269080 2916
rect 270500 2864 270552 2916
rect 288256 2864 288308 2916
rect 290740 2864 290792 2916
rect 297824 2864 297876 2916
rect 300308 2864 300360 2916
rect 384948 2864 385000 2916
rect 391848 2864 391900 2916
rect 491116 2864 491168 2916
rect 494152 2864 494204 2916
rect 528928 2864 528980 2916
rect 546500 2864 546552 2916
rect 546592 2864 546644 2916
rect 547696 2864 547748 2916
rect 548156 2864 548208 2916
rect 554964 2932 555016 2984
rect 564348 2932 564400 2984
rect 572628 2932 572680 2984
rect 565544 2864 565596 2916
rect 19524 2796 19576 2848
rect 26148 2796 26200 2848
rect 30288 2796 30340 2848
rect 34520 2796 34572 2848
rect 39764 2796 39816 2848
rect 45468 2796 45520 2848
rect 278412 2796 278464 2848
rect 280068 2796 280120 2848
rect 308220 2796 308272 2848
rect 312176 2796 312228 2848
rect 355508 2796 355560 2848
rect 360752 2796 360804 2848
rect 532332 2796 532384 2848
rect 550088 2796 550140 2848
rect 550548 2796 550600 2848
rect 567844 2796 567896 2848
rect 18822 2694 18874 2746
rect 18886 2694 18938 2746
rect 18950 2694 19002 2746
rect 19014 2694 19066 2746
rect 19078 2694 19130 2746
rect 19142 2694 19194 2746
rect 19206 2694 19258 2746
rect 19270 2694 19322 2746
rect 19334 2694 19386 2746
rect 54822 2694 54874 2746
rect 54886 2694 54938 2746
rect 54950 2694 55002 2746
rect 55014 2694 55066 2746
rect 55078 2694 55130 2746
rect 55142 2694 55194 2746
rect 55206 2694 55258 2746
rect 55270 2694 55322 2746
rect 55334 2694 55386 2746
rect 90822 2694 90874 2746
rect 90886 2694 90938 2746
rect 90950 2694 91002 2746
rect 91014 2694 91066 2746
rect 91078 2694 91130 2746
rect 91142 2694 91194 2746
rect 91206 2694 91258 2746
rect 91270 2694 91322 2746
rect 91334 2694 91386 2746
rect 126822 2694 126874 2746
rect 126886 2694 126938 2746
rect 126950 2694 127002 2746
rect 127014 2694 127066 2746
rect 127078 2694 127130 2746
rect 127142 2694 127194 2746
rect 127206 2694 127258 2746
rect 127270 2694 127322 2746
rect 127334 2694 127386 2746
rect 162822 2694 162874 2746
rect 162886 2694 162938 2746
rect 162950 2694 163002 2746
rect 163014 2694 163066 2746
rect 163078 2694 163130 2746
rect 163142 2694 163194 2746
rect 163206 2694 163258 2746
rect 163270 2694 163322 2746
rect 163334 2694 163386 2746
rect 198822 2694 198874 2746
rect 198886 2694 198938 2746
rect 198950 2694 199002 2746
rect 199014 2694 199066 2746
rect 199078 2694 199130 2746
rect 199142 2694 199194 2746
rect 199206 2694 199258 2746
rect 199270 2694 199322 2746
rect 199334 2694 199386 2746
rect 234822 2694 234874 2746
rect 234886 2694 234938 2746
rect 234950 2694 235002 2746
rect 235014 2694 235066 2746
rect 235078 2694 235130 2746
rect 235142 2694 235194 2746
rect 235206 2694 235258 2746
rect 235270 2694 235322 2746
rect 235334 2694 235386 2746
rect 270822 2694 270874 2746
rect 270886 2694 270938 2746
rect 270950 2694 271002 2746
rect 271014 2694 271066 2746
rect 271078 2694 271130 2746
rect 271142 2694 271194 2746
rect 271206 2694 271258 2746
rect 271270 2694 271322 2746
rect 271334 2694 271386 2746
rect 306822 2694 306874 2746
rect 306886 2694 306938 2746
rect 306950 2694 307002 2746
rect 307014 2694 307066 2746
rect 307078 2694 307130 2746
rect 307142 2694 307194 2746
rect 307206 2694 307258 2746
rect 307270 2694 307322 2746
rect 307334 2694 307386 2746
rect 342822 2694 342874 2746
rect 342886 2694 342938 2746
rect 342950 2694 343002 2746
rect 343014 2694 343066 2746
rect 343078 2694 343130 2746
rect 343142 2694 343194 2746
rect 343206 2694 343258 2746
rect 343270 2694 343322 2746
rect 343334 2694 343386 2746
rect 378822 2694 378874 2746
rect 378886 2694 378938 2746
rect 378950 2694 379002 2746
rect 379014 2694 379066 2746
rect 379078 2694 379130 2746
rect 379142 2694 379194 2746
rect 379206 2694 379258 2746
rect 379270 2694 379322 2746
rect 379334 2694 379386 2746
rect 414822 2694 414874 2746
rect 414886 2694 414938 2746
rect 414950 2694 415002 2746
rect 415014 2694 415066 2746
rect 415078 2694 415130 2746
rect 415142 2694 415194 2746
rect 415206 2694 415258 2746
rect 415270 2694 415322 2746
rect 415334 2694 415386 2746
rect 450822 2694 450874 2746
rect 450886 2694 450938 2746
rect 450950 2694 451002 2746
rect 451014 2694 451066 2746
rect 451078 2694 451130 2746
rect 451142 2694 451194 2746
rect 451206 2694 451258 2746
rect 451270 2694 451322 2746
rect 451334 2694 451386 2746
rect 486822 2694 486874 2746
rect 486886 2694 486938 2746
rect 486950 2694 487002 2746
rect 487014 2694 487066 2746
rect 487078 2694 487130 2746
rect 487142 2694 487194 2746
rect 487206 2694 487258 2746
rect 487270 2694 487322 2746
rect 487334 2694 487386 2746
rect 522822 2694 522874 2746
rect 522886 2694 522938 2746
rect 522950 2694 523002 2746
rect 523014 2694 523066 2746
rect 523078 2694 523130 2746
rect 523142 2694 523194 2746
rect 523206 2694 523258 2746
rect 523270 2694 523322 2746
rect 523334 2694 523386 2746
rect 558822 2694 558874 2746
rect 558886 2694 558938 2746
rect 558950 2694 559002 2746
rect 559014 2694 559066 2746
rect 559078 2694 559130 2746
rect 559142 2694 559194 2746
rect 559206 2694 559258 2746
rect 559270 2694 559322 2746
rect 559334 2694 559386 2746
rect 554780 2592 554832 2644
rect 36822 2150 36874 2202
rect 36886 2150 36938 2202
rect 36950 2150 37002 2202
rect 37014 2150 37066 2202
rect 37078 2150 37130 2202
rect 37142 2150 37194 2202
rect 37206 2150 37258 2202
rect 37270 2150 37322 2202
rect 37334 2150 37386 2202
rect 72822 2150 72874 2202
rect 72886 2150 72938 2202
rect 72950 2150 73002 2202
rect 73014 2150 73066 2202
rect 73078 2150 73130 2202
rect 73142 2150 73194 2202
rect 73206 2150 73258 2202
rect 73270 2150 73322 2202
rect 73334 2150 73386 2202
rect 108822 2150 108874 2202
rect 108886 2150 108938 2202
rect 108950 2150 109002 2202
rect 109014 2150 109066 2202
rect 109078 2150 109130 2202
rect 109142 2150 109194 2202
rect 109206 2150 109258 2202
rect 109270 2150 109322 2202
rect 109334 2150 109386 2202
rect 144822 2150 144874 2202
rect 144886 2150 144938 2202
rect 144950 2150 145002 2202
rect 145014 2150 145066 2202
rect 145078 2150 145130 2202
rect 145142 2150 145194 2202
rect 145206 2150 145258 2202
rect 145270 2150 145322 2202
rect 145334 2150 145386 2202
rect 180822 2150 180874 2202
rect 180886 2150 180938 2202
rect 180950 2150 181002 2202
rect 181014 2150 181066 2202
rect 181078 2150 181130 2202
rect 181142 2150 181194 2202
rect 181206 2150 181258 2202
rect 181270 2150 181322 2202
rect 181334 2150 181386 2202
rect 216822 2150 216874 2202
rect 216886 2150 216938 2202
rect 216950 2150 217002 2202
rect 217014 2150 217066 2202
rect 217078 2150 217130 2202
rect 217142 2150 217194 2202
rect 217206 2150 217258 2202
rect 217270 2150 217322 2202
rect 217334 2150 217386 2202
rect 252822 2150 252874 2202
rect 252886 2150 252938 2202
rect 252950 2150 253002 2202
rect 253014 2150 253066 2202
rect 253078 2150 253130 2202
rect 253142 2150 253194 2202
rect 253206 2150 253258 2202
rect 253270 2150 253322 2202
rect 253334 2150 253386 2202
rect 288822 2150 288874 2202
rect 288886 2150 288938 2202
rect 288950 2150 289002 2202
rect 289014 2150 289066 2202
rect 289078 2150 289130 2202
rect 289142 2150 289194 2202
rect 289206 2150 289258 2202
rect 289270 2150 289322 2202
rect 289334 2150 289386 2202
rect 324822 2150 324874 2202
rect 324886 2150 324938 2202
rect 324950 2150 325002 2202
rect 325014 2150 325066 2202
rect 325078 2150 325130 2202
rect 325142 2150 325194 2202
rect 325206 2150 325258 2202
rect 325270 2150 325322 2202
rect 325334 2150 325386 2202
rect 360822 2150 360874 2202
rect 360886 2150 360938 2202
rect 360950 2150 361002 2202
rect 361014 2150 361066 2202
rect 361078 2150 361130 2202
rect 361142 2150 361194 2202
rect 361206 2150 361258 2202
rect 361270 2150 361322 2202
rect 361334 2150 361386 2202
rect 396822 2150 396874 2202
rect 396886 2150 396938 2202
rect 396950 2150 397002 2202
rect 397014 2150 397066 2202
rect 397078 2150 397130 2202
rect 397142 2150 397194 2202
rect 397206 2150 397258 2202
rect 397270 2150 397322 2202
rect 397334 2150 397386 2202
rect 432822 2150 432874 2202
rect 432886 2150 432938 2202
rect 432950 2150 433002 2202
rect 433014 2150 433066 2202
rect 433078 2150 433130 2202
rect 433142 2150 433194 2202
rect 433206 2150 433258 2202
rect 433270 2150 433322 2202
rect 433334 2150 433386 2202
rect 468822 2150 468874 2202
rect 468886 2150 468938 2202
rect 468950 2150 469002 2202
rect 469014 2150 469066 2202
rect 469078 2150 469130 2202
rect 469142 2150 469194 2202
rect 469206 2150 469258 2202
rect 469270 2150 469322 2202
rect 469334 2150 469386 2202
rect 504822 2150 504874 2202
rect 504886 2150 504938 2202
rect 504950 2150 505002 2202
rect 505014 2150 505066 2202
rect 505078 2150 505130 2202
rect 505142 2150 505194 2202
rect 505206 2150 505258 2202
rect 505270 2150 505322 2202
rect 505334 2150 505386 2202
rect 540822 2150 540874 2202
rect 540886 2150 540938 2202
rect 540950 2150 541002 2202
rect 541014 2150 541066 2202
rect 541078 2150 541130 2202
rect 541142 2150 541194 2202
rect 541206 2150 541258 2202
rect 541270 2150 541322 2202
rect 541334 2150 541386 2202
rect 576822 2150 576874 2202
rect 576886 2150 576938 2202
rect 576950 2150 577002 2202
rect 577014 2150 577066 2202
rect 577078 2150 577130 2202
rect 577142 2150 577194 2202
rect 577206 2150 577258 2202
rect 577270 2150 577322 2202
rect 577334 2150 577386 2202
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 700369 8156 703520
rect 18822 701244 19386 701264
rect 18822 701242 18836 701244
rect 18892 701242 18916 701244
rect 18972 701242 18996 701244
rect 19052 701242 19076 701244
rect 19132 701242 19156 701244
rect 19212 701242 19236 701244
rect 19292 701242 19316 701244
rect 19372 701242 19386 701244
rect 19066 701190 19076 701242
rect 19132 701190 19142 701242
rect 18822 701188 18836 701190
rect 18892 701188 18916 701190
rect 18972 701188 18996 701190
rect 19052 701188 19076 701190
rect 19132 701188 19156 701190
rect 19212 701188 19236 701190
rect 19292 701188 19316 701190
rect 19372 701188 19386 701190
rect 18822 701168 19386 701188
rect 24320 700505 24348 703520
rect 36822 701788 37386 701808
rect 36822 701786 36836 701788
rect 36892 701786 36916 701788
rect 36972 701786 36996 701788
rect 37052 701786 37076 701788
rect 37132 701786 37156 701788
rect 37212 701786 37236 701788
rect 37292 701786 37316 701788
rect 37372 701786 37386 701788
rect 37066 701734 37076 701786
rect 37132 701734 37142 701786
rect 36822 701732 36836 701734
rect 36892 701732 36916 701734
rect 36972 701732 36996 701734
rect 37052 701732 37076 701734
rect 37132 701732 37156 701734
rect 37212 701732 37236 701734
rect 37292 701732 37316 701734
rect 37372 701732 37386 701734
rect 36822 701712 37386 701732
rect 40512 701049 40540 703520
rect 72988 701978 73016 703520
rect 72712 701950 73016 701978
rect 54822 701244 55386 701264
rect 54822 701242 54836 701244
rect 54892 701242 54916 701244
rect 54972 701242 54996 701244
rect 55052 701242 55076 701244
rect 55132 701242 55156 701244
rect 55212 701242 55236 701244
rect 55292 701242 55316 701244
rect 55372 701242 55386 701244
rect 55066 701190 55076 701242
rect 55132 701190 55142 701242
rect 54822 701188 54836 701190
rect 54892 701188 54916 701190
rect 54972 701188 54996 701190
rect 55052 701188 55076 701190
rect 55132 701188 55156 701190
rect 55212 701188 55236 701190
rect 55292 701188 55316 701190
rect 55372 701188 55386 701190
rect 54822 701168 55386 701188
rect 40498 701040 40554 701049
rect 40498 700975 40554 700984
rect 36822 700700 37386 700720
rect 36822 700698 36836 700700
rect 36892 700698 36916 700700
rect 36972 700698 36996 700700
rect 37052 700698 37076 700700
rect 37132 700698 37156 700700
rect 37212 700698 37236 700700
rect 37292 700698 37316 700700
rect 37372 700698 37386 700700
rect 37066 700646 37076 700698
rect 37132 700646 37142 700698
rect 36822 700644 36836 700646
rect 36892 700644 36916 700646
rect 36972 700644 36996 700646
rect 37052 700644 37076 700646
rect 37132 700644 37156 700646
rect 37212 700644 37236 700646
rect 37292 700644 37316 700646
rect 37372 700644 37386 700646
rect 36822 700624 37386 700644
rect 24306 700496 24362 700505
rect 24306 700431 24362 700440
rect 8114 700360 8170 700369
rect 72712 700330 72740 701950
rect 72822 701788 73386 701808
rect 72822 701786 72836 701788
rect 72892 701786 72916 701788
rect 72972 701786 72996 701788
rect 73052 701786 73076 701788
rect 73132 701786 73156 701788
rect 73212 701786 73236 701788
rect 73292 701786 73316 701788
rect 73372 701786 73386 701788
rect 73066 701734 73076 701786
rect 73132 701734 73142 701786
rect 72822 701732 72836 701734
rect 72892 701732 72916 701734
rect 72972 701732 72996 701734
rect 73052 701732 73076 701734
rect 73132 701732 73156 701734
rect 73212 701732 73236 701734
rect 73292 701732 73316 701734
rect 73372 701732 73386 701734
rect 72822 701712 73386 701732
rect 72822 700700 73386 700720
rect 72822 700698 72836 700700
rect 72892 700698 72916 700700
rect 72972 700698 72996 700700
rect 73052 700698 73076 700700
rect 73132 700698 73156 700700
rect 73212 700698 73236 700700
rect 73292 700698 73316 700700
rect 73372 700698 73386 700700
rect 73066 700646 73076 700698
rect 73132 700646 73142 700698
rect 72822 700644 72836 700646
rect 72892 700644 72916 700646
rect 72972 700644 72996 700646
rect 73052 700644 73076 700646
rect 73132 700644 73156 700646
rect 73212 700644 73236 700646
rect 73292 700644 73316 700646
rect 73372 700644 73386 700646
rect 72822 700624 73386 700644
rect 89180 700466 89208 703520
rect 90822 701244 91386 701264
rect 90822 701242 90836 701244
rect 90892 701242 90916 701244
rect 90972 701242 90996 701244
rect 91052 701242 91076 701244
rect 91132 701242 91156 701244
rect 91212 701242 91236 701244
rect 91292 701242 91316 701244
rect 91372 701242 91386 701244
rect 91066 701190 91076 701242
rect 91132 701190 91142 701242
rect 90822 701188 90836 701190
rect 90892 701188 90916 701190
rect 90972 701188 90996 701190
rect 91052 701188 91076 701190
rect 91132 701188 91156 701190
rect 91212 701188 91236 701190
rect 91292 701188 91316 701190
rect 91372 701188 91386 701190
rect 90822 701168 91386 701188
rect 105464 700806 105492 703520
rect 108822 701788 109386 701808
rect 108822 701786 108836 701788
rect 108892 701786 108916 701788
rect 108972 701786 108996 701788
rect 109052 701786 109076 701788
rect 109132 701786 109156 701788
rect 109212 701786 109236 701788
rect 109292 701786 109316 701788
rect 109372 701786 109386 701788
rect 109066 701734 109076 701786
rect 109132 701734 109142 701786
rect 108822 701732 108836 701734
rect 108892 701732 108916 701734
rect 108972 701732 108996 701734
rect 109052 701732 109076 701734
rect 109132 701732 109156 701734
rect 109212 701732 109236 701734
rect 109292 701732 109316 701734
rect 109372 701732 109386 701734
rect 108822 701712 109386 701732
rect 126822 701244 127386 701264
rect 126822 701242 126836 701244
rect 126892 701242 126916 701244
rect 126972 701242 126996 701244
rect 127052 701242 127076 701244
rect 127132 701242 127156 701244
rect 127212 701242 127236 701244
rect 127292 701242 127316 701244
rect 127372 701242 127386 701244
rect 127066 701190 127076 701242
rect 127132 701190 127142 701242
rect 126822 701188 126836 701190
rect 126892 701188 126916 701190
rect 126972 701188 126996 701190
rect 127052 701188 127076 701190
rect 127132 701188 127156 701190
rect 127212 701188 127236 701190
rect 127292 701188 127316 701190
rect 127372 701188 127386 701190
rect 126822 701168 127386 701188
rect 137848 700874 137876 703520
rect 144822 701788 145386 701808
rect 144822 701786 144836 701788
rect 144892 701786 144916 701788
rect 144972 701786 144996 701788
rect 145052 701786 145076 701788
rect 145132 701786 145156 701788
rect 145212 701786 145236 701788
rect 145292 701786 145316 701788
rect 145372 701786 145386 701788
rect 145066 701734 145076 701786
rect 145132 701734 145142 701786
rect 144822 701732 144836 701734
rect 144892 701732 144916 701734
rect 144972 701732 144996 701734
rect 145052 701732 145076 701734
rect 145132 701732 145156 701734
rect 145212 701732 145236 701734
rect 145292 701732 145316 701734
rect 145372 701732 145386 701734
rect 144822 701712 145386 701732
rect 154132 700942 154160 703520
rect 162822 701244 163386 701264
rect 162822 701242 162836 701244
rect 162892 701242 162916 701244
rect 162972 701242 162996 701244
rect 163052 701242 163076 701244
rect 163132 701242 163156 701244
rect 163212 701242 163236 701244
rect 163292 701242 163316 701244
rect 163372 701242 163386 701244
rect 163066 701190 163076 701242
rect 163132 701190 163142 701242
rect 162822 701188 162836 701190
rect 162892 701188 162916 701190
rect 162972 701188 162996 701190
rect 163052 701188 163076 701190
rect 163132 701188 163156 701190
rect 163212 701188 163236 701190
rect 163292 701188 163316 701190
rect 163372 701188 163386 701190
rect 162822 701168 163386 701188
rect 154120 700936 154172 700942
rect 154120 700878 154172 700884
rect 137836 700868 137888 700874
rect 137836 700810 137888 700816
rect 105452 700800 105504 700806
rect 105452 700742 105504 700748
rect 108822 700700 109386 700720
rect 108822 700698 108836 700700
rect 108892 700698 108916 700700
rect 108972 700698 108996 700700
rect 109052 700698 109076 700700
rect 109132 700698 109156 700700
rect 109212 700698 109236 700700
rect 109292 700698 109316 700700
rect 109372 700698 109386 700700
rect 109066 700646 109076 700698
rect 109132 700646 109142 700698
rect 108822 700644 108836 700646
rect 108892 700644 108916 700646
rect 108972 700644 108996 700646
rect 109052 700644 109076 700646
rect 109132 700644 109156 700646
rect 109212 700644 109236 700646
rect 109292 700644 109316 700646
rect 109372 700644 109386 700646
rect 108822 700624 109386 700644
rect 144822 700700 145386 700720
rect 144822 700698 144836 700700
rect 144892 700698 144916 700700
rect 144972 700698 144996 700700
rect 145052 700698 145076 700700
rect 145132 700698 145156 700700
rect 145212 700698 145236 700700
rect 145292 700698 145316 700700
rect 145372 700698 145386 700700
rect 145066 700646 145076 700698
rect 145132 700646 145142 700698
rect 144822 700644 144836 700646
rect 144892 700644 144916 700646
rect 144972 700644 144996 700646
rect 145052 700644 145076 700646
rect 145132 700644 145156 700646
rect 145212 700644 145236 700646
rect 145292 700644 145316 700646
rect 145372 700644 145386 700646
rect 144822 700624 145386 700644
rect 89168 700460 89220 700466
rect 89168 700402 89220 700408
rect 8114 700295 8170 700304
rect 72700 700324 72752 700330
rect 72700 700266 72752 700272
rect 18822 700156 19386 700176
rect 18822 700154 18836 700156
rect 18892 700154 18916 700156
rect 18972 700154 18996 700156
rect 19052 700154 19076 700156
rect 19132 700154 19156 700156
rect 19212 700154 19236 700156
rect 19292 700154 19316 700156
rect 19372 700154 19386 700156
rect 19066 700102 19076 700154
rect 19132 700102 19142 700154
rect 18822 700100 18836 700102
rect 18892 700100 18916 700102
rect 18972 700100 18996 700102
rect 19052 700100 19076 700102
rect 19132 700100 19156 700102
rect 19212 700100 19236 700102
rect 19292 700100 19316 700102
rect 19372 700100 19386 700102
rect 18822 700080 19386 700100
rect 54822 700156 55386 700176
rect 54822 700154 54836 700156
rect 54892 700154 54916 700156
rect 54972 700154 54996 700156
rect 55052 700154 55076 700156
rect 55132 700154 55156 700156
rect 55212 700154 55236 700156
rect 55292 700154 55316 700156
rect 55372 700154 55386 700156
rect 55066 700102 55076 700154
rect 55132 700102 55142 700154
rect 54822 700100 54836 700102
rect 54892 700100 54916 700102
rect 54972 700100 54996 700102
rect 55052 700100 55076 700102
rect 55132 700100 55156 700102
rect 55212 700100 55236 700102
rect 55292 700100 55316 700102
rect 55372 700100 55386 700102
rect 54822 700080 55386 700100
rect 90822 700156 91386 700176
rect 90822 700154 90836 700156
rect 90892 700154 90916 700156
rect 90972 700154 90996 700156
rect 91052 700154 91076 700156
rect 91132 700154 91156 700156
rect 91212 700154 91236 700156
rect 91292 700154 91316 700156
rect 91372 700154 91386 700156
rect 91066 700102 91076 700154
rect 91132 700102 91142 700154
rect 90822 700100 90836 700102
rect 90892 700100 90916 700102
rect 90972 700100 90996 700102
rect 91052 700100 91076 700102
rect 91132 700100 91156 700102
rect 91212 700100 91236 700102
rect 91292 700100 91316 700102
rect 91372 700100 91386 700102
rect 90822 700080 91386 700100
rect 126822 700156 127386 700176
rect 126822 700154 126836 700156
rect 126892 700154 126916 700156
rect 126972 700154 126996 700156
rect 127052 700154 127076 700156
rect 127132 700154 127156 700156
rect 127212 700154 127236 700156
rect 127292 700154 127316 700156
rect 127372 700154 127386 700156
rect 127066 700102 127076 700154
rect 127132 700102 127142 700154
rect 126822 700100 126836 700102
rect 126892 700100 126916 700102
rect 126972 700100 126996 700102
rect 127052 700100 127076 700102
rect 127132 700100 127156 700102
rect 127212 700100 127236 700102
rect 127292 700100 127316 700102
rect 127372 700100 127386 700102
rect 126822 700080 127386 700100
rect 162822 700156 163386 700176
rect 162822 700154 162836 700156
rect 162892 700154 162916 700156
rect 162972 700154 162996 700156
rect 163052 700154 163076 700156
rect 163132 700154 163156 700156
rect 163212 700154 163236 700156
rect 163292 700154 163316 700156
rect 163372 700154 163386 700156
rect 163066 700102 163076 700154
rect 163132 700102 163142 700154
rect 162822 700100 162836 700102
rect 162892 700100 162916 700102
rect 162972 700100 162996 700102
rect 163052 700100 163076 700102
rect 163132 700100 163156 700102
rect 163212 700100 163236 700102
rect 163292 700100 163316 700102
rect 163372 700100 163386 700102
rect 162822 700080 163386 700100
rect 170324 700058 170352 703520
rect 180822 701788 181386 701808
rect 180822 701786 180836 701788
rect 180892 701786 180916 701788
rect 180972 701786 180996 701788
rect 181052 701786 181076 701788
rect 181132 701786 181156 701788
rect 181212 701786 181236 701788
rect 181292 701786 181316 701788
rect 181372 701786 181386 701788
rect 181066 701734 181076 701786
rect 181132 701734 181142 701786
rect 180822 701732 180836 701734
rect 180892 701732 180916 701734
rect 180972 701732 180996 701734
rect 181052 701732 181076 701734
rect 181132 701732 181156 701734
rect 181212 701732 181236 701734
rect 181292 701732 181316 701734
rect 181372 701732 181386 701734
rect 180822 701712 181386 701732
rect 198822 701244 199386 701264
rect 198822 701242 198836 701244
rect 198892 701242 198916 701244
rect 198972 701242 198996 701244
rect 199052 701242 199076 701244
rect 199132 701242 199156 701244
rect 199212 701242 199236 701244
rect 199292 701242 199316 701244
rect 199372 701242 199386 701244
rect 199066 701190 199076 701242
rect 199132 701190 199142 701242
rect 198822 701188 198836 701190
rect 198892 701188 198916 701190
rect 198972 701188 198996 701190
rect 199052 701188 199076 701190
rect 199132 701188 199156 701190
rect 199212 701188 199236 701190
rect 199292 701188 199316 701190
rect 199372 701188 199386 701190
rect 198822 701168 199386 701188
rect 180822 700700 181386 700720
rect 180822 700698 180836 700700
rect 180892 700698 180916 700700
rect 180972 700698 180996 700700
rect 181052 700698 181076 700700
rect 181132 700698 181156 700700
rect 181212 700698 181236 700700
rect 181292 700698 181316 700700
rect 181372 700698 181386 700700
rect 181066 700646 181076 700698
rect 181132 700646 181142 700698
rect 180822 700644 180836 700646
rect 180892 700644 180916 700646
rect 180972 700644 180996 700646
rect 181052 700644 181076 700646
rect 181132 700644 181156 700646
rect 181212 700644 181236 700646
rect 181292 700644 181316 700646
rect 181372 700644 181386 700646
rect 180822 700624 181386 700644
rect 202800 700398 202828 703520
rect 216822 701788 217386 701808
rect 216822 701786 216836 701788
rect 216892 701786 216916 701788
rect 216972 701786 216996 701788
rect 217052 701786 217076 701788
rect 217132 701786 217156 701788
rect 217212 701786 217236 701788
rect 217292 701786 217316 701788
rect 217372 701786 217386 701788
rect 217066 701734 217076 701786
rect 217132 701734 217142 701786
rect 216822 701732 216836 701734
rect 216892 701732 216916 701734
rect 216972 701732 216996 701734
rect 217052 701732 217076 701734
rect 217132 701732 217156 701734
rect 217212 701732 217236 701734
rect 217292 701732 217316 701734
rect 217372 701732 217386 701734
rect 216822 701712 217386 701732
rect 216822 700700 217386 700720
rect 216822 700698 216836 700700
rect 216892 700698 216916 700700
rect 216972 700698 216996 700700
rect 217052 700698 217076 700700
rect 217132 700698 217156 700700
rect 217212 700698 217236 700700
rect 217292 700698 217316 700700
rect 217372 700698 217386 700700
rect 217066 700646 217076 700698
rect 217132 700646 217142 700698
rect 216822 700644 216836 700646
rect 216892 700644 216916 700646
rect 216972 700644 216996 700646
rect 217052 700644 217076 700646
rect 217132 700644 217156 700646
rect 217212 700644 217236 700646
rect 217292 700644 217316 700646
rect 217372 700644 217386 700646
rect 216822 700624 217386 700644
rect 202788 700392 202840 700398
rect 202788 700334 202840 700340
rect 198822 700156 199386 700176
rect 198822 700154 198836 700156
rect 198892 700154 198916 700156
rect 198972 700154 198996 700156
rect 199052 700154 199076 700156
rect 199132 700154 199156 700156
rect 199212 700154 199236 700156
rect 199292 700154 199316 700156
rect 199372 700154 199386 700156
rect 199066 700102 199076 700154
rect 199132 700102 199142 700154
rect 198822 700100 198836 700102
rect 198892 700100 198916 700102
rect 198972 700100 198996 700102
rect 199052 700100 199076 700102
rect 199132 700100 199156 700102
rect 199212 700100 199236 700102
rect 199292 700100 199316 700102
rect 199372 700100 199386 700102
rect 198822 700080 199386 700100
rect 170312 700052 170364 700058
rect 170312 699994 170364 700000
rect 218992 699922 219020 703520
rect 223304 701888 223356 701894
rect 223304 701830 223356 701836
rect 218980 699916 219032 699922
rect 218980 699858 219032 699864
rect 36822 699612 37386 699632
rect 36822 699610 36836 699612
rect 36892 699610 36916 699612
rect 36972 699610 36996 699612
rect 37052 699610 37076 699612
rect 37132 699610 37156 699612
rect 37212 699610 37236 699612
rect 37292 699610 37316 699612
rect 37372 699610 37386 699612
rect 37066 699558 37076 699610
rect 37132 699558 37142 699610
rect 36822 699556 36836 699558
rect 36892 699556 36916 699558
rect 36972 699556 36996 699558
rect 37052 699556 37076 699558
rect 37132 699556 37156 699558
rect 37212 699556 37236 699558
rect 37292 699556 37316 699558
rect 37372 699556 37386 699558
rect 36822 699536 37386 699556
rect 72822 699612 73386 699632
rect 72822 699610 72836 699612
rect 72892 699610 72916 699612
rect 72972 699610 72996 699612
rect 73052 699610 73076 699612
rect 73132 699610 73156 699612
rect 73212 699610 73236 699612
rect 73292 699610 73316 699612
rect 73372 699610 73386 699612
rect 73066 699558 73076 699610
rect 73132 699558 73142 699610
rect 72822 699556 72836 699558
rect 72892 699556 72916 699558
rect 72972 699556 72996 699558
rect 73052 699556 73076 699558
rect 73132 699556 73156 699558
rect 73212 699556 73236 699558
rect 73292 699556 73316 699558
rect 73372 699556 73386 699558
rect 72822 699536 73386 699556
rect 108822 699612 109386 699632
rect 108822 699610 108836 699612
rect 108892 699610 108916 699612
rect 108972 699610 108996 699612
rect 109052 699610 109076 699612
rect 109132 699610 109156 699612
rect 109212 699610 109236 699612
rect 109292 699610 109316 699612
rect 109372 699610 109386 699612
rect 109066 699558 109076 699610
rect 109132 699558 109142 699610
rect 108822 699556 108836 699558
rect 108892 699556 108916 699558
rect 108972 699556 108996 699558
rect 109052 699556 109076 699558
rect 109132 699556 109156 699558
rect 109212 699556 109236 699558
rect 109292 699556 109316 699558
rect 109372 699556 109386 699558
rect 108822 699536 109386 699556
rect 144822 699612 145386 699632
rect 144822 699610 144836 699612
rect 144892 699610 144916 699612
rect 144972 699610 144996 699612
rect 145052 699610 145076 699612
rect 145132 699610 145156 699612
rect 145212 699610 145236 699612
rect 145292 699610 145316 699612
rect 145372 699610 145386 699612
rect 145066 699558 145076 699610
rect 145132 699558 145142 699610
rect 144822 699556 144836 699558
rect 144892 699556 144916 699558
rect 144972 699556 144996 699558
rect 145052 699556 145076 699558
rect 145132 699556 145156 699558
rect 145212 699556 145236 699558
rect 145292 699556 145316 699558
rect 145372 699556 145386 699558
rect 144822 699536 145386 699556
rect 180822 699612 181386 699632
rect 180822 699610 180836 699612
rect 180892 699610 180916 699612
rect 180972 699610 180996 699612
rect 181052 699610 181076 699612
rect 181132 699610 181156 699612
rect 181212 699610 181236 699612
rect 181292 699610 181316 699612
rect 181372 699610 181386 699612
rect 181066 699558 181076 699610
rect 181132 699558 181142 699610
rect 180822 699556 180836 699558
rect 180892 699556 180916 699558
rect 180972 699556 180996 699558
rect 181052 699556 181076 699558
rect 181132 699556 181156 699558
rect 181212 699556 181236 699558
rect 181292 699556 181316 699558
rect 181372 699556 181386 699558
rect 180822 699536 181386 699556
rect 216822 699612 217386 699632
rect 216822 699610 216836 699612
rect 216892 699610 216916 699612
rect 216972 699610 216996 699612
rect 217052 699610 217076 699612
rect 217132 699610 217156 699612
rect 217212 699610 217236 699612
rect 217292 699610 217316 699612
rect 217372 699610 217386 699612
rect 217066 699558 217076 699610
rect 217132 699558 217142 699610
rect 216822 699556 216836 699558
rect 216892 699556 216916 699558
rect 216972 699556 216996 699558
rect 217052 699556 217076 699558
rect 217132 699556 217156 699558
rect 217212 699556 217236 699558
rect 217292 699556 217316 699558
rect 217372 699556 217386 699558
rect 216822 699536 217386 699556
rect 142804 699508 142856 699514
rect 142804 699450 142856 699456
rect 71780 699440 71832 699446
rect 71780 699382 71832 699388
rect 48136 699236 48188 699242
rect 48136 699178 48188 699184
rect 5080 699168 5132 699174
rect 5080 699110 5132 699116
rect 4802 698864 4858 698873
rect 4802 698799 4858 698808
rect 4068 696720 4120 696726
rect 4068 696662 4120 696668
rect 3148 696516 3200 696522
rect 3148 696458 3200 696464
rect 2964 682576 3016 682582
rect 2964 682518 3016 682524
rect 2976 682281 3004 682518
rect 2962 682272 3018 682281
rect 2962 682207 3018 682216
rect 2780 668228 2832 668234
rect 2780 668170 2832 668176
rect 2792 668001 2820 668170
rect 2778 667992 2834 668001
rect 2778 667927 2834 667936
rect 3056 654016 3108 654022
rect 3056 653958 3108 653964
rect 3068 653585 3096 653958
rect 3054 653576 3110 653585
rect 3054 653511 3110 653520
rect 2964 624912 3016 624918
rect 2962 624880 2964 624889
rect 3016 624880 3018 624889
rect 2962 624815 3018 624824
rect 3160 610473 3188 696458
rect 3884 696244 3936 696250
rect 3884 696186 3936 696192
rect 3332 696176 3384 696182
rect 3332 696118 3384 696124
rect 3240 695360 3292 695366
rect 3240 695302 3292 695308
rect 3146 610464 3202 610473
rect 3146 610399 3202 610408
rect 3148 596080 3200 596086
rect 3146 596048 3148 596057
rect 3200 596048 3202 596057
rect 3146 595983 3202 595992
rect 3056 567656 3108 567662
rect 3056 567598 3108 567604
rect 3068 567361 3096 567598
rect 3054 567352 3110 567361
rect 3054 567287 3110 567296
rect 3252 538665 3280 695302
rect 3238 538656 3294 538665
rect 3238 538591 3294 538600
rect 3056 510400 3108 510406
rect 3056 510342 3108 510348
rect 3068 509969 3096 510342
rect 3054 509960 3110 509969
rect 3054 509895 3110 509904
rect 3344 495553 3372 696118
rect 3792 695904 3844 695910
rect 3792 695846 3844 695852
rect 3516 695564 3568 695570
rect 3516 695506 3568 695512
rect 3422 693832 3478 693841
rect 3422 693767 3478 693776
rect 3330 495544 3386 495553
rect 3330 495479 3386 495488
rect 3332 481160 3384 481166
rect 3330 481128 3332 481137
rect 3384 481128 3386 481137
rect 3330 481063 3386 481072
rect 3332 452464 3384 452470
rect 3330 452432 3332 452441
rect 3384 452432 3386 452441
rect 3330 452367 3386 452376
rect 3332 438932 3384 438938
rect 3332 438874 3384 438880
rect 2872 423904 2924 423910
rect 2872 423846 2924 423852
rect 2884 423745 2912 423846
rect 2870 423736 2926 423745
rect 2870 423671 2926 423680
rect 3240 395752 3292 395758
rect 3240 395694 3292 395700
rect 3252 395049 3280 395694
rect 3238 395040 3294 395049
rect 3238 394975 3294 394984
rect 2780 380656 2832 380662
rect 2778 380624 2780 380633
rect 2832 380624 2834 380633
rect 2778 380559 2834 380568
rect 3240 367056 3292 367062
rect 3240 366998 3292 367004
rect 3252 366217 3280 366998
rect 3238 366208 3294 366217
rect 3238 366143 3294 366152
rect 3240 337680 3292 337686
rect 3240 337622 3292 337628
rect 3252 337521 3280 337622
rect 3238 337512 3294 337521
rect 3238 337447 3294 337456
rect 3240 308916 3292 308922
rect 3240 308858 3292 308864
rect 3252 308825 3280 308858
rect 3238 308816 3294 308825
rect 3238 308751 3294 308760
rect 3240 294772 3292 294778
rect 3240 294714 3292 294720
rect 3252 294409 3280 294714
rect 3238 294400 3294 294409
rect 3238 294335 3294 294344
rect 2778 280120 2834 280129
rect 2778 280055 2780 280064
rect 2832 280055 2834 280064
rect 2780 280026 2832 280032
rect 2964 266348 3016 266354
rect 2964 266290 3016 266296
rect 2976 265713 3004 266290
rect 2962 265704 3018 265713
rect 2962 265639 3018 265648
rect 3240 252544 3292 252550
rect 3240 252486 3292 252492
rect 3252 251297 3280 252486
rect 3238 251288 3294 251297
rect 3238 251223 3294 251232
rect 3344 237017 3372 438874
rect 3330 237008 3386 237017
rect 3330 236943 3386 236952
rect 3332 208208 3384 208214
rect 3330 208176 3332 208185
rect 3384 208176 3386 208185
rect 3330 208111 3386 208120
rect 2780 194472 2832 194478
rect 2780 194414 2832 194420
rect 2792 193905 2820 194414
rect 2778 193896 2834 193905
rect 2778 193831 2834 193840
rect 3332 165096 3384 165102
rect 3330 165064 3332 165073
rect 3384 165064 3386 165073
rect 3330 164999 3386 165008
rect 3332 136400 3384 136406
rect 3330 136368 3332 136377
rect 3384 136368 3386 136377
rect 3330 136303 3386 136312
rect 3332 122188 3384 122194
rect 3332 122130 3384 122136
rect 3344 122097 3372 122130
rect 3330 122088 3386 122097
rect 3330 122023 3386 122032
rect 2780 108044 2832 108050
rect 2780 107986 2832 107992
rect 2792 107681 2820 107986
rect 2778 107672 2834 107681
rect 2778 107607 2834 107616
rect 3056 79892 3108 79898
rect 3056 79834 3108 79840
rect 3068 78985 3096 79834
rect 3054 78976 3110 78985
rect 3054 78911 3110 78920
rect 3436 50153 3464 693767
rect 3528 64569 3556 695506
rect 3700 694612 3752 694618
rect 3700 694554 3752 694560
rect 3608 694340 3660 694346
rect 3608 694282 3660 694288
rect 3620 93265 3648 694282
rect 3712 179489 3740 694554
rect 3804 222601 3832 695846
rect 3896 553081 3924 696186
rect 3976 695088 4028 695094
rect 3976 695030 4028 695036
rect 3882 553072 3938 553081
rect 3882 553007 3938 553016
rect 3884 539436 3936 539442
rect 3884 539378 3936 539384
rect 3790 222592 3846 222601
rect 3790 222527 3846 222536
rect 3698 179480 3754 179489
rect 3698 179415 3754 179424
rect 3896 150793 3924 539378
rect 3988 323105 4016 695030
rect 4080 438025 4108 696662
rect 4066 438016 4122 438025
rect 4066 437951 4122 437960
rect 3974 323096 4030 323105
rect 3974 323031 4030 323040
rect 3882 150784 3938 150793
rect 3882 150719 3938 150728
rect 3606 93256 3662 93265
rect 3606 93191 3662 93200
rect 3514 64560 3570 64569
rect 3514 64495 3570 64504
rect 3422 50144 3478 50153
rect 3422 50079 3478 50088
rect 3422 35864 3478 35873
rect 3422 35799 3424 35808
rect 3476 35799 3478 35808
rect 3424 35770 3476 35776
rect 4816 21894 4844 698799
rect 4986 698728 5042 698737
rect 4986 698663 5042 698672
rect 4896 695700 4948 695706
rect 4896 695642 4948 695648
rect 4908 194478 4936 695642
rect 4896 194472 4948 194478
rect 4896 194414 4948 194420
rect 5000 108050 5028 698663
rect 5092 280090 5120 699110
rect 18822 699068 19386 699088
rect 18822 699066 18836 699068
rect 18892 699066 18916 699068
rect 18972 699066 18996 699068
rect 19052 699066 19076 699068
rect 19132 699066 19156 699068
rect 19212 699066 19236 699068
rect 19292 699066 19316 699068
rect 19372 699066 19386 699068
rect 19066 699014 19076 699066
rect 19132 699014 19142 699066
rect 18822 699012 18836 699014
rect 18892 699012 18916 699014
rect 18972 699012 18996 699014
rect 19052 699012 19076 699014
rect 19132 699012 19156 699014
rect 19212 699012 19236 699014
rect 19292 699012 19316 699014
rect 19372 699012 19386 699014
rect 18822 698992 19386 699012
rect 5264 698828 5316 698834
rect 5264 698770 5316 698776
rect 5172 696040 5224 696046
rect 5172 695982 5224 695988
rect 5184 380662 5212 695982
rect 5276 438938 5304 698770
rect 33968 698760 34020 698766
rect 33968 698702 34020 698708
rect 5356 698624 5408 698630
rect 5356 698566 5408 698572
rect 5368 539442 5396 698566
rect 5816 698284 5868 698290
rect 5816 698226 5868 698232
rect 5448 696652 5500 696658
rect 5448 696594 5500 696600
rect 5460 668234 5488 696594
rect 5828 682582 5856 698226
rect 5908 698216 5960 698222
rect 5908 698158 5960 698164
rect 5816 682576 5868 682582
rect 5816 682518 5868 682524
rect 5448 668228 5500 668234
rect 5448 668170 5500 668176
rect 5920 624918 5948 698158
rect 6012 698018 6132 698034
rect 6012 698012 6144 698018
rect 6012 698006 6092 698012
rect 5908 624912 5960 624918
rect 5908 624854 5960 624860
rect 6012 567662 6040 698006
rect 6092 697954 6144 697960
rect 6092 697876 6144 697882
rect 6092 697818 6144 697824
rect 6000 567656 6052 567662
rect 6000 567598 6052 567604
rect 5356 539436 5408 539442
rect 5356 539378 5408 539384
rect 6104 510406 6132 697818
rect 7472 697808 7524 697814
rect 7472 697750 7524 697756
rect 6828 697672 6880 697678
rect 6828 697614 6880 697620
rect 6736 697536 6788 697542
rect 6736 697478 6788 697484
rect 6552 697400 6604 697406
rect 6552 697342 6604 697348
rect 6368 697332 6420 697338
rect 6368 697274 6420 697280
rect 6276 697264 6328 697270
rect 6276 697206 6328 697212
rect 6182 697096 6238 697105
rect 6182 697031 6238 697040
rect 6092 510400 6144 510406
rect 6092 510342 6144 510348
rect 5264 438932 5316 438938
rect 5264 438874 5316 438880
rect 5172 380656 5224 380662
rect 5172 380598 5224 380604
rect 5080 280084 5132 280090
rect 5080 280026 5132 280032
rect 4988 108044 5040 108050
rect 4988 107986 5040 107992
rect 2780 21888 2832 21894
rect 2780 21830 2832 21836
rect 4804 21888 4856 21894
rect 4804 21830 4856 21836
rect 2792 21457 2820 21830
rect 2778 21448 2834 21457
rect 2778 21383 2834 21392
rect 6196 7206 6224 697031
rect 6288 252550 6316 697206
rect 6380 266354 6408 697274
rect 6460 695972 6512 695978
rect 6460 695914 6512 695920
rect 6472 294778 6500 695914
rect 6564 337686 6592 697342
rect 6642 694104 6698 694113
rect 6642 694039 6698 694048
rect 6656 367062 6684 694039
rect 6748 395758 6776 697478
rect 6840 452470 6868 697614
rect 7288 695496 7340 695502
rect 7288 695438 7340 695444
rect 7300 654022 7328 695438
rect 7380 695428 7432 695434
rect 7380 695370 7432 695376
rect 7288 654016 7340 654022
rect 7288 653958 7340 653964
rect 7392 596086 7420 695370
rect 7380 596080 7432 596086
rect 7380 596022 7432 596028
rect 7484 481166 7512 697750
rect 7932 697196 7984 697202
rect 7932 697138 7984 697144
rect 7564 697128 7616 697134
rect 7564 697070 7616 697076
rect 7472 481160 7524 481166
rect 7472 481102 7524 481108
rect 6828 452464 6880 452470
rect 6828 452406 6880 452412
rect 6736 395752 6788 395758
rect 6736 395694 6788 395700
rect 6644 367056 6696 367062
rect 6644 366998 6696 367004
rect 6552 337680 6604 337686
rect 6552 337622 6604 337628
rect 6460 294772 6512 294778
rect 6460 294714 6512 294720
rect 6368 266348 6420 266354
rect 6368 266290 6420 266296
rect 6276 252544 6328 252550
rect 6276 252486 6328 252492
rect 7576 35834 7604 697070
rect 7748 695700 7800 695706
rect 7748 695642 7800 695648
rect 7654 693696 7710 693705
rect 7654 693631 7710 693640
rect 7668 79898 7696 693631
rect 7760 122194 7788 695642
rect 7840 694612 7892 694618
rect 7840 694554 7892 694560
rect 7852 136406 7880 694554
rect 7944 165102 7972 697138
rect 24492 696992 24544 696998
rect 10322 696960 10378 696969
rect 24492 696934 24544 696940
rect 10322 696895 10378 696904
rect 8208 696108 8260 696114
rect 8208 696050 8260 696056
rect 8024 695836 8076 695842
rect 8024 695778 8076 695784
rect 8036 208214 8064 695778
rect 8116 695088 8168 695094
rect 8116 695030 8168 695036
rect 8128 308922 8156 695030
rect 8220 423910 8248 696050
rect 10336 695980 10364 696895
rect 19982 696008 20038 696017
rect 19734 695966 19982 695994
rect 24504 695980 24532 696934
rect 33980 695980 34008 698702
rect 36822 698524 37386 698544
rect 36822 698522 36836 698524
rect 36892 698522 36916 698524
rect 36972 698522 36996 698524
rect 37052 698522 37076 698524
rect 37132 698522 37156 698524
rect 37212 698522 37236 698524
rect 37292 698522 37316 698524
rect 37372 698522 37386 698524
rect 37066 698470 37076 698522
rect 37132 698470 37142 698522
rect 36822 698468 36836 698470
rect 36892 698468 36916 698470
rect 36972 698468 36996 698470
rect 37052 698468 37076 698470
rect 37132 698468 37156 698470
rect 37212 698468 37236 698470
rect 37292 698468 37316 698470
rect 37372 698468 37386 698470
rect 36822 698448 37386 698468
rect 38660 697060 38712 697066
rect 38660 697002 38712 697008
rect 38672 695980 38700 697002
rect 48148 695980 48176 699178
rect 54822 699068 55386 699088
rect 54822 699066 54836 699068
rect 54892 699066 54916 699068
rect 54972 699066 54996 699068
rect 55052 699066 55076 699068
rect 55132 699066 55156 699068
rect 55212 699066 55236 699068
rect 55292 699066 55316 699068
rect 55372 699066 55386 699068
rect 55066 699014 55076 699066
rect 55132 699014 55142 699066
rect 54822 699012 54836 699014
rect 54892 699012 54916 699014
rect 54972 699012 54996 699014
rect 55052 699012 55076 699014
rect 55132 699012 55156 699014
rect 55212 699012 55236 699014
rect 55292 699012 55316 699014
rect 55372 699012 55386 699014
rect 54822 698992 55386 699012
rect 57612 698896 57664 698902
rect 57612 698838 57664 698844
rect 57624 695980 57652 698838
rect 62304 698352 62356 698358
rect 62304 698294 62356 698300
rect 62316 695980 62344 698294
rect 71792 695980 71820 699382
rect 100208 699372 100260 699378
rect 100208 699314 100260 699320
rect 90822 699068 91386 699088
rect 90822 699066 90836 699068
rect 90892 699066 90916 699068
rect 90972 699066 90996 699068
rect 91052 699066 91076 699068
rect 91132 699066 91156 699068
rect 91212 699066 91236 699068
rect 91292 699066 91316 699068
rect 91372 699066 91386 699068
rect 91066 699014 91076 699066
rect 91132 699014 91142 699066
rect 90822 699012 90836 699014
rect 90892 699012 90916 699014
rect 90972 699012 90996 699014
rect 91052 699012 91076 699014
rect 91132 699012 91156 699014
rect 91212 699012 91236 699014
rect 91292 699012 91316 699014
rect 91372 699012 91386 699014
rect 90822 698992 91386 699012
rect 89720 698760 89772 698766
rect 89720 698702 89772 698708
rect 72822 698524 73386 698544
rect 72822 698522 72836 698524
rect 72892 698522 72916 698524
rect 72972 698522 72996 698524
rect 73052 698522 73076 698524
rect 73132 698522 73156 698524
rect 73212 698522 73236 698524
rect 73292 698522 73316 698524
rect 73372 698522 73386 698524
rect 73066 698470 73076 698522
rect 73132 698470 73142 698522
rect 72822 698468 72836 698470
rect 72892 698468 72916 698470
rect 72972 698468 72996 698470
rect 73052 698468 73076 698470
rect 73132 698468 73156 698470
rect 73212 698468 73236 698470
rect 73292 698468 73316 698470
rect 73372 698468 73386 698470
rect 72822 698448 73386 698468
rect 76564 698420 76616 698426
rect 76564 698362 76616 698368
rect 76576 695980 76604 698362
rect 81256 696244 81308 696250
rect 81256 696186 81308 696192
rect 81268 695980 81296 696186
rect 89732 696153 89760 698702
rect 90732 698692 90784 698698
rect 90732 698634 90784 698640
rect 89718 696144 89774 696153
rect 89718 696079 89774 696088
rect 90744 695980 90772 698634
rect 100220 695980 100248 699314
rect 133328 699304 133380 699310
rect 133328 699246 133380 699252
rect 126822 699068 127386 699088
rect 126822 699066 126836 699068
rect 126892 699066 126916 699068
rect 126972 699066 126996 699068
rect 127052 699066 127076 699068
rect 127132 699066 127156 699068
rect 127212 699066 127236 699068
rect 127292 699066 127316 699068
rect 127372 699066 127386 699068
rect 127066 699014 127076 699066
rect 127132 699014 127142 699066
rect 126822 699012 126836 699014
rect 126892 699012 126916 699014
rect 126972 699012 126996 699014
rect 127052 699012 127076 699014
rect 127132 699012 127156 699014
rect 127212 699012 127236 699014
rect 127292 699012 127316 699014
rect 127372 699012 127386 699014
rect 126822 698992 127386 699012
rect 119160 698964 119212 698970
rect 119160 698906 119212 698912
rect 107568 698896 107620 698902
rect 107568 698838 107620 698844
rect 114376 698896 114428 698902
rect 114376 698838 114428 698844
rect 104992 698760 105044 698766
rect 104992 698702 105044 698708
rect 105004 695980 105032 698702
rect 107580 696250 107608 698838
rect 108822 698524 109386 698544
rect 108822 698522 108836 698524
rect 108892 698522 108916 698524
rect 108972 698522 108996 698524
rect 109052 698522 109076 698524
rect 109132 698522 109156 698524
rect 109212 698522 109236 698524
rect 109292 698522 109316 698524
rect 109372 698522 109386 698524
rect 109066 698470 109076 698522
rect 109132 698470 109142 698522
rect 108822 698468 108836 698470
rect 108892 698468 108916 698470
rect 108972 698468 108996 698470
rect 109052 698468 109076 698470
rect 109132 698468 109156 698470
rect 109212 698468 109236 698470
rect 109292 698468 109316 698470
rect 109372 698468 109386 698470
rect 108822 698448 109386 698468
rect 107568 696244 107620 696250
rect 107568 696186 107620 696192
rect 114388 695980 114416 698838
rect 119172 695980 119200 698906
rect 133340 695980 133368 699246
rect 142712 699236 142764 699242
rect 142712 699178 142764 699184
rect 142724 696590 142752 699178
rect 142712 696584 142764 696590
rect 142712 696526 142764 696532
rect 142816 695980 142844 699450
rect 146944 699304 146996 699310
rect 146944 699246 146996 699252
rect 161756 699304 161808 699310
rect 161756 699246 161808 699252
rect 186134 699272 186190 699281
rect 144822 698524 145386 698544
rect 144822 698522 144836 698524
rect 144892 698522 144916 698524
rect 144972 698522 144996 698524
rect 145052 698522 145076 698524
rect 145132 698522 145156 698524
rect 145212 698522 145236 698524
rect 145292 698522 145316 698524
rect 145372 698522 145386 698524
rect 145066 698470 145076 698522
rect 145132 698470 145142 698522
rect 144822 698468 144836 698470
rect 144892 698468 144916 698470
rect 144972 698468 144996 698470
rect 145052 698468 145076 698470
rect 145132 698468 145156 698470
rect 145212 698468 145236 698470
rect 145292 698468 145316 698470
rect 145372 698468 145386 698470
rect 144822 698448 145386 698468
rect 146956 696658 146984 699246
rect 147588 699236 147640 699242
rect 147588 699178 147640 699184
rect 146944 696652 146996 696658
rect 146944 696594 146996 696600
rect 147600 695980 147628 699178
rect 152280 697468 152332 697474
rect 152280 697410 152332 697416
rect 152292 695980 152320 697410
rect 160100 696788 160152 696794
rect 160100 696730 160152 696736
rect 160192 696788 160244 696794
rect 160192 696730 160244 696736
rect 160112 696674 160140 696730
rect 160204 696674 160232 696730
rect 160112 696646 160232 696674
rect 161768 695980 161796 699246
rect 186134 699207 186136 699216
rect 186188 699207 186190 699216
rect 186136 699178 186188 699184
rect 162822 699068 163386 699088
rect 162822 699066 162836 699068
rect 162892 699066 162916 699068
rect 162972 699066 162996 699068
rect 163052 699066 163076 699068
rect 163132 699066 163156 699068
rect 163212 699066 163236 699068
rect 163292 699066 163316 699068
rect 163372 699066 163386 699068
rect 163066 699014 163076 699066
rect 163132 699014 163142 699066
rect 162822 699012 162836 699014
rect 162892 699012 162916 699014
rect 162972 699012 162996 699014
rect 163052 699012 163076 699014
rect 163132 699012 163156 699014
rect 163212 699012 163236 699014
rect 163292 699012 163316 699014
rect 163372 699012 163386 699014
rect 162822 698992 163386 699012
rect 198822 699068 199386 699088
rect 198822 699066 198836 699068
rect 198892 699066 198916 699068
rect 198972 699066 198996 699068
rect 199052 699066 199076 699068
rect 199132 699066 199156 699068
rect 199212 699066 199236 699068
rect 199292 699066 199316 699068
rect 199372 699066 199386 699068
rect 199066 699014 199076 699066
rect 199132 699014 199142 699066
rect 198822 699012 198836 699014
rect 198892 699012 198916 699014
rect 198972 699012 198996 699014
rect 199052 699012 199076 699014
rect 199132 699012 199156 699014
rect 199212 699012 199236 699014
rect 199292 699012 199316 699014
rect 199372 699012 199386 699014
rect 198822 698992 199386 699012
rect 180822 698524 181386 698544
rect 180822 698522 180836 698524
rect 180892 698522 180916 698524
rect 180972 698522 180996 698524
rect 181052 698522 181076 698524
rect 181132 698522 181156 698524
rect 181212 698522 181236 698524
rect 181292 698522 181316 698524
rect 181372 698522 181386 698524
rect 181066 698470 181076 698522
rect 181132 698470 181142 698522
rect 180822 698468 180836 698470
rect 180892 698468 180916 698470
rect 180972 698468 180996 698470
rect 181052 698468 181076 698470
rect 181132 698468 181156 698470
rect 181212 698468 181236 698470
rect 181292 698468 181316 698470
rect 181372 698468 181386 698470
rect 180822 698448 181386 698468
rect 216822 698524 217386 698544
rect 216822 698522 216836 698524
rect 216892 698522 216916 698524
rect 216972 698522 216996 698524
rect 217052 698522 217076 698524
rect 217132 698522 217156 698524
rect 217212 698522 217236 698524
rect 217292 698522 217316 698524
rect 217372 698522 217386 698524
rect 217066 698470 217076 698522
rect 217132 698470 217142 698522
rect 216822 698468 216836 698470
rect 216892 698468 216916 698470
rect 216972 698468 216996 698470
rect 217052 698468 217076 698470
rect 217132 698468 217156 698470
rect 217212 698468 217236 698470
rect 217292 698468 217316 698470
rect 217372 698468 217386 698470
rect 216822 698448 217386 698468
rect 218058 698456 218114 698465
rect 218058 698391 218060 698400
rect 218112 698391 218114 698400
rect 218426 698456 218482 698465
rect 218426 698391 218428 698400
rect 218060 698362 218112 698368
rect 218480 698391 218482 698400
rect 218428 698362 218480 698368
rect 218058 698320 218114 698329
rect 218058 698255 218060 698264
rect 218112 698255 218114 698264
rect 218426 698320 218482 698329
rect 218426 698255 218428 698264
rect 218060 698226 218112 698232
rect 218480 698255 218482 698264
rect 218428 698226 218480 698232
rect 215116 698216 215168 698222
rect 208950 698184 209006 698193
rect 193312 698148 193364 698154
rect 193312 698090 193364 698096
rect 202788 698148 202840 698154
rect 215114 698184 215116 698193
rect 218152 698216 218204 698222
rect 215168 698184 215170 698193
rect 208950 698119 208952 698128
rect 202788 698090 202840 698096
rect 209004 698119 209006 698128
rect 209044 698148 209096 698154
rect 208952 698090 209004 698096
rect 218336 698216 218388 698222
rect 218204 698164 218336 698170
rect 218152 698158 218388 698164
rect 218164 698142 218376 698158
rect 215114 698119 215170 698128
rect 209044 698090 209096 698096
rect 193324 698057 193352 698090
rect 202800 698057 202828 698090
rect 193310 698048 193366 698057
rect 193310 697983 193366 697992
rect 202786 698048 202842 698057
rect 202786 697983 202842 697992
rect 194876 697944 194928 697950
rect 194876 697886 194928 697892
rect 180708 697740 180760 697746
rect 180708 697682 180760 697688
rect 166448 697604 166500 697610
rect 166448 697546 166500 697552
rect 165528 696448 165580 696454
rect 165528 696390 165580 696396
rect 165712 696448 165764 696454
rect 165712 696390 165764 696396
rect 165540 696266 165568 696390
rect 165724 696266 165752 696390
rect 165540 696238 165752 696266
rect 166460 695980 166488 697546
rect 180720 695980 180748 697682
rect 190184 696312 190236 696318
rect 190184 696254 190236 696260
rect 190196 695980 190224 696254
rect 194888 695980 194916 697886
rect 204352 696448 204404 696454
rect 204352 696390 204404 696396
rect 204364 695980 204392 696390
rect 205546 696008 205602 696017
rect 19982 695943 20038 695952
rect 209056 695980 209084 698090
rect 213828 698080 213880 698086
rect 213828 698022 213880 698028
rect 213734 696008 213790 696017
rect 205546 695943 205602 695952
rect 213840 695980 213868 698022
rect 218520 696720 218572 696726
rect 218520 696662 218572 696668
rect 218532 695980 218560 696662
rect 223316 695980 223344 701830
rect 235184 701690 235212 703520
rect 251640 702024 251692 702030
rect 251640 701966 251692 701972
rect 237472 701956 237524 701962
rect 237472 701898 237524 701904
rect 235172 701684 235224 701690
rect 235172 701626 235224 701632
rect 234822 701244 235386 701264
rect 234822 701242 234836 701244
rect 234892 701242 234916 701244
rect 234972 701242 234996 701244
rect 235052 701242 235076 701244
rect 235132 701242 235156 701244
rect 235212 701242 235236 701244
rect 235292 701242 235316 701244
rect 235372 701242 235386 701244
rect 235066 701190 235076 701242
rect 235132 701190 235142 701242
rect 234822 701188 234836 701190
rect 234892 701188 234916 701190
rect 234972 701188 234996 701190
rect 235052 701188 235076 701190
rect 235132 701188 235156 701190
rect 235212 701188 235236 701190
rect 235292 701188 235316 701190
rect 235372 701188 235386 701190
rect 234822 701168 235386 701188
rect 227994 700904 228050 700913
rect 227994 700839 228050 700848
rect 226338 698320 226394 698329
rect 226338 698255 226394 698264
rect 226352 698222 226380 698255
rect 226340 698216 226392 698222
rect 226340 698158 226392 698164
rect 224958 696416 225014 696425
rect 224958 696351 224960 696360
rect 225012 696351 225014 696360
rect 224960 696322 225012 696328
rect 228008 695980 228036 700839
rect 234822 700156 235386 700176
rect 234822 700154 234836 700156
rect 234892 700154 234916 700156
rect 234972 700154 234996 700156
rect 235052 700154 235076 700156
rect 235132 700154 235156 700156
rect 235212 700154 235236 700156
rect 235292 700154 235316 700156
rect 235372 700154 235386 700156
rect 235066 700102 235076 700154
rect 235132 700102 235142 700154
rect 234822 700100 234836 700102
rect 234892 700100 234916 700102
rect 234972 700100 234996 700102
rect 235052 700100 235076 700102
rect 235132 700100 235156 700102
rect 235212 700100 235236 700102
rect 235292 700100 235316 700102
rect 235372 700100 235386 700102
rect 234822 700080 235386 700100
rect 234822 699068 235386 699088
rect 234822 699066 234836 699068
rect 234892 699066 234916 699068
rect 234972 699066 234996 699068
rect 235052 699066 235076 699068
rect 235132 699066 235156 699068
rect 235212 699066 235236 699068
rect 235292 699066 235316 699068
rect 235372 699066 235386 699068
rect 235066 699014 235076 699066
rect 235132 699014 235142 699066
rect 234822 699012 234836 699014
rect 234892 699012 234916 699014
rect 234972 699012 234996 699014
rect 235052 699012 235076 699014
rect 235132 699012 235156 699014
rect 235212 699012 235236 699014
rect 235292 699012 235316 699014
rect 235372 699012 235386 699014
rect 234822 698992 235386 699012
rect 235906 698320 235962 698329
rect 235906 698255 235962 698264
rect 235920 698222 235948 698255
rect 235908 698216 235960 698222
rect 237380 698216 237432 698222
rect 235908 698158 235960 698164
rect 237378 698184 237380 698193
rect 237432 698184 237434 698193
rect 237378 698119 237434 698128
rect 232964 696924 233016 696930
rect 232964 696866 233016 696872
rect 233056 696924 233108 696930
rect 233056 696866 233108 696872
rect 232976 696833 233004 696866
rect 232962 696824 233018 696833
rect 232962 696759 233018 696768
rect 229006 696008 229062 696017
rect 213734 695943 213790 695952
rect 229006 695943 229062 695952
rect 230386 696008 230442 696017
rect 233068 695994 233096 696866
rect 234526 696824 234582 696833
rect 234526 696759 234528 696768
rect 234580 696759 234582 696768
rect 234528 696730 234580 696736
rect 234526 696416 234582 696425
rect 234526 696351 234528 696360
rect 234580 696351 234582 696360
rect 234528 696322 234580 696328
rect 232806 695966 233096 695994
rect 237484 695980 237512 701898
rect 242256 700596 242308 700602
rect 242256 700538 242308 700544
rect 237564 698216 237616 698222
rect 237562 698184 237564 698193
rect 237616 698184 237618 698193
rect 237562 698119 237618 698128
rect 242268 695980 242296 700538
rect 246948 700528 247000 700534
rect 246948 700470 247000 700476
rect 244094 699272 244150 699281
rect 244278 699272 244334 699281
rect 244150 699230 244228 699258
rect 244094 699207 244150 699216
rect 244094 699000 244150 699009
rect 244200 698970 244228 699230
rect 244278 699207 244334 699216
rect 244292 698970 244320 699207
rect 244370 699000 244426 699009
rect 244094 698935 244096 698944
rect 244148 698935 244150 698944
rect 244188 698964 244240 698970
rect 244096 698906 244148 698912
rect 244188 698906 244240 698912
rect 244280 698964 244332 698970
rect 244370 698935 244372 698944
rect 244280 698906 244332 698912
rect 244424 698935 244426 698944
rect 244372 698906 244424 698912
rect 244278 696824 244334 696833
rect 244278 696759 244280 696768
rect 244332 696759 244334 696768
rect 244280 696730 244332 696736
rect 244278 696416 244334 696425
rect 244278 696351 244280 696360
rect 244332 696351 244334 696360
rect 244280 696322 244332 696328
rect 246960 695980 246988 700470
rect 251088 699848 251140 699854
rect 251088 699790 251140 699796
rect 251100 699718 251128 699790
rect 251088 699712 251140 699718
rect 251088 699654 251140 699660
rect 248326 698320 248382 698329
rect 248326 698255 248382 698264
rect 248340 696930 248368 698255
rect 248328 696924 248380 696930
rect 248328 696866 248380 696872
rect 248420 696924 248472 696930
rect 248420 696866 248472 696872
rect 248432 696833 248460 696866
rect 248418 696824 248474 696833
rect 248418 696759 248474 696768
rect 251086 696008 251142 696017
rect 230386 695943 230442 695952
rect 251652 695980 251680 701966
rect 252822 701788 253386 701808
rect 252822 701786 252836 701788
rect 252892 701786 252916 701788
rect 252972 701786 252996 701788
rect 253052 701786 253076 701788
rect 253132 701786 253156 701788
rect 253212 701786 253236 701788
rect 253292 701786 253316 701788
rect 253372 701786 253386 701788
rect 253066 701734 253076 701786
rect 253132 701734 253142 701786
rect 252822 701732 252836 701734
rect 252892 701732 252916 701734
rect 252972 701732 252996 701734
rect 253052 701732 253076 701734
rect 253132 701732 253156 701734
rect 253212 701732 253236 701734
rect 253292 701732 253316 701734
rect 253372 701732 253386 701734
rect 252822 701712 253386 701732
rect 261116 701004 261168 701010
rect 261116 700946 261168 700952
rect 252822 700700 253386 700720
rect 252822 700698 252836 700700
rect 252892 700698 252916 700700
rect 252972 700698 252996 700700
rect 253052 700698 253076 700700
rect 253132 700698 253156 700700
rect 253212 700698 253236 700700
rect 253292 700698 253316 700700
rect 253372 700698 253386 700700
rect 253066 700646 253076 700698
rect 253132 700646 253142 700698
rect 252822 700644 252836 700646
rect 252892 700644 252916 700646
rect 252972 700644 252996 700646
rect 253052 700644 253076 700646
rect 253132 700644 253156 700646
rect 253212 700644 253236 700646
rect 253292 700644 253316 700646
rect 253372 700644 253386 700646
rect 252822 700624 253386 700644
rect 256424 700256 256476 700262
rect 256424 700198 256476 700204
rect 252822 699612 253386 699632
rect 252822 699610 252836 699612
rect 252892 699610 252916 699612
rect 252972 699610 252996 699612
rect 253052 699610 253076 699612
rect 253132 699610 253156 699612
rect 253212 699610 253236 699612
rect 253292 699610 253316 699612
rect 253372 699610 253386 699612
rect 253066 699558 253076 699610
rect 253132 699558 253142 699610
rect 252822 699556 252836 699558
rect 252892 699556 252916 699558
rect 252972 699556 252996 699558
rect 253052 699556 253076 699558
rect 253132 699556 253156 699558
rect 253212 699556 253236 699558
rect 253292 699556 253316 699558
rect 253372 699556 253386 699558
rect 252822 699536 253386 699556
rect 253754 699000 253810 699009
rect 253754 698935 253756 698944
rect 253808 698935 253810 698944
rect 253848 698964 253900 698970
rect 253756 698906 253808 698912
rect 253848 698906 253900 698912
rect 252822 698524 253386 698544
rect 252822 698522 252836 698524
rect 252892 698522 252916 698524
rect 252972 698522 252996 698524
rect 253052 698522 253076 698524
rect 253132 698522 253156 698524
rect 253212 698522 253236 698524
rect 253292 698522 253316 698524
rect 253372 698522 253386 698524
rect 253066 698470 253076 698522
rect 253132 698470 253142 698522
rect 252822 698468 252836 698470
rect 252892 698468 252916 698470
rect 252972 698468 252996 698470
rect 253052 698468 253076 698470
rect 253132 698468 253156 698470
rect 253212 698468 253236 698470
rect 253292 698468 253316 698470
rect 253372 698468 253386 698470
rect 252822 698448 253386 698468
rect 253860 698329 253888 698906
rect 253846 698320 253902 698329
rect 253846 698255 253902 698264
rect 253848 698216 253900 698222
rect 253846 698184 253848 698193
rect 254032 698216 254084 698222
rect 253900 698184 253902 698193
rect 253846 698119 253902 698128
rect 254030 698184 254032 698193
rect 254084 698184 254086 698193
rect 254030 698119 254086 698128
rect 253846 696416 253902 696425
rect 253846 696351 253848 696360
rect 253900 696351 253902 696360
rect 253848 696322 253900 696328
rect 256436 695980 256464 700198
rect 259460 699780 259512 699786
rect 259460 699722 259512 699728
rect 259472 699553 259500 699722
rect 259458 699544 259514 699553
rect 259458 699479 259514 699488
rect 261128 695980 261156 700946
rect 265900 699984 265952 699990
rect 265900 699926 265952 699932
rect 263598 696416 263654 696425
rect 263598 696351 263600 696360
rect 263652 696351 263654 696360
rect 263600 696322 263652 696328
rect 265622 696008 265678 696017
rect 251086 695943 251142 695952
rect 265912 695980 265940 699926
rect 267660 699854 267688 703520
rect 270822 701244 271386 701264
rect 270822 701242 270836 701244
rect 270892 701242 270916 701244
rect 270972 701242 270996 701244
rect 271052 701242 271076 701244
rect 271132 701242 271156 701244
rect 271212 701242 271236 701244
rect 271292 701242 271316 701244
rect 271372 701242 271386 701244
rect 271066 701190 271076 701242
rect 271132 701190 271142 701242
rect 270822 701188 270836 701190
rect 270892 701188 270916 701190
rect 270972 701188 270996 701190
rect 271052 701188 271076 701190
rect 271132 701188 271156 701190
rect 271212 701188 271236 701190
rect 271292 701188 271316 701190
rect 271372 701188 271386 701190
rect 270822 701168 271386 701188
rect 270822 700156 271386 700176
rect 270822 700154 270836 700156
rect 270892 700154 270916 700156
rect 270972 700154 270996 700156
rect 271052 700154 271076 700156
rect 271132 700154 271156 700156
rect 271212 700154 271236 700156
rect 271292 700154 271316 700156
rect 271372 700154 271386 700156
rect 271066 700102 271076 700154
rect 271132 700102 271142 700154
rect 270822 700100 270836 700102
rect 270892 700100 270916 700102
rect 270972 700100 270996 700102
rect 271052 700100 271076 700102
rect 271132 700100 271156 700102
rect 271212 700100 271236 700102
rect 271292 700100 271316 700102
rect 271372 700100 271386 700102
rect 270822 700080 271386 700100
rect 283102 700088 283158 700097
rect 283102 700023 283158 700032
rect 267648 699848 267700 699854
rect 267648 699790 267700 699796
rect 273260 699848 273312 699854
rect 273260 699790 273312 699796
rect 273902 699816 273958 699825
rect 270592 699780 270644 699786
rect 270592 699722 270644 699728
rect 267646 699272 267702 699281
rect 267646 699207 267648 699216
rect 267700 699207 267702 699216
rect 267648 699178 267700 699184
rect 270604 695980 270632 699722
rect 273272 699417 273300 699790
rect 273902 699751 273904 699760
rect 273956 699751 273958 699760
rect 273904 699722 273956 699728
rect 282920 699712 282972 699718
rect 280066 699680 280122 699689
rect 283012 699712 283064 699718
rect 282920 699654 282972 699660
rect 283010 699680 283012 699689
rect 283064 699680 283066 699689
rect 280066 699615 280122 699624
rect 273258 699408 273314 699417
rect 273258 699343 273314 699352
rect 273352 699372 273404 699378
rect 273352 699314 273404 699320
rect 273364 699281 273392 699314
rect 273350 699272 273406 699281
rect 273350 699207 273406 699216
rect 277398 699272 277454 699281
rect 277398 699207 277454 699216
rect 270822 699068 271386 699088
rect 270822 699066 270836 699068
rect 270892 699066 270916 699068
rect 270972 699066 270996 699068
rect 271052 699066 271076 699068
rect 271132 699066 271156 699068
rect 271212 699066 271236 699068
rect 271292 699066 271316 699068
rect 271372 699066 271386 699068
rect 271066 699014 271076 699066
rect 271132 699014 271142 699066
rect 270822 699012 270836 699014
rect 270892 699012 270916 699014
rect 270972 699012 270996 699014
rect 271052 699012 271076 699014
rect 271132 699012 271156 699014
rect 271212 699012 271236 699014
rect 271292 699012 271316 699014
rect 271372 699012 271386 699014
rect 270822 698992 271386 699012
rect 277412 698193 277440 699207
rect 275742 698184 275798 698193
rect 275742 698119 275798 698128
rect 277398 698184 277454 698193
rect 277398 698119 277454 698128
rect 273166 696416 273222 696425
rect 273166 696351 273168 696360
rect 273220 696351 273222 696360
rect 273168 696322 273220 696328
rect 275756 695994 275784 698119
rect 275402 695966 275784 695994
rect 280080 695980 280108 699615
rect 282932 699145 282960 699654
rect 283010 699615 283066 699624
rect 283010 699408 283066 699417
rect 283010 699343 283012 699352
rect 283064 699343 283066 699352
rect 283012 699314 283064 699320
rect 282918 699136 282974 699145
rect 282918 699071 282974 699080
rect 283116 698986 283144 700023
rect 283746 699816 283802 699825
rect 283852 699786 283880 703520
rect 288822 701788 289386 701808
rect 288822 701786 288836 701788
rect 288892 701786 288916 701788
rect 288972 701786 288996 701788
rect 289052 701786 289076 701788
rect 289132 701786 289156 701788
rect 289212 701786 289236 701788
rect 289292 701786 289316 701788
rect 289372 701786 289386 701788
rect 289066 701734 289076 701786
rect 289132 701734 289142 701786
rect 288822 701732 288836 701734
rect 288892 701732 288916 701734
rect 288972 701732 288996 701734
rect 289052 701732 289076 701734
rect 289132 701732 289156 701734
rect 289212 701732 289236 701734
rect 289292 701732 289316 701734
rect 289372 701732 289386 701734
rect 288822 701712 289386 701732
rect 288822 700700 289386 700720
rect 288822 700698 288836 700700
rect 288892 700698 288916 700700
rect 288972 700698 288996 700700
rect 289052 700698 289076 700700
rect 289132 700698 289156 700700
rect 289212 700698 289236 700700
rect 289292 700698 289316 700700
rect 289372 700698 289386 700700
rect 289066 700646 289076 700698
rect 289132 700646 289142 700698
rect 288822 700644 288836 700646
rect 288892 700644 288916 700646
rect 288972 700644 288996 700646
rect 289052 700644 289076 700646
rect 289132 700644 289156 700646
rect 289212 700644 289236 700646
rect 289292 700644 289316 700646
rect 289372 700644 289386 700646
rect 288822 700624 289386 700644
rect 296536 700392 296588 700398
rect 296536 700334 296588 700340
rect 296628 700392 296680 700398
rect 296628 700334 296680 700340
rect 296548 700233 296576 700334
rect 296534 700224 296590 700233
rect 296534 700159 296590 700168
rect 296640 700097 296668 700334
rect 298650 700224 298706 700233
rect 298650 700159 298706 700168
rect 296626 700088 296682 700097
rect 296626 700023 296682 700032
rect 298006 699952 298062 699961
rect 296720 699916 296772 699922
rect 298006 699887 298008 699896
rect 296720 699858 296772 699864
rect 298060 699887 298062 699896
rect 298008 699858 298060 699864
rect 296732 699825 296760 699858
rect 288714 699816 288770 699825
rect 283746 699751 283748 699760
rect 283800 699751 283802 699760
rect 283840 699780 283892 699786
rect 283748 699722 283800 699728
rect 283840 699722 283892 699728
rect 288532 699780 288584 699786
rect 288714 699751 288770 699760
rect 296718 699816 296774 699825
rect 296718 699751 296774 699760
rect 296904 699780 296956 699786
rect 288532 699722 288584 699728
rect 282932 698970 283144 698986
rect 282920 698964 283144 698970
rect 282972 698958 283144 698964
rect 282920 698906 282972 698912
rect 284484 696924 284536 696930
rect 284484 696866 284536 696872
rect 282918 696416 282974 696425
rect 282918 696351 282920 696360
rect 282972 696351 282974 696360
rect 282920 696322 282972 696328
rect 284496 695994 284524 696866
rect 288544 696538 288572 699722
rect 288728 699718 288756 699751
rect 296904 699722 296956 699728
rect 288716 699712 288768 699718
rect 288716 699654 288768 699660
rect 292396 699712 292448 699718
rect 292396 699654 292448 699660
rect 292488 699712 292540 699718
rect 292488 699654 292540 699660
rect 288822 699612 289386 699632
rect 288822 699610 288836 699612
rect 288892 699610 288916 699612
rect 288972 699610 288996 699612
rect 289052 699610 289076 699612
rect 289132 699610 289156 699612
rect 289212 699610 289236 699612
rect 289292 699610 289316 699612
rect 289372 699610 289386 699612
rect 289066 699558 289076 699610
rect 289132 699558 289142 699610
rect 288822 699556 288836 699558
rect 288892 699556 288916 699558
rect 288972 699556 288996 699558
rect 289052 699556 289076 699558
rect 289132 699556 289156 699558
rect 289212 699556 289236 699558
rect 289292 699556 289316 699558
rect 289372 699556 289386 699558
rect 288822 699536 289386 699556
rect 289726 699544 289782 699553
rect 289726 699479 289782 699488
rect 288822 698524 289386 698544
rect 288822 698522 288836 698524
rect 288892 698522 288916 698524
rect 288972 698522 288996 698524
rect 289052 698522 289076 698524
rect 289132 698522 289156 698524
rect 289212 698522 289236 698524
rect 289292 698522 289316 698524
rect 289372 698522 289386 698524
rect 289066 698470 289076 698522
rect 289132 698470 289142 698522
rect 288822 698468 288836 698470
rect 288892 698468 288916 698470
rect 288972 698468 288996 698470
rect 289052 698468 289076 698470
rect 289132 698468 289156 698470
rect 289212 698468 289236 698470
rect 289292 698468 289316 698470
rect 289372 698468 289386 698470
rect 288822 698448 289386 698468
rect 289740 696862 289768 699479
rect 292408 699417 292436 699654
rect 292394 699408 292450 699417
rect 292394 699343 292450 699352
rect 292500 699281 292528 699654
rect 296916 699553 296944 699722
rect 296902 699544 296958 699553
rect 296902 699479 296958 699488
rect 294050 699408 294106 699417
rect 294050 699343 294106 699352
rect 296536 699372 296588 699378
rect 292486 699272 292542 699281
rect 292486 699207 292542 699216
rect 289728 696856 289780 696862
rect 289728 696798 289780 696804
rect 288544 696510 289124 696538
rect 284496 695966 284878 695994
rect 265622 695943 265678 695952
rect 119986 695736 120042 695745
rect 119986 695671 120042 695680
rect 53288 695632 53340 695638
rect 52946 695580 53288 695586
rect 52946 695574 53340 695580
rect 120000 695586 120028 695671
rect 205560 695609 205588 695943
rect 213748 695609 213776 695943
rect 120170 695600 120226 695609
rect 52946 695558 53328 695574
rect 120000 695558 120170 695586
rect 176198 695600 176254 695609
rect 175950 695558 176198 695586
rect 120170 695535 120226 695544
rect 176198 695535 176254 695544
rect 205546 695600 205602 695609
rect 205546 695535 205602 695544
rect 213734 695600 213790 695609
rect 213734 695535 213790 695544
rect 215206 695600 215262 695609
rect 215262 695558 215340 695586
rect 215206 695535 215262 695544
rect 215312 695473 215340 695558
rect 229020 695473 229048 695943
rect 230400 695609 230428 695943
rect 234618 695736 234674 695745
rect 234618 695671 234674 695680
rect 230386 695600 230442 695609
rect 230386 695535 230442 695544
rect 234526 695600 234582 695609
rect 234632 695586 234660 695671
rect 251100 695609 251128 695943
rect 265636 695745 265664 695943
rect 289096 695858 289124 696510
rect 292486 696416 292542 696425
rect 292486 696351 292488 696360
rect 292540 696351 292542 696360
rect 292488 696322 292540 696328
rect 294064 695994 294092 699343
rect 296536 699314 296588 699320
rect 296628 699372 296680 699378
rect 296628 699314 296680 699320
rect 296548 699281 296576 699314
rect 296534 699272 296590 699281
rect 296534 699207 296590 699216
rect 296640 699145 296668 699314
rect 296626 699136 296682 699145
rect 296626 699071 296682 699080
rect 298664 695994 298692 700159
rect 300136 699961 300164 703520
rect 324822 701788 325386 701808
rect 324822 701786 324836 701788
rect 324892 701786 324916 701788
rect 324972 701786 324996 701788
rect 325052 701786 325076 701788
rect 325132 701786 325156 701788
rect 325212 701786 325236 701788
rect 325292 701786 325316 701788
rect 325372 701786 325386 701788
rect 325066 701734 325076 701786
rect 325132 701734 325142 701786
rect 324822 701732 324836 701734
rect 324892 701732 324916 701734
rect 324972 701732 324996 701734
rect 325052 701732 325076 701734
rect 325132 701732 325156 701734
rect 325212 701732 325236 701734
rect 325292 701732 325316 701734
rect 325372 701732 325386 701734
rect 324822 701712 325386 701732
rect 306822 701244 307386 701264
rect 306822 701242 306836 701244
rect 306892 701242 306916 701244
rect 306972 701242 306996 701244
rect 307052 701242 307076 701244
rect 307132 701242 307156 701244
rect 307212 701242 307236 701244
rect 307292 701242 307316 701244
rect 307372 701242 307386 701244
rect 307066 701190 307076 701242
rect 307132 701190 307142 701242
rect 306822 701188 306836 701190
rect 306892 701188 306916 701190
rect 306972 701188 306996 701190
rect 307052 701188 307076 701190
rect 307132 701188 307156 701190
rect 307212 701188 307236 701190
rect 307292 701188 307316 701190
rect 307372 701188 307386 701190
rect 306822 701168 307386 701188
rect 317972 700936 318024 700942
rect 317972 700878 318024 700884
rect 313188 700868 313240 700874
rect 313188 700810 313240 700816
rect 306822 700156 307386 700176
rect 306822 700154 306836 700156
rect 306892 700154 306916 700156
rect 306972 700154 306996 700156
rect 307052 700154 307076 700156
rect 307132 700154 307156 700156
rect 307212 700154 307236 700156
rect 307292 700154 307316 700156
rect 307372 700154 307386 700156
rect 307066 700102 307076 700154
rect 307132 700102 307142 700154
rect 306822 700100 306836 700102
rect 306892 700100 306916 700102
rect 306972 700100 306996 700102
rect 307052 700100 307076 700102
rect 307132 700100 307156 700102
rect 307212 700100 307236 700102
rect 307292 700100 307316 700102
rect 307372 700100 307386 700102
rect 306822 700080 307386 700100
rect 308496 700052 308548 700058
rect 308496 699994 308548 700000
rect 308588 700052 308640 700058
rect 308588 699994 308640 700000
rect 300122 699952 300178 699961
rect 300122 699887 300178 699896
rect 302330 699952 302386 699961
rect 302330 699887 302386 699896
rect 302344 699718 302372 699887
rect 303618 699816 303674 699825
rect 303618 699751 303674 699760
rect 302332 699712 302384 699718
rect 302332 699654 302384 699660
rect 302330 699272 302386 699281
rect 302330 699207 302332 699216
rect 302384 699207 302386 699216
rect 302332 699178 302384 699184
rect 299480 696788 299532 696794
rect 299480 696730 299532 696736
rect 299492 696697 299520 696730
rect 299478 696688 299534 696697
rect 299478 696623 299534 696632
rect 303632 695994 303660 699751
rect 306822 699068 307386 699088
rect 306822 699066 306836 699068
rect 306892 699066 306916 699068
rect 306972 699066 306996 699068
rect 307052 699066 307076 699068
rect 307132 699066 307156 699068
rect 307212 699066 307236 699068
rect 307292 699066 307316 699068
rect 307372 699066 307386 699068
rect 307066 699014 307076 699066
rect 307132 699014 307142 699066
rect 306822 699012 306836 699014
rect 306892 699012 306916 699014
rect 306972 699012 306996 699014
rect 307052 699012 307076 699014
rect 307132 699012 307156 699014
rect 307212 699012 307236 699014
rect 307292 699012 307316 699014
rect 307372 699012 307386 699014
rect 306822 698992 307386 699012
rect 294064 695966 294354 695994
rect 298664 695966 299046 695994
rect 303632 695966 303738 695994
rect 308508 695980 308536 699994
rect 308600 699961 308628 699994
rect 308586 699952 308642 699961
rect 308586 699887 308642 699896
rect 311992 699712 312044 699718
rect 311992 699654 312044 699660
rect 312004 699281 312032 699654
rect 311990 699272 312046 699281
rect 311716 699236 311768 699242
rect 311990 699207 312046 699216
rect 311716 699178 311768 699184
rect 311728 698986 311756 699178
rect 311990 699000 312046 699009
rect 311728 698958 311990 698986
rect 311990 698935 312046 698944
rect 309140 696856 309192 696862
rect 309138 696824 309140 696833
rect 309192 696824 309194 696833
rect 309048 696788 309100 696794
rect 309138 696759 309194 696768
rect 309048 696730 309100 696736
rect 309060 696697 309088 696730
rect 309046 696688 309102 696697
rect 309046 696623 309102 696632
rect 313200 695980 313228 700810
rect 317984 695980 318012 700878
rect 322664 700800 322716 700806
rect 322664 700742 322716 700748
rect 321650 699272 321706 699281
rect 321650 699207 321706 699216
rect 321664 699174 321692 699207
rect 321652 699168 321704 699174
rect 321558 699136 321614 699145
rect 321652 699110 321704 699116
rect 321558 699071 321614 699080
rect 321572 698970 321600 699071
rect 321650 699000 321706 699009
rect 321560 698964 321612 698970
rect 321650 698935 321652 698944
rect 321560 698906 321612 698912
rect 321704 698935 321706 698944
rect 321652 698906 321704 698912
rect 318614 696824 318670 696833
rect 318614 696759 318670 696768
rect 321560 696788 321612 696794
rect 318628 696674 318656 696759
rect 321560 696730 321612 696736
rect 321572 696697 321600 696730
rect 318798 696688 318854 696697
rect 318628 696646 318798 696674
rect 318798 696623 318854 696632
rect 321558 696688 321614 696697
rect 321558 696623 321614 696632
rect 322676 695980 322704 700742
rect 324822 700700 325386 700720
rect 324822 700698 324836 700700
rect 324892 700698 324916 700700
rect 324972 700698 324996 700700
rect 325052 700698 325076 700700
rect 325132 700698 325156 700700
rect 325212 700698 325236 700700
rect 325292 700698 325316 700700
rect 325372 700698 325386 700700
rect 325066 700646 325076 700698
rect 325132 700646 325142 700698
rect 324822 700644 324836 700646
rect 324892 700644 324916 700646
rect 324972 700644 324996 700646
rect 325052 700644 325076 700646
rect 325132 700644 325156 700646
rect 325212 700644 325236 700646
rect 325292 700644 325316 700646
rect 325372 700644 325386 700646
rect 324822 700624 325386 700644
rect 332140 700460 332192 700466
rect 332140 700402 332192 700408
rect 327448 700324 327500 700330
rect 327448 700266 327500 700272
rect 324822 699612 325386 699632
rect 324822 699610 324836 699612
rect 324892 699610 324916 699612
rect 324972 699610 324996 699612
rect 325052 699610 325076 699612
rect 325132 699610 325156 699612
rect 325212 699610 325236 699612
rect 325292 699610 325316 699612
rect 325372 699610 325386 699612
rect 325066 699558 325076 699610
rect 325132 699558 325142 699610
rect 324822 699556 324836 699558
rect 324892 699556 324916 699558
rect 324972 699556 324996 699558
rect 325052 699556 325076 699558
rect 325132 699556 325156 699558
rect 325212 699556 325236 699558
rect 325292 699556 325316 699558
rect 325372 699556 325386 699558
rect 324822 699536 325386 699556
rect 324822 698524 325386 698544
rect 324822 698522 324836 698524
rect 324892 698522 324916 698524
rect 324972 698522 324996 698524
rect 325052 698522 325076 698524
rect 325132 698522 325156 698524
rect 325212 698522 325236 698524
rect 325292 698522 325316 698524
rect 325372 698522 325386 698524
rect 325066 698470 325076 698522
rect 325132 698470 325142 698522
rect 324822 698468 324836 698470
rect 324892 698468 324916 698470
rect 324972 698468 324996 698470
rect 325052 698468 325076 698470
rect 325132 698468 325156 698470
rect 325212 698468 325236 698470
rect 325292 698468 325316 698470
rect 325372 698468 325386 698470
rect 324822 698448 325386 698468
rect 327460 695980 327488 700266
rect 331312 699916 331364 699922
rect 331312 699858 331364 699864
rect 331324 699281 331352 699858
rect 331034 699272 331090 699281
rect 331034 699207 331090 699216
rect 331310 699272 331366 699281
rect 331310 699207 331366 699216
rect 331048 699174 331076 699207
rect 331036 699168 331088 699174
rect 331128 699168 331180 699174
rect 331036 699110 331088 699116
rect 331126 699136 331128 699145
rect 331180 699136 331182 699145
rect 331126 699071 331182 699080
rect 328460 696788 328512 696794
rect 328460 696730 328512 696736
rect 328472 696697 328500 696730
rect 328458 696688 328514 696697
rect 328458 696623 328514 696632
rect 328366 696008 328422 696017
rect 332152 695980 332180 700402
rect 332520 699854 332548 703520
rect 342822 701244 343386 701264
rect 342822 701242 342836 701244
rect 342892 701242 342916 701244
rect 342972 701242 342996 701244
rect 343052 701242 343076 701244
rect 343132 701242 343156 701244
rect 343212 701242 343236 701244
rect 343292 701242 343316 701244
rect 343372 701242 343386 701244
rect 343066 701190 343076 701242
rect 343132 701190 343142 701242
rect 342822 701188 342836 701190
rect 342892 701188 342916 701190
rect 342972 701188 342996 701190
rect 343052 701188 343076 701190
rect 343132 701188 343156 701190
rect 343212 701188 343236 701190
rect 343292 701188 343316 701190
rect 343372 701188 343386 701190
rect 342822 701168 343386 701188
rect 336922 701040 336978 701049
rect 336922 700975 336978 700984
rect 332508 699848 332560 699854
rect 332508 699790 332560 699796
rect 336936 695980 336964 700975
rect 346306 700496 346362 700505
rect 346306 700431 346362 700440
rect 341614 700360 341670 700369
rect 341614 700295 341670 700304
rect 340694 699272 340750 699281
rect 340694 699207 340750 699216
rect 340708 699174 340736 699207
rect 340696 699168 340748 699174
rect 340696 699110 340748 699116
rect 338118 696824 338174 696833
rect 338118 696759 338174 696768
rect 338026 696688 338082 696697
rect 338132 696674 338160 696759
rect 338082 696646 338160 696674
rect 338026 696623 338082 696632
rect 341628 695980 341656 700295
rect 342822 700156 343386 700176
rect 342822 700154 342836 700156
rect 342892 700154 342916 700156
rect 342972 700154 342996 700156
rect 343052 700154 343076 700156
rect 343132 700154 343156 700156
rect 343212 700154 343236 700156
rect 343292 700154 343316 700156
rect 343372 700154 343386 700156
rect 343066 700102 343076 700154
rect 343132 700102 343142 700154
rect 342822 700100 342836 700102
rect 342892 700100 342916 700102
rect 342972 700100 342996 700102
rect 343052 700100 343076 700102
rect 343132 700100 343156 700102
rect 343212 700100 343236 700102
rect 343292 700100 343316 700102
rect 343372 700100 343386 700102
rect 342822 700080 343386 700100
rect 344926 699272 344982 699281
rect 344926 699207 344982 699216
rect 342822 699068 343386 699088
rect 342822 699066 342836 699068
rect 342892 699066 342916 699068
rect 342972 699066 342996 699068
rect 343052 699066 343076 699068
rect 343132 699066 343156 699068
rect 343212 699066 343236 699068
rect 343292 699066 343316 699068
rect 343372 699066 343386 699068
rect 343066 699014 343076 699066
rect 343132 699014 343142 699066
rect 342822 699012 342836 699014
rect 342892 699012 342916 699014
rect 342972 699012 342996 699014
rect 343052 699012 343076 699014
rect 343132 699012 343156 699014
rect 343212 699012 343236 699014
rect 343292 699012 343316 699014
rect 343372 699012 343386 699014
rect 342822 698992 343386 699012
rect 344940 698970 344968 699207
rect 344928 698964 344980 698970
rect 344928 698906 344980 698912
rect 342626 696824 342682 696833
rect 342626 696759 342628 696768
rect 342680 696759 342682 696768
rect 342628 696730 342680 696736
rect 346320 695980 346348 700431
rect 348804 699922 348832 703520
rect 360822 701788 361386 701808
rect 360822 701786 360836 701788
rect 360892 701786 360916 701788
rect 360972 701786 360996 701788
rect 361052 701786 361076 701788
rect 361132 701786 361156 701788
rect 361212 701786 361236 701788
rect 361292 701786 361316 701788
rect 361372 701786 361386 701788
rect 361066 701734 361076 701786
rect 361132 701734 361142 701786
rect 360822 701732 360836 701734
rect 360892 701732 360916 701734
rect 360972 701732 360996 701734
rect 361052 701732 361076 701734
rect 361132 701732 361156 701734
rect 361212 701732 361236 701734
rect 361292 701732 361316 701734
rect 361372 701732 361386 701734
rect 360822 701712 361386 701732
rect 360822 700700 361386 700720
rect 360822 700698 360836 700700
rect 360892 700698 360916 700700
rect 360972 700698 360996 700700
rect 361052 700698 361076 700700
rect 361132 700698 361156 700700
rect 361212 700698 361236 700700
rect 361292 700698 361316 700700
rect 361372 700698 361386 700700
rect 361066 700646 361076 700698
rect 361132 700646 361142 700698
rect 360822 700644 360836 700646
rect 360892 700644 360916 700646
rect 360972 700644 360996 700646
rect 361052 700644 361076 700646
rect 361132 700644 361156 700646
rect 361212 700644 361236 700646
rect 361292 700644 361316 700646
rect 361372 700644 361386 700646
rect 360822 700624 361386 700644
rect 364996 699990 365024 703520
rect 396822 701788 397386 701808
rect 396822 701786 396836 701788
rect 396892 701786 396916 701788
rect 396972 701786 396996 701788
rect 397052 701786 397076 701788
rect 397132 701786 397156 701788
rect 397212 701786 397236 701788
rect 397292 701786 397316 701788
rect 397372 701786 397386 701788
rect 397066 701734 397076 701786
rect 397132 701734 397142 701786
rect 396822 701732 396836 701734
rect 396892 701732 396916 701734
rect 396972 701732 396996 701734
rect 397052 701732 397076 701734
rect 397132 701732 397156 701734
rect 397212 701732 397236 701734
rect 397292 701732 397316 701734
rect 397372 701732 397386 701734
rect 396822 701712 397386 701732
rect 378822 701244 379386 701264
rect 378822 701242 378836 701244
rect 378892 701242 378916 701244
rect 378972 701242 378996 701244
rect 379052 701242 379076 701244
rect 379132 701242 379156 701244
rect 379212 701242 379236 701244
rect 379292 701242 379316 701244
rect 379372 701242 379386 701244
rect 379066 701190 379076 701242
rect 379132 701190 379142 701242
rect 378822 701188 378836 701190
rect 378892 701188 378916 701190
rect 378972 701188 378996 701190
rect 379052 701188 379076 701190
rect 379132 701188 379156 701190
rect 379212 701188 379236 701190
rect 379292 701188 379316 701190
rect 379372 701188 379386 701190
rect 378822 701168 379386 701188
rect 396822 700700 397386 700720
rect 396822 700698 396836 700700
rect 396892 700698 396916 700700
rect 396972 700698 396996 700700
rect 397052 700698 397076 700700
rect 397132 700698 397156 700700
rect 397212 700698 397236 700700
rect 397292 700698 397316 700700
rect 397372 700698 397386 700700
rect 397066 700646 397076 700698
rect 397132 700646 397142 700698
rect 396822 700644 396836 700646
rect 396892 700644 396916 700646
rect 396972 700644 396996 700646
rect 397052 700644 397076 700646
rect 397132 700644 397156 700646
rect 397212 700644 397236 700646
rect 397292 700644 397316 700646
rect 397372 700644 397386 700646
rect 396822 700624 397386 700644
rect 397472 700262 397500 703520
rect 413664 701010 413692 703520
rect 429856 702030 429884 703520
rect 429844 702024 429896 702030
rect 429844 701966 429896 701972
rect 432822 701788 433386 701808
rect 432822 701786 432836 701788
rect 432892 701786 432916 701788
rect 432972 701786 432996 701788
rect 433052 701786 433076 701788
rect 433132 701786 433156 701788
rect 433212 701786 433236 701788
rect 433292 701786 433316 701788
rect 433372 701786 433386 701788
rect 433066 701734 433076 701786
rect 433132 701734 433142 701786
rect 432822 701732 432836 701734
rect 432892 701732 432916 701734
rect 432972 701732 432996 701734
rect 433052 701732 433076 701734
rect 433132 701732 433156 701734
rect 433212 701732 433236 701734
rect 433292 701732 433316 701734
rect 433372 701732 433386 701734
rect 432822 701712 433386 701732
rect 414822 701244 415386 701264
rect 414822 701242 414836 701244
rect 414892 701242 414916 701244
rect 414972 701242 414996 701244
rect 415052 701242 415076 701244
rect 415132 701242 415156 701244
rect 415212 701242 415236 701244
rect 415292 701242 415316 701244
rect 415372 701242 415386 701244
rect 415066 701190 415076 701242
rect 415132 701190 415142 701242
rect 414822 701188 414836 701190
rect 414892 701188 414916 701190
rect 414972 701188 414996 701190
rect 415052 701188 415076 701190
rect 415132 701188 415156 701190
rect 415212 701188 415236 701190
rect 415292 701188 415316 701190
rect 415372 701188 415386 701190
rect 414822 701168 415386 701188
rect 450822 701244 451386 701264
rect 450822 701242 450836 701244
rect 450892 701242 450916 701244
rect 450972 701242 450996 701244
rect 451052 701242 451076 701244
rect 451132 701242 451156 701244
rect 451212 701242 451236 701244
rect 451292 701242 451316 701244
rect 451372 701242 451386 701244
rect 451066 701190 451076 701242
rect 451132 701190 451142 701242
rect 450822 701188 450836 701190
rect 450892 701188 450916 701190
rect 450972 701188 450996 701190
rect 451052 701188 451076 701190
rect 451132 701188 451156 701190
rect 451212 701188 451236 701190
rect 451292 701188 451316 701190
rect 451372 701188 451386 701190
rect 450822 701168 451386 701188
rect 413652 701004 413704 701010
rect 413652 700946 413704 700952
rect 432822 700700 433386 700720
rect 432822 700698 432836 700700
rect 432892 700698 432916 700700
rect 432972 700698 432996 700700
rect 433052 700698 433076 700700
rect 433132 700698 433156 700700
rect 433212 700698 433236 700700
rect 433292 700698 433316 700700
rect 433372 700698 433386 700700
rect 433066 700646 433076 700698
rect 433132 700646 433142 700698
rect 432822 700644 432836 700646
rect 432892 700644 432916 700646
rect 432972 700644 432996 700646
rect 433052 700644 433076 700646
rect 433132 700644 433156 700646
rect 433212 700644 433236 700646
rect 433292 700644 433316 700646
rect 433372 700644 433386 700646
rect 432822 700624 433386 700644
rect 462332 700602 462360 703520
rect 468822 701788 469386 701808
rect 468822 701786 468836 701788
rect 468892 701786 468916 701788
rect 468972 701786 468996 701788
rect 469052 701786 469076 701788
rect 469132 701786 469156 701788
rect 469212 701786 469236 701788
rect 469292 701786 469316 701788
rect 469372 701786 469386 701788
rect 469066 701734 469076 701786
rect 469132 701734 469142 701786
rect 468822 701732 468836 701734
rect 468892 701732 468916 701734
rect 468972 701732 468996 701734
rect 469052 701732 469076 701734
rect 469132 701732 469156 701734
rect 469212 701732 469236 701734
rect 469292 701732 469316 701734
rect 469372 701732 469386 701734
rect 468822 701712 469386 701732
rect 468822 700700 469386 700720
rect 468822 700698 468836 700700
rect 468892 700698 468916 700700
rect 468972 700698 468996 700700
rect 469052 700698 469076 700700
rect 469132 700698 469156 700700
rect 469212 700698 469236 700700
rect 469292 700698 469316 700700
rect 469372 700698 469386 700700
rect 469066 700646 469076 700698
rect 469132 700646 469142 700698
rect 468822 700644 468836 700646
rect 468892 700644 468916 700646
rect 468972 700644 468996 700646
rect 469052 700644 469076 700646
rect 469132 700644 469156 700646
rect 469212 700644 469236 700646
rect 469292 700644 469316 700646
rect 469372 700644 469386 700646
rect 468822 700624 469386 700644
rect 462320 700596 462372 700602
rect 462320 700538 462372 700544
rect 478524 700534 478552 703520
rect 494808 701962 494836 703520
rect 494796 701956 494848 701962
rect 494796 701898 494848 701904
rect 504822 701788 505386 701808
rect 504822 701786 504836 701788
rect 504892 701786 504916 701788
rect 504972 701786 504996 701788
rect 505052 701786 505076 701788
rect 505132 701786 505156 701788
rect 505212 701786 505236 701788
rect 505292 701786 505316 701788
rect 505372 701786 505386 701788
rect 505066 701734 505076 701786
rect 505132 701734 505142 701786
rect 504822 701732 504836 701734
rect 504892 701732 504916 701734
rect 504972 701732 504996 701734
rect 505052 701732 505076 701734
rect 505132 701732 505156 701734
rect 505212 701732 505236 701734
rect 505292 701732 505316 701734
rect 505372 701732 505386 701734
rect 504822 701712 505386 701732
rect 486822 701244 487386 701264
rect 486822 701242 486836 701244
rect 486892 701242 486916 701244
rect 486972 701242 486996 701244
rect 487052 701242 487076 701244
rect 487132 701242 487156 701244
rect 487212 701242 487236 701244
rect 487292 701242 487316 701244
rect 487372 701242 487386 701244
rect 487066 701190 487076 701242
rect 487132 701190 487142 701242
rect 486822 701188 486836 701190
rect 486892 701188 486916 701190
rect 486972 701188 486996 701190
rect 487052 701188 487076 701190
rect 487132 701188 487156 701190
rect 487212 701188 487236 701190
rect 487292 701188 487316 701190
rect 487372 701188 487386 701190
rect 486822 701168 487386 701188
rect 522822 701244 523386 701264
rect 522822 701242 522836 701244
rect 522892 701242 522916 701244
rect 522972 701242 522996 701244
rect 523052 701242 523076 701244
rect 523132 701242 523156 701244
rect 523212 701242 523236 701244
rect 523292 701242 523316 701244
rect 523372 701242 523386 701244
rect 523066 701190 523076 701242
rect 523132 701190 523142 701242
rect 522822 701188 522836 701190
rect 522892 701188 522916 701190
rect 522972 701188 522996 701190
rect 523052 701188 523076 701190
rect 523132 701188 523156 701190
rect 523212 701188 523236 701190
rect 523292 701188 523316 701190
rect 523372 701188 523386 701190
rect 522822 701168 523386 701188
rect 527192 700913 527220 703520
rect 540822 701788 541386 701808
rect 540822 701786 540836 701788
rect 540892 701786 540916 701788
rect 540972 701786 540996 701788
rect 541052 701786 541076 701788
rect 541132 701786 541156 701788
rect 541212 701786 541236 701788
rect 541292 701786 541316 701788
rect 541372 701786 541386 701788
rect 541066 701734 541076 701786
rect 541132 701734 541142 701786
rect 540822 701732 540836 701734
rect 540892 701732 540916 701734
rect 540972 701732 540996 701734
rect 541052 701732 541076 701734
rect 541132 701732 541156 701734
rect 541212 701732 541236 701734
rect 541292 701732 541316 701734
rect 541372 701732 541386 701734
rect 540822 701712 541386 701732
rect 527178 700904 527234 700913
rect 527178 700839 527234 700848
rect 504822 700700 505386 700720
rect 504822 700698 504836 700700
rect 504892 700698 504916 700700
rect 504972 700698 504996 700700
rect 505052 700698 505076 700700
rect 505132 700698 505156 700700
rect 505212 700698 505236 700700
rect 505292 700698 505316 700700
rect 505372 700698 505386 700700
rect 505066 700646 505076 700698
rect 505132 700646 505142 700698
rect 504822 700644 504836 700646
rect 504892 700644 504916 700646
rect 504972 700644 504996 700646
rect 505052 700644 505076 700646
rect 505132 700644 505156 700646
rect 505212 700644 505236 700646
rect 505292 700644 505316 700646
rect 505372 700644 505386 700646
rect 504822 700624 505386 700644
rect 540822 700700 541386 700720
rect 540822 700698 540836 700700
rect 540892 700698 540916 700700
rect 540972 700698 540996 700700
rect 541052 700698 541076 700700
rect 541132 700698 541156 700700
rect 541212 700698 541236 700700
rect 541292 700698 541316 700700
rect 541372 700698 541386 700700
rect 541066 700646 541076 700698
rect 541132 700646 541142 700698
rect 540822 700644 540836 700646
rect 540892 700644 540916 700646
rect 540972 700644 540996 700646
rect 541052 700644 541076 700646
rect 541132 700644 541156 700646
rect 541212 700644 541236 700646
rect 541292 700644 541316 700646
rect 541372 700644 541386 700646
rect 540822 700624 541386 700644
rect 478512 700528 478564 700534
rect 478512 700470 478564 700476
rect 543476 700398 543504 703520
rect 559668 701894 559696 703520
rect 559656 701888 559708 701894
rect 559656 701830 559708 701836
rect 576822 701788 577386 701808
rect 576822 701786 576836 701788
rect 576892 701786 576916 701788
rect 576972 701786 576996 701788
rect 577052 701786 577076 701788
rect 577132 701786 577156 701788
rect 577212 701786 577236 701788
rect 577292 701786 577316 701788
rect 577372 701786 577386 701788
rect 577066 701734 577076 701786
rect 577132 701734 577142 701786
rect 576822 701732 576836 701734
rect 576892 701732 576916 701734
rect 576972 701732 576996 701734
rect 577052 701732 577076 701734
rect 577132 701732 577156 701734
rect 577212 701732 577236 701734
rect 577292 701732 577316 701734
rect 577372 701732 577386 701734
rect 576822 701712 577386 701732
rect 558822 701244 559386 701264
rect 558822 701242 558836 701244
rect 558892 701242 558916 701244
rect 558972 701242 558996 701244
rect 559052 701242 559076 701244
rect 559132 701242 559156 701244
rect 559212 701242 559236 701244
rect 559292 701242 559316 701244
rect 559372 701242 559386 701244
rect 559066 701190 559076 701242
rect 559132 701190 559142 701242
rect 558822 701188 558836 701190
rect 558892 701188 558916 701190
rect 558972 701188 558996 701190
rect 559052 701188 559076 701190
rect 559132 701188 559156 701190
rect 559212 701188 559236 701190
rect 559292 701188 559316 701190
rect 559372 701188 559386 701190
rect 558822 701168 559386 701188
rect 576822 700700 577386 700720
rect 576822 700698 576836 700700
rect 576892 700698 576916 700700
rect 576972 700698 576996 700700
rect 577052 700698 577076 700700
rect 577132 700698 577156 700700
rect 577212 700698 577236 700700
rect 577292 700698 577316 700700
rect 577372 700698 577386 700700
rect 577066 700646 577076 700698
rect 577132 700646 577142 700698
rect 576822 700644 576836 700646
rect 576892 700644 576916 700646
rect 576972 700644 576996 700646
rect 577052 700644 577076 700646
rect 577132 700644 577156 700646
rect 577212 700644 577236 700646
rect 577292 700644 577316 700646
rect 577372 700644 577386 700646
rect 576822 700624 577386 700644
rect 543464 700392 543516 700398
rect 543464 700334 543516 700340
rect 397460 700256 397512 700262
rect 397460 700198 397512 700204
rect 378822 700156 379386 700176
rect 378822 700154 378836 700156
rect 378892 700154 378916 700156
rect 378972 700154 378996 700156
rect 379052 700154 379076 700156
rect 379132 700154 379156 700156
rect 379212 700154 379236 700156
rect 379292 700154 379316 700156
rect 379372 700154 379386 700156
rect 379066 700102 379076 700154
rect 379132 700102 379142 700154
rect 378822 700100 378836 700102
rect 378892 700100 378916 700102
rect 378972 700100 378996 700102
rect 379052 700100 379076 700102
rect 379132 700100 379156 700102
rect 379212 700100 379236 700102
rect 379292 700100 379316 700102
rect 379372 700100 379386 700102
rect 378822 700080 379386 700100
rect 414822 700156 415386 700176
rect 414822 700154 414836 700156
rect 414892 700154 414916 700156
rect 414972 700154 414996 700156
rect 415052 700154 415076 700156
rect 415132 700154 415156 700156
rect 415212 700154 415236 700156
rect 415292 700154 415316 700156
rect 415372 700154 415386 700156
rect 415066 700102 415076 700154
rect 415132 700102 415142 700154
rect 414822 700100 414836 700102
rect 414892 700100 414916 700102
rect 414972 700100 414996 700102
rect 415052 700100 415076 700102
rect 415132 700100 415156 700102
rect 415212 700100 415236 700102
rect 415292 700100 415316 700102
rect 415372 700100 415386 700102
rect 414822 700080 415386 700100
rect 450822 700156 451386 700176
rect 450822 700154 450836 700156
rect 450892 700154 450916 700156
rect 450972 700154 450996 700156
rect 451052 700154 451076 700156
rect 451132 700154 451156 700156
rect 451212 700154 451236 700156
rect 451292 700154 451316 700156
rect 451372 700154 451386 700156
rect 451066 700102 451076 700154
rect 451132 700102 451142 700154
rect 450822 700100 450836 700102
rect 450892 700100 450916 700102
rect 450972 700100 450996 700102
rect 451052 700100 451076 700102
rect 451132 700100 451156 700102
rect 451212 700100 451236 700102
rect 451292 700100 451316 700102
rect 451372 700100 451386 700102
rect 450822 700080 451386 700100
rect 486822 700156 487386 700176
rect 486822 700154 486836 700156
rect 486892 700154 486916 700156
rect 486972 700154 486996 700156
rect 487052 700154 487076 700156
rect 487132 700154 487156 700156
rect 487212 700154 487236 700156
rect 487292 700154 487316 700156
rect 487372 700154 487386 700156
rect 487066 700102 487076 700154
rect 487132 700102 487142 700154
rect 486822 700100 486836 700102
rect 486892 700100 486916 700102
rect 486972 700100 486996 700102
rect 487052 700100 487076 700102
rect 487132 700100 487156 700102
rect 487212 700100 487236 700102
rect 487292 700100 487316 700102
rect 487372 700100 487386 700102
rect 486822 700080 487386 700100
rect 522822 700156 523386 700176
rect 522822 700154 522836 700156
rect 522892 700154 522916 700156
rect 522972 700154 522996 700156
rect 523052 700154 523076 700156
rect 523132 700154 523156 700156
rect 523212 700154 523236 700156
rect 523292 700154 523316 700156
rect 523372 700154 523386 700156
rect 523066 700102 523076 700154
rect 523132 700102 523142 700154
rect 522822 700100 522836 700102
rect 522892 700100 522916 700102
rect 522972 700100 522996 700102
rect 523052 700100 523076 700102
rect 523132 700100 523156 700102
rect 523212 700100 523236 700102
rect 523292 700100 523316 700102
rect 523372 700100 523386 700102
rect 522822 700080 523386 700100
rect 558822 700156 559386 700176
rect 558822 700154 558836 700156
rect 558892 700154 558916 700156
rect 558972 700154 558996 700156
rect 559052 700154 559076 700156
rect 559132 700154 559156 700156
rect 559212 700154 559236 700156
rect 559292 700154 559316 700156
rect 559372 700154 559386 700156
rect 559066 700102 559076 700154
rect 559132 700102 559142 700154
rect 558822 700100 558836 700102
rect 558892 700100 558916 700102
rect 558972 700100 558996 700102
rect 559052 700100 559076 700102
rect 559132 700100 559156 700102
rect 559212 700100 559236 700102
rect 559292 700100 559316 700102
rect 559372 700100 559386 700102
rect 558822 700080 559386 700100
rect 364984 699984 365036 699990
rect 364984 699926 365036 699932
rect 348792 699916 348844 699922
rect 348792 699858 348844 699864
rect 360822 699612 361386 699632
rect 360822 699610 360836 699612
rect 360892 699610 360916 699612
rect 360972 699610 360996 699612
rect 361052 699610 361076 699612
rect 361132 699610 361156 699612
rect 361212 699610 361236 699612
rect 361292 699610 361316 699612
rect 361372 699610 361386 699612
rect 361066 699558 361076 699610
rect 361132 699558 361142 699610
rect 360822 699556 360836 699558
rect 360892 699556 360916 699558
rect 360972 699556 360996 699558
rect 361052 699556 361076 699558
rect 361132 699556 361156 699558
rect 361212 699556 361236 699558
rect 361292 699556 361316 699558
rect 361372 699556 361386 699558
rect 360822 699536 361386 699556
rect 396822 699612 397386 699632
rect 396822 699610 396836 699612
rect 396892 699610 396916 699612
rect 396972 699610 396996 699612
rect 397052 699610 397076 699612
rect 397132 699610 397156 699612
rect 397212 699610 397236 699612
rect 397292 699610 397316 699612
rect 397372 699610 397386 699612
rect 397066 699558 397076 699610
rect 397132 699558 397142 699610
rect 396822 699556 396836 699558
rect 396892 699556 396916 699558
rect 396972 699556 396996 699558
rect 397052 699556 397076 699558
rect 397132 699556 397156 699558
rect 397212 699556 397236 699558
rect 397292 699556 397316 699558
rect 397372 699556 397386 699558
rect 396822 699536 397386 699556
rect 432822 699612 433386 699632
rect 432822 699610 432836 699612
rect 432892 699610 432916 699612
rect 432972 699610 432996 699612
rect 433052 699610 433076 699612
rect 433132 699610 433156 699612
rect 433212 699610 433236 699612
rect 433292 699610 433316 699612
rect 433372 699610 433386 699612
rect 433066 699558 433076 699610
rect 433132 699558 433142 699610
rect 432822 699556 432836 699558
rect 432892 699556 432916 699558
rect 432972 699556 432996 699558
rect 433052 699556 433076 699558
rect 433132 699556 433156 699558
rect 433212 699556 433236 699558
rect 433292 699556 433316 699558
rect 433372 699556 433386 699558
rect 432822 699536 433386 699556
rect 468822 699612 469386 699632
rect 468822 699610 468836 699612
rect 468892 699610 468916 699612
rect 468972 699610 468996 699612
rect 469052 699610 469076 699612
rect 469132 699610 469156 699612
rect 469212 699610 469236 699612
rect 469292 699610 469316 699612
rect 469372 699610 469386 699612
rect 469066 699558 469076 699610
rect 469132 699558 469142 699610
rect 468822 699556 468836 699558
rect 468892 699556 468916 699558
rect 468972 699556 468996 699558
rect 469052 699556 469076 699558
rect 469132 699556 469156 699558
rect 469212 699556 469236 699558
rect 469292 699556 469316 699558
rect 469372 699556 469386 699558
rect 468822 699536 469386 699556
rect 504822 699612 505386 699632
rect 504822 699610 504836 699612
rect 504892 699610 504916 699612
rect 504972 699610 504996 699612
rect 505052 699610 505076 699612
rect 505132 699610 505156 699612
rect 505212 699610 505236 699612
rect 505292 699610 505316 699612
rect 505372 699610 505386 699612
rect 505066 699558 505076 699610
rect 505132 699558 505142 699610
rect 504822 699556 504836 699558
rect 504892 699556 504916 699558
rect 504972 699556 504996 699558
rect 505052 699556 505076 699558
rect 505132 699556 505156 699558
rect 505212 699556 505236 699558
rect 505292 699556 505316 699558
rect 505372 699556 505386 699558
rect 504822 699536 505386 699556
rect 540822 699612 541386 699632
rect 540822 699610 540836 699612
rect 540892 699610 540916 699612
rect 540972 699610 540996 699612
rect 541052 699610 541076 699612
rect 541132 699610 541156 699612
rect 541212 699610 541236 699612
rect 541292 699610 541316 699612
rect 541372 699610 541386 699612
rect 541066 699558 541076 699610
rect 541132 699558 541142 699610
rect 540822 699556 540836 699558
rect 540892 699556 540916 699558
rect 540972 699556 540996 699558
rect 541052 699556 541076 699558
rect 541132 699556 541156 699558
rect 541212 699556 541236 699558
rect 541292 699556 541316 699558
rect 541372 699556 541386 699558
rect 540822 699536 541386 699556
rect 576822 699612 577386 699632
rect 576822 699610 576836 699612
rect 576892 699610 576916 699612
rect 576972 699610 576996 699612
rect 577052 699610 577076 699612
rect 577132 699610 577156 699612
rect 577212 699610 577236 699612
rect 577292 699610 577316 699612
rect 577372 699610 577386 699612
rect 577066 699558 577076 699610
rect 577132 699558 577142 699610
rect 576822 699556 576836 699558
rect 576892 699556 576916 699558
rect 576972 699556 576996 699558
rect 577052 699556 577076 699558
rect 577132 699556 577156 699558
rect 577212 699556 577236 699558
rect 577292 699556 577316 699558
rect 577372 699556 577386 699558
rect 576822 699536 577386 699556
rect 403348 699508 403400 699514
rect 403348 699450 403400 699456
rect 364338 699272 364394 699281
rect 364338 699207 364340 699216
rect 364392 699207 364394 699216
rect 373906 699272 373962 699281
rect 374090 699272 374146 699281
rect 373906 699207 373908 699216
rect 364340 699178 364392 699184
rect 373960 699207 373962 699216
rect 374000 699236 374052 699242
rect 373908 699178 373960 699184
rect 374052 699216 374090 699224
rect 374052 699207 374146 699216
rect 383566 699272 383622 699281
rect 383566 699207 383568 699216
rect 374052 699196 374132 699207
rect 374000 699178 374052 699184
rect 383620 699207 383622 699216
rect 383568 699178 383620 699184
rect 378822 699068 379386 699088
rect 378822 699066 378836 699068
rect 378892 699066 378916 699068
rect 378972 699066 378996 699068
rect 379052 699066 379076 699068
rect 379132 699066 379156 699068
rect 379212 699066 379236 699068
rect 379292 699066 379316 699068
rect 379372 699066 379386 699068
rect 379066 699014 379076 699066
rect 379132 699014 379142 699066
rect 378822 699012 378836 699014
rect 378892 699012 378916 699014
rect 378972 699012 378996 699014
rect 379052 699012 379076 699014
rect 379132 699012 379156 699014
rect 379212 699012 379236 699014
rect 379292 699012 379316 699014
rect 379372 699012 379386 699014
rect 378822 698992 379386 699012
rect 360822 698524 361386 698544
rect 360822 698522 360836 698524
rect 360892 698522 360916 698524
rect 360972 698522 360996 698524
rect 361052 698522 361076 698524
rect 361132 698522 361156 698524
rect 361212 698522 361236 698524
rect 361292 698522 361316 698524
rect 361372 698522 361386 698524
rect 361066 698470 361076 698522
rect 361132 698470 361142 698522
rect 360822 698468 360836 698470
rect 360892 698468 360916 698470
rect 360972 698468 360996 698470
rect 361052 698468 361076 698470
rect 361132 698468 361156 698470
rect 361212 698468 361236 698470
rect 361292 698468 361316 698470
rect 361372 698468 361386 698470
rect 360822 698448 361386 698468
rect 396822 698524 397386 698544
rect 396822 698522 396836 698524
rect 396892 698522 396916 698524
rect 396972 698522 396996 698524
rect 397052 698522 397076 698524
rect 397132 698522 397156 698524
rect 397212 698522 397236 698524
rect 397292 698522 397316 698524
rect 397372 698522 397386 698524
rect 397066 698470 397076 698522
rect 397132 698470 397142 698522
rect 396822 698468 396836 698470
rect 396892 698468 396916 698470
rect 396972 698468 396996 698470
rect 397052 698468 397076 698470
rect 397132 698468 397156 698470
rect 397212 698468 397236 698470
rect 397292 698468 397316 698470
rect 397372 698468 397386 698470
rect 396822 698448 397386 698468
rect 350724 698284 350776 698290
rect 350724 698226 350776 698232
rect 365260 698284 365312 698290
rect 365260 698226 365312 698232
rect 393964 698284 394016 698290
rect 393964 698226 394016 698232
rect 350448 698216 350500 698222
rect 350446 698184 350448 698193
rect 350736 698193 350764 698226
rect 351092 698216 351144 698222
rect 350500 698184 350502 698193
rect 350446 698119 350502 698128
rect 350722 698184 350778 698193
rect 351092 698158 351144 698164
rect 350722 698119 350778 698128
rect 351104 695980 351132 698158
rect 360200 696924 360252 696930
rect 360200 696866 360252 696872
rect 360212 695994 360240 696866
rect 360212 695966 360594 695994
rect 365272 695980 365300 698226
rect 379520 698012 379572 698018
rect 379520 697954 379572 697960
rect 374736 696516 374788 696522
rect 374736 696458 374788 696464
rect 371882 696008 371938 696017
rect 328366 695943 328422 695952
rect 374748 695980 374776 696458
rect 379532 695980 379560 697954
rect 393976 697882 394004 698226
rect 393688 697876 393740 697882
rect 393688 697818 393740 697824
rect 393964 697876 394016 697882
rect 393964 697818 394016 697824
rect 388996 696788 389048 696794
rect 388996 696730 389048 696736
rect 389008 695980 389036 696730
rect 393700 695980 393728 697818
rect 398380 697808 398432 697814
rect 398380 697750 398432 697756
rect 398392 695980 398420 697750
rect 403360 696522 403388 699450
rect 417332 699440 417384 699446
rect 417332 699382 417384 699388
rect 414822 699068 415386 699088
rect 414822 699066 414836 699068
rect 414892 699066 414916 699068
rect 414972 699066 414996 699068
rect 415052 699066 415076 699068
rect 415132 699066 415156 699068
rect 415212 699066 415236 699068
rect 415292 699066 415316 699068
rect 415372 699066 415386 699068
rect 415066 699014 415076 699066
rect 415132 699014 415142 699066
rect 414822 699012 414836 699014
rect 414892 699012 414916 699014
rect 414972 699012 414996 699014
rect 415052 699012 415076 699014
rect 415132 699012 415156 699014
rect 415212 699012 415236 699014
rect 415292 699012 415316 699014
rect 415372 699012 415386 699014
rect 414822 698992 415386 699012
rect 407856 697672 407908 697678
rect 407856 697614 407908 697620
rect 403348 696516 403400 696522
rect 403348 696458 403400 696464
rect 403164 696176 403216 696182
rect 403164 696118 403216 696124
rect 403176 695980 403204 696118
rect 407868 695980 407896 697614
rect 412640 696108 412692 696114
rect 412640 696050 412692 696056
rect 412652 695980 412680 696050
rect 417344 695980 417372 699382
rect 445760 699372 445812 699378
rect 445760 699314 445812 699320
rect 432822 698524 433386 698544
rect 432822 698522 432836 698524
rect 432892 698522 432916 698524
rect 432972 698522 432996 698524
rect 433052 698522 433076 698524
rect 433132 698522 433156 698524
rect 433212 698522 433236 698524
rect 433292 698522 433316 698524
rect 433372 698522 433386 698524
rect 433066 698470 433076 698522
rect 433132 698470 433142 698522
rect 432822 698468 432836 698470
rect 432892 698468 432916 698470
rect 432972 698468 432996 698470
rect 433052 698468 433076 698470
rect 433132 698468 433156 698470
rect 433212 698468 433236 698470
rect 433292 698468 433316 698470
rect 433372 698468 433386 698470
rect 432822 698448 433386 698468
rect 422116 697536 422168 697542
rect 422116 697478 422168 697484
rect 422128 695980 422156 697478
rect 436284 697400 436336 697406
rect 436284 697342 436336 697348
rect 425152 696108 425204 696114
rect 425152 696050 425204 696056
rect 426900 696108 426952 696114
rect 426900 696050 426952 696056
rect 371882 695943 371938 695952
rect 292670 695872 292726 695881
rect 289096 695830 289570 695858
rect 292670 695807 292726 695816
rect 299386 695872 299442 695881
rect 299386 695807 299442 695816
rect 253938 695736 253994 695745
rect 253938 695671 253994 695680
rect 265622 695736 265678 695745
rect 265622 695671 265678 695680
rect 292486 695736 292542 695745
rect 292684 695722 292712 695807
rect 292542 695694 292712 695722
rect 292486 695671 292542 695680
rect 234582 695558 234660 695586
rect 251086 695600 251142 695609
rect 234526 695535 234582 695544
rect 251086 695535 251142 695544
rect 253846 695600 253902 695609
rect 253952 695586 253980 695671
rect 299400 695609 299428 695807
rect 309230 695736 309286 695745
rect 309230 695671 309286 695680
rect 253902 695558 253980 695586
rect 299386 695600 299442 695609
rect 253846 695535 253902 695544
rect 299386 695535 299442 695544
rect 309138 695600 309194 695609
rect 309244 695586 309272 695671
rect 328380 695609 328408 695943
rect 331218 695736 331274 695745
rect 360290 695736 360346 695745
rect 331218 695671 331274 695680
rect 360120 695694 360290 695722
rect 309194 695558 309272 695586
rect 328366 695600 328422 695609
rect 309138 695535 309194 695544
rect 328366 695535 328422 695544
rect 331126 695600 331182 695609
rect 331232 695586 331260 695671
rect 360120 695609 360148 695694
rect 360290 695671 360346 695680
rect 371896 695609 371924 695943
rect 422206 695872 422262 695881
rect 422206 695807 422262 695816
rect 425058 695872 425114 695881
rect 425058 695807 425114 695816
rect 384946 695736 385002 695745
rect 386602 695736 386658 695745
rect 384946 695671 385002 695680
rect 386524 695694 386602 695722
rect 331182 695558 331260 695586
rect 357438 695600 357494 695609
rect 331126 695535 331182 695544
rect 357622 695600 357678 695609
rect 357494 695558 357622 695586
rect 357438 695535 357494 695544
rect 357622 695535 357678 695544
rect 360106 695600 360162 695609
rect 360106 695535 360162 695544
rect 371882 695600 371938 695609
rect 371882 695535 371938 695544
rect 375378 695600 375434 695609
rect 375378 695535 375434 695544
rect 375392 695502 375420 695535
rect 384960 695502 384988 695671
rect 386524 695609 386552 695694
rect 386602 695671 386658 695680
rect 398746 695736 398802 695745
rect 398746 695671 398802 695680
rect 403070 695736 403126 695745
rect 403070 695671 403126 695680
rect 386510 695600 386566 695609
rect 398760 695586 398788 695671
rect 398930 695600 398986 695609
rect 398760 695558 398930 695586
rect 386510 695535 386566 695544
rect 398930 695535 398986 695544
rect 402978 695600 403034 695609
rect 402978 695535 403034 695544
rect 355508 695496 355560 695502
rect 215298 695464 215354 695473
rect 215298 695399 215354 695408
rect 229006 695464 229062 695473
rect 375380 695496 375432 695502
rect 355560 695444 355810 695450
rect 355508 695438 355810 695444
rect 355520 695422 355810 695438
rect 369964 695434 370070 695450
rect 375380 695438 375432 695444
rect 384948 695496 385000 695502
rect 384948 695438 385000 695444
rect 402992 695450 403020 695535
rect 403084 695450 403112 695671
rect 369952 695428 370070 695434
rect 229006 695399 229062 695408
rect 370004 695422 370070 695428
rect 402992 695422 403112 695450
rect 369952 695370 370004 695376
rect 383844 695360 383896 695366
rect 15382 695328 15438 695337
rect 15042 695286 15382 695314
rect 157062 695328 157118 695337
rect 29210 695298 29592 695314
rect 43470 695298 43760 695314
rect 67114 695298 67496 695314
rect 86066 695298 86448 695314
rect 95542 695298 95832 695314
rect 109710 695298 110000 695314
rect 123878 695298 124168 695314
rect 128662 695298 128952 695314
rect 138138 695298 138520 695314
rect 29210 695292 29604 695298
rect 29210 695286 29552 695292
rect 15382 695263 15438 695272
rect 43470 695292 43772 695298
rect 43470 695286 43720 695292
rect 29552 695234 29604 695240
rect 67114 695292 67508 695298
rect 67114 695286 67456 695292
rect 43720 695234 43772 695240
rect 86066 695292 86460 695298
rect 86066 695286 86408 695292
rect 67456 695234 67508 695240
rect 95542 695292 95844 695298
rect 95542 695286 95792 695292
rect 86408 695234 86460 695240
rect 109710 695292 110012 695298
rect 109710 695286 109960 695292
rect 95792 695234 95844 695240
rect 123878 695292 124180 695298
rect 123878 695286 124128 695292
rect 109960 695234 110012 695240
rect 128662 695292 128964 695298
rect 128662 695286 128912 695292
rect 124128 695234 124180 695240
rect 138138 695292 138532 695298
rect 138138 695286 138480 695292
rect 128912 695234 128964 695240
rect 156998 695286 157062 695314
rect 171258 695298 171640 695314
rect 185426 695298 185808 695314
rect 199686 695298 199976 695314
rect 422220 695337 422248 695807
rect 425072 695722 425100 695807
rect 425164 695722 425192 696050
rect 425072 695694 425192 695722
rect 426912 695609 426940 696050
rect 431316 696040 431368 696046
rect 431368 695988 431618 695994
rect 431316 695982 431618 695988
rect 431328 695966 431618 695982
rect 436296 695980 436324 697342
rect 445772 695980 445800 699314
rect 579344 699304 579396 699310
rect 526258 699272 526314 699281
rect 579344 699246 579396 699252
rect 526258 699207 526314 699216
rect 579252 699236 579304 699242
rect 459928 699168 459980 699174
rect 459928 699110 459980 699116
rect 450822 699068 451386 699088
rect 450822 699066 450836 699068
rect 450892 699066 450916 699068
rect 450972 699066 450996 699068
rect 451052 699066 451076 699068
rect 451132 699066 451156 699068
rect 451212 699066 451236 699068
rect 451292 699066 451316 699068
rect 451372 699066 451386 699068
rect 451066 699014 451076 699066
rect 451132 699014 451142 699066
rect 450822 699012 450836 699014
rect 450892 699012 450916 699014
rect 450972 699012 450996 699014
rect 451052 699012 451076 699014
rect 451132 699012 451156 699014
rect 451212 699012 451236 699014
rect 451292 699012 451316 699014
rect 451372 699012 451386 699014
rect 450822 698992 451386 699012
rect 455236 697332 455288 697338
rect 455236 697274 455288 697280
rect 450096 695978 450478 695994
rect 455248 695980 455276 697274
rect 459940 695980 459968 699110
rect 486822 699068 487386 699088
rect 486822 699066 486836 699068
rect 486892 699066 486916 699068
rect 486972 699066 486996 699068
rect 487052 699066 487076 699068
rect 487132 699066 487156 699068
rect 487212 699066 487236 699068
rect 487292 699066 487316 699068
rect 487372 699066 487386 699068
rect 487066 699014 487076 699066
rect 487132 699014 487142 699066
rect 486822 699012 486836 699014
rect 486892 699012 486916 699014
rect 486972 699012 486996 699014
rect 487052 699012 487076 699014
rect 487132 699012 487156 699014
rect 487212 699012 487236 699014
rect 487292 699012 487316 699014
rect 487372 699012 487386 699014
rect 486822 698992 487386 699012
rect 522822 699068 523386 699088
rect 522822 699066 522836 699068
rect 522892 699066 522916 699068
rect 522972 699066 522996 699068
rect 523052 699066 523076 699068
rect 523132 699066 523156 699068
rect 523212 699066 523236 699068
rect 523292 699066 523316 699068
rect 523372 699066 523386 699068
rect 523066 699014 523076 699066
rect 523132 699014 523142 699066
rect 522822 699012 522836 699014
rect 522892 699012 522916 699014
rect 522972 699012 522996 699014
rect 523052 699012 523076 699014
rect 523132 699012 523156 699014
rect 523212 699012 523236 699014
rect 523292 699012 523316 699014
rect 523372 699012 523386 699014
rect 522822 698992 523386 699012
rect 474188 698828 474240 698834
rect 474188 698770 474240 698776
rect 468822 698524 469386 698544
rect 468822 698522 468836 698524
rect 468892 698522 468916 698524
rect 468972 698522 468996 698524
rect 469052 698522 469076 698524
rect 469132 698522 469156 698524
rect 469212 698522 469236 698524
rect 469292 698522 469316 698524
rect 469372 698522 469386 698524
rect 469066 698470 469076 698522
rect 469132 698470 469142 698522
rect 468822 698468 468836 698470
rect 468892 698468 468916 698470
rect 468972 698468 468996 698470
rect 469052 698468 469076 698470
rect 469132 698468 469156 698470
rect 469212 698468 469236 698470
rect 469292 698468 469316 698470
rect 469372 698468 469386 698470
rect 468822 698448 469386 698468
rect 464712 697264 464764 697270
rect 464712 697206 464764 697212
rect 464724 695980 464752 697206
rect 468482 696008 468538 696017
rect 450084 695972 450478 695978
rect 450136 695966 450478 695972
rect 474200 695980 474228 698770
rect 516782 698728 516838 698737
rect 516782 698663 516838 698672
rect 502524 698624 502576 698630
rect 502524 698566 502576 698572
rect 493048 697196 493100 697202
rect 493048 697138 493100 697144
rect 482926 696008 482982 696017
rect 468482 695943 468538 695952
rect 493060 695980 493088 697138
rect 502536 695980 502564 698566
rect 504822 698524 505386 698544
rect 504822 698522 504836 698524
rect 504892 698522 504916 698524
rect 504972 698522 504996 698524
rect 505052 698522 505076 698524
rect 505132 698522 505156 698524
rect 505212 698522 505236 698524
rect 505292 698522 505316 698524
rect 505372 698522 505386 698524
rect 505066 698470 505076 698522
rect 505132 698470 505142 698522
rect 504822 698468 504836 698470
rect 504892 698468 504916 698470
rect 504972 698468 504996 698470
rect 505052 698468 505076 698470
rect 505132 698468 505156 698470
rect 505212 698468 505236 698470
rect 505292 698468 505316 698470
rect 505372 698468 505386 698470
rect 504822 698448 505386 698468
rect 516796 695980 516824 698663
rect 526272 695980 526300 699207
rect 579252 699178 579304 699184
rect 558822 699068 559386 699088
rect 558822 699066 558836 699068
rect 558892 699066 558916 699068
rect 558972 699066 558996 699068
rect 559052 699066 559076 699068
rect 559132 699066 559156 699068
rect 559212 699066 559236 699068
rect 559292 699066 559316 699068
rect 559372 699066 559386 699068
rect 559066 699014 559076 699066
rect 559132 699014 559142 699066
rect 558822 699012 558836 699014
rect 558892 699012 558916 699014
rect 558972 699012 558996 699014
rect 559052 699012 559076 699014
rect 559132 699012 559156 699014
rect 559212 699012 559236 699014
rect 559292 699012 559316 699014
rect 559372 699012 559386 699014
rect 558822 698992 559386 699012
rect 579160 698964 579212 698970
rect 579160 698906 579212 698912
rect 577780 698896 577832 698902
rect 545118 698864 545174 698873
rect 577780 698838 577832 698844
rect 545118 698799 545174 698808
rect 540822 698524 541386 698544
rect 540822 698522 540836 698524
rect 540892 698522 540916 698524
rect 540972 698522 540996 698524
rect 541052 698522 541076 698524
rect 541132 698522 541156 698524
rect 541212 698522 541236 698524
rect 541292 698522 541316 698524
rect 541372 698522 541386 698524
rect 541066 698470 541076 698522
rect 541132 698470 541142 698522
rect 540822 698468 540836 698470
rect 540892 698468 540916 698470
rect 540972 698468 540996 698470
rect 541052 698468 541076 698470
rect 541132 698468 541156 698470
rect 541212 698468 541236 698470
rect 541292 698468 541316 698470
rect 541372 698468 541386 698470
rect 540822 698448 541386 698468
rect 535644 697128 535696 697134
rect 535644 697070 535696 697076
rect 540426 697096 540482 697105
rect 535656 695980 535684 697070
rect 540426 697031 540482 697040
rect 540440 695980 540468 697031
rect 545132 695980 545160 698799
rect 576822 698524 577386 698544
rect 576822 698522 576836 698524
rect 576892 698522 576916 698524
rect 576972 698522 576996 698524
rect 577052 698522 577076 698524
rect 577132 698522 577156 698524
rect 577212 698522 577236 698524
rect 577292 698522 577316 698524
rect 577372 698522 577386 698524
rect 577066 698470 577076 698522
rect 577132 698470 577142 698522
rect 576822 698468 576836 698470
rect 576892 698468 576916 698470
rect 576972 698468 576996 698470
rect 577052 698468 577076 698470
rect 577132 698468 577156 698470
rect 577212 698468 577236 698470
rect 577292 698468 577316 698470
rect 577372 698468 577386 698470
rect 576822 698448 577386 698468
rect 577596 698352 577648 698358
rect 577596 698294 577648 698300
rect 576032 698148 576084 698154
rect 576032 698090 576084 698096
rect 574652 697944 574704 697950
rect 574652 697886 574704 697892
rect 482926 695943 482982 695952
rect 450084 695914 450136 695920
rect 437294 695872 437350 695881
rect 437478 695872 437534 695881
rect 437350 695830 437478 695858
rect 437294 695807 437350 695816
rect 437478 695807 437534 695816
rect 452566 695736 452622 695745
rect 452566 695671 452622 695680
rect 426530 695600 426586 695609
rect 426898 695600 426954 695609
rect 426586 695558 426834 695586
rect 426530 695535 426586 695544
rect 426898 695535 426954 695544
rect 452580 695473 452608 695671
rect 468496 695609 468524 695943
rect 469220 695904 469272 695910
rect 469272 695852 469430 695858
rect 469220 695846 469430 695852
rect 469232 695830 469430 695846
rect 478800 695842 478906 695858
rect 478788 695836 478906 695842
rect 478840 695830 478906 695836
rect 478788 695778 478840 695784
rect 482940 695745 482968 695943
rect 485780 695836 485832 695842
rect 485780 695778 485832 695784
rect 492588 695836 492640 695842
rect 492588 695778 492640 695784
rect 485792 695745 485820 695778
rect 487988 695768 488040 695774
rect 482926 695736 482982 695745
rect 482926 695671 482982 695680
rect 485778 695736 485834 695745
rect 488040 695716 488382 695722
rect 487988 695710 488382 695716
rect 488000 695694 488382 695710
rect 485778 695671 485834 695680
rect 492600 695609 492628 695778
rect 562324 695768 562376 695774
rect 543830 695736 543886 695745
rect 506952 695706 507334 695722
rect 506940 695700 507334 695706
rect 506992 695694 507334 695700
rect 540980 695700 541032 695706
rect 506940 695642 506992 695648
rect 543830 695671 543832 695680
rect 540980 695642 541032 695648
rect 543884 695671 543886 695680
rect 553214 695736 553270 695745
rect 553398 695736 553454 695745
rect 553270 695694 553398 695722
rect 553214 695671 553270 695680
rect 553398 695671 553454 695680
rect 562322 695736 562324 695745
rect 567108 695768 567160 695774
rect 562376 695736 562378 695745
rect 562322 695671 562378 695680
rect 567106 695736 567108 695745
rect 567160 695736 567162 695745
rect 567106 695671 567162 695680
rect 569314 695736 569370 695745
rect 569314 695671 569370 695680
rect 543832 695642 543884 695648
rect 540992 695609 541020 695642
rect 468482 695600 468538 695609
rect 468482 695535 468538 695544
rect 492586 695600 492642 695609
rect 540978 695600 541034 695609
rect 530688 695570 530978 695586
rect 492586 695535 492642 695544
rect 530676 695564 530978 695570
rect 530728 695558 530978 695564
rect 540978 695535 541034 695544
rect 530676 695506 530728 695512
rect 452566 695464 452622 695473
rect 452566 695399 452622 695408
rect 440700 695360 440752 695366
rect 422206 695328 422262 695337
rect 383896 695308 384238 695314
rect 383844 695302 384238 695308
rect 171258 695292 171652 695298
rect 171258 695286 171600 695292
rect 157062 695263 157118 695272
rect 138480 695234 138532 695240
rect 185426 695292 185820 695298
rect 185426 695286 185768 695292
rect 171600 695234 171652 695240
rect 199686 695292 199988 695298
rect 199686 695286 199936 695292
rect 185768 695234 185820 695240
rect 383856 695286 384238 695302
rect 483388 695360 483440 695366
rect 440752 695308 441002 695314
rect 440700 695302 441002 695308
rect 497556 695360 497608 695366
rect 483440 695308 483690 695314
rect 483388 695302 483690 695308
rect 511908 695360 511960 695366
rect 497608 695308 497858 695314
rect 497556 695302 497858 695308
rect 521382 695328 521438 695337
rect 511960 695308 512026 695314
rect 511908 695302 512026 695308
rect 440712 695286 441002 695302
rect 483400 695286 483690 695302
rect 497568 695286 497858 695302
rect 511920 695286 512026 695302
rect 422206 695263 422262 695272
rect 521438 695286 521502 695314
rect 521382 695263 521438 695272
rect 199936 695234 199988 695240
rect 569328 694754 569356 695671
rect 569316 694748 569368 694754
rect 569316 694690 569368 694696
rect 568486 693832 568542 693841
rect 568486 693767 568542 693776
rect 568500 693433 568528 693767
rect 568486 693424 568542 693433
rect 568486 693359 568542 693368
rect 574664 628017 574692 697886
rect 575388 697740 575440 697746
rect 575388 697682 575440 697688
rect 575296 697604 575348 697610
rect 575296 697546 575348 697552
rect 575204 697468 575256 697474
rect 575204 697410 575256 697416
rect 574928 697060 574980 697066
rect 574928 697002 574980 697008
rect 574836 696992 574888 696998
rect 574742 696960 574798 696969
rect 574836 696934 574888 696940
rect 574742 696895 574798 696904
rect 574650 628008 574706 628017
rect 574650 627943 574706 627952
rect 8208 423904 8260 423910
rect 8208 423846 8260 423852
rect 8116 308916 8168 308922
rect 8116 308858 8168 308864
rect 8024 208208 8076 208214
rect 8024 208150 8076 208156
rect 7932 165096 7984 165102
rect 7932 165038 7984 165044
rect 7840 136400 7892 136406
rect 7840 136342 7892 136348
rect 7748 122188 7800 122194
rect 7748 122130 7800 122136
rect 7656 79892 7708 79898
rect 7656 79834 7708 79840
rect 7564 35828 7616 35834
rect 7564 35770 7616 35776
rect 574756 17762 574784 696895
rect 574848 66178 574876 696934
rect 574940 111790 574968 697002
rect 575020 695632 575072 695638
rect 575020 695574 575072 695580
rect 575032 158710 575060 695574
rect 575112 694408 575164 694414
rect 575112 694350 575164 694356
rect 575124 205562 575152 694350
rect 575216 487150 575244 697410
rect 575308 534070 575336 697546
rect 575400 580922 575428 697682
rect 576044 674830 576072 698090
rect 577412 695292 577464 695298
rect 577412 695234 577464 695240
rect 576768 695020 576820 695026
rect 576768 694962 576820 694968
rect 576676 694884 576728 694890
rect 576676 694826 576728 694832
rect 576584 694816 576636 694822
rect 576584 694758 576636 694764
rect 576492 694680 576544 694686
rect 576492 694622 576544 694628
rect 576400 694476 576452 694482
rect 576400 694418 576452 694424
rect 576122 694376 576178 694385
rect 576122 694311 576178 694320
rect 576032 674824 576084 674830
rect 576032 674766 576084 674772
rect 575478 628008 575534 628017
rect 575478 627943 575534 627952
rect 575492 627910 575520 627943
rect 575480 627904 575532 627910
rect 575480 627846 575532 627852
rect 575388 580916 575440 580922
rect 575388 580858 575440 580864
rect 575296 534064 575348 534070
rect 575296 534006 575348 534012
rect 575204 487144 575256 487150
rect 575204 487086 575256 487092
rect 575112 205556 575164 205562
rect 575112 205498 575164 205504
rect 575020 158704 575072 158710
rect 575020 158646 575072 158652
rect 574928 111784 574980 111790
rect 574928 111726 574980 111732
rect 574848 66150 574968 66178
rect 574940 64870 574968 66150
rect 574928 64864 574980 64870
rect 574928 64806 574980 64812
rect 576136 41274 576164 694311
rect 576308 694272 576360 694278
rect 576308 694214 576360 694220
rect 576216 694204 576268 694210
rect 576216 694146 576268 694152
rect 576228 88330 576256 694146
rect 576320 135250 576348 694214
rect 576412 252550 576440 694418
rect 576504 299470 576532 694622
rect 576596 346390 576624 694758
rect 576688 393242 576716 694826
rect 576780 440230 576808 694962
rect 577424 651370 577452 695234
rect 577504 694748 577556 694754
rect 577504 694690 577556 694696
rect 577412 651364 577464 651370
rect 577412 651306 577464 651312
rect 576768 440224 576820 440230
rect 576768 440166 576820 440172
rect 576676 393236 576728 393242
rect 576676 393178 576728 393184
rect 576584 346384 576636 346390
rect 576584 346326 576636 346332
rect 576492 299464 576544 299470
rect 576492 299406 576544 299412
rect 576400 252544 576452 252550
rect 576400 252486 576452 252492
rect 576308 135244 576360 135250
rect 576308 135186 576360 135192
rect 576216 88324 576268 88330
rect 576216 88266 576268 88272
rect 576124 41268 576176 41274
rect 576124 41210 576176 41216
rect 577516 30326 577544 694690
rect 577608 170678 577636 698294
rect 577688 694544 577740 694550
rect 577688 694486 577740 694492
rect 577700 276010 577728 694486
rect 577792 369850 577820 698838
rect 579068 698760 579120 698766
rect 579068 698702 579120 698708
rect 578976 698692 579028 698698
rect 578976 698634 579028 698640
rect 578884 698420 578936 698426
rect 578884 698362 578936 698368
rect 578700 696720 578752 696726
rect 578700 696662 578752 696668
rect 578148 695360 578200 695366
rect 578148 695302 578200 695308
rect 578056 695156 578108 695162
rect 578056 695098 578108 695104
rect 577872 694952 577924 694958
rect 577872 694894 577924 694900
rect 577884 416634 577912 694894
rect 577962 693968 578018 693977
rect 577962 693903 578018 693912
rect 577976 510610 578004 693903
rect 578068 557394 578096 695098
rect 578160 604314 578188 695302
rect 578712 687206 578740 696662
rect 578792 696448 578844 696454
rect 578792 696390 578844 696396
rect 578700 687200 578752 687206
rect 578700 687142 578752 687148
rect 578804 640218 578832 696390
rect 578792 640212 578844 640218
rect 578792 640154 578844 640160
rect 578148 604308 578200 604314
rect 578148 604250 578200 604256
rect 578056 557388 578108 557394
rect 578056 557330 578108 557336
rect 577964 510604 578016 510610
rect 577964 510546 578016 510552
rect 577872 416628 577924 416634
rect 577872 416570 577924 416576
rect 577780 369844 577832 369850
rect 577780 369786 577832 369792
rect 577688 276004 577740 276010
rect 577688 275946 577740 275952
rect 578896 217025 578924 698362
rect 578988 263945 579016 698634
rect 579080 310865 579108 698702
rect 579172 357921 579200 698906
rect 579264 451761 579292 699178
rect 579356 498681 579384 699246
rect 580540 698216 580592 698222
rect 580540 698158 580592 698164
rect 579620 698080 579672 698086
rect 579618 698048 579620 698057
rect 579672 698048 579674 698057
rect 579618 697983 579674 697992
rect 580356 696584 580408 696590
rect 580356 696526 580408 696532
rect 579528 696176 579580 696182
rect 579528 696118 579580 696124
rect 580262 696144 580318 696153
rect 579434 693560 579490 693569
rect 579434 693495 579490 693504
rect 579448 545601 579476 693495
rect 579540 592521 579568 696118
rect 580262 696079 580318 696088
rect 579804 674824 579856 674830
rect 579804 674766 579856 674772
rect 579816 674665 579844 674766
rect 579802 674656 579858 674665
rect 579802 674591 579858 674600
rect 579620 651364 579672 651370
rect 579620 651306 579672 651312
rect 579632 651137 579660 651306
rect 579618 651128 579674 651137
rect 579618 651063 579674 651072
rect 579804 627904 579856 627910
rect 579804 627846 579856 627852
rect 579816 627745 579844 627846
rect 579802 627736 579858 627745
rect 579802 627671 579858 627680
rect 579620 604308 579672 604314
rect 579620 604250 579672 604256
rect 579632 604217 579660 604250
rect 579618 604208 579674 604217
rect 579618 604143 579674 604152
rect 579526 592512 579582 592521
rect 579526 592447 579582 592456
rect 580172 580916 580224 580922
rect 580172 580858 580224 580864
rect 580184 580825 580212 580858
rect 580170 580816 580226 580825
rect 580170 580751 580226 580760
rect 579620 557388 579672 557394
rect 579620 557330 579672 557336
rect 579632 557297 579660 557330
rect 579618 557288 579674 557297
rect 579618 557223 579674 557232
rect 579434 545592 579490 545601
rect 579434 545527 579490 545536
rect 579804 534064 579856 534070
rect 579804 534006 579856 534012
rect 579816 533905 579844 534006
rect 579802 533896 579858 533905
rect 579802 533831 579858 533840
rect 580080 510604 580132 510610
rect 580080 510546 580132 510552
rect 580092 510377 580120 510546
rect 580078 510368 580134 510377
rect 580078 510303 580134 510312
rect 579342 498672 579398 498681
rect 579342 498607 579398 498616
rect 580172 487144 580224 487150
rect 580172 487086 580224 487092
rect 580184 486849 580212 487086
rect 580170 486840 580226 486849
rect 580170 486775 580226 486784
rect 579250 451752 579306 451761
rect 579250 451687 579306 451696
rect 579988 440224 580040 440230
rect 579988 440166 580040 440172
rect 580000 439929 580028 440166
rect 579986 439920 580042 439929
rect 579986 439855 580042 439864
rect 579620 416628 579672 416634
rect 579620 416570 579672 416576
rect 579632 416537 579660 416570
rect 579618 416528 579674 416537
rect 579618 416463 579674 416472
rect 579620 393236 579672 393242
rect 579620 393178 579672 393184
rect 579632 393009 579660 393178
rect 579618 393000 579674 393009
rect 579618 392935 579674 392944
rect 579158 357912 579214 357921
rect 579158 357847 579214 357856
rect 580172 346384 580224 346390
rect 580172 346326 580224 346332
rect 580184 346089 580212 346326
rect 580170 346080 580226 346089
rect 580170 346015 580226 346024
rect 579066 310856 579122 310865
rect 579066 310791 579122 310800
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 299169 580212 299406
rect 580170 299160 580226 299169
rect 580170 299095 580226 299104
rect 579620 276004 579672 276010
rect 579620 275946 579672 275952
rect 579632 275777 579660 275946
rect 579618 275768 579674 275777
rect 579618 275703 579674 275712
rect 578974 263936 579030 263945
rect 578974 263871 579030 263880
rect 580172 252544 580224 252550
rect 580172 252486 580224 252492
rect 580184 252249 580212 252486
rect 580170 252240 580226 252249
rect 580170 252175 580226 252184
rect 578882 217016 578938 217025
rect 578882 216951 578938 216960
rect 580172 205556 580224 205562
rect 580172 205498 580224 205504
rect 580184 205329 580212 205498
rect 580170 205320 580226 205329
rect 580170 205255 580226 205264
rect 577596 170672 577648 170678
rect 577596 170614 577648 170620
rect 579620 158704 579672 158710
rect 579620 158646 579672 158652
rect 579632 158409 579660 158646
rect 579618 158400 579674 158409
rect 579618 158335 579674 158344
rect 580172 135244 580224 135250
rect 580172 135186 580224 135192
rect 580184 134881 580212 135186
rect 580170 134872 580226 134881
rect 580170 134807 580226 134816
rect 580172 111784 580224 111790
rect 580172 111726 580224 111732
rect 580184 111489 580212 111726
rect 580170 111480 580226 111489
rect 580170 111415 580226 111424
rect 579896 88324 579948 88330
rect 579896 88266 579948 88272
rect 579908 87961 579936 88266
rect 579894 87952 579950 87961
rect 579894 87887 579950 87896
rect 580276 76265 580304 696079
rect 580368 123185 580396 696526
rect 580448 696244 580500 696250
rect 580448 696186 580500 696192
rect 580460 181937 580488 696186
rect 580552 228857 580580 698158
rect 580632 697876 580684 697882
rect 580632 697818 580684 697824
rect 580644 322697 580672 697818
rect 580724 696652 580776 696658
rect 580724 696594 580776 696600
rect 580736 404841 580764 696594
rect 580816 696516 580868 696522
rect 580816 696458 580868 696464
rect 580828 463457 580856 696458
rect 580908 687200 580960 687206
rect 580908 687142 580960 687148
rect 580920 686361 580948 687142
rect 580906 686352 580962 686361
rect 580906 686287 580962 686296
rect 580908 640212 580960 640218
rect 580908 640154 580960 640160
rect 580920 639441 580948 640154
rect 580906 639432 580962 639441
rect 580906 639367 580962 639376
rect 580814 463448 580870 463457
rect 580814 463383 580870 463392
rect 580722 404832 580778 404841
rect 580722 404767 580778 404776
rect 580724 369844 580776 369850
rect 580724 369786 580776 369792
rect 580736 369617 580764 369786
rect 580722 369608 580778 369617
rect 580722 369543 580778 369552
rect 580630 322688 580686 322697
rect 580630 322623 580686 322632
rect 580538 228848 580594 228857
rect 580538 228783 580594 228792
rect 580446 181928 580502 181937
rect 580446 181863 580502 181872
rect 580632 170672 580684 170678
rect 580632 170614 580684 170620
rect 580644 170105 580672 170614
rect 580630 170096 580686 170105
rect 580630 170031 580686 170040
rect 580354 123176 580410 123185
rect 580354 123111 580410 123120
rect 580262 76256 580318 76265
rect 580262 76191 580318 76200
rect 579804 64864 579856 64870
rect 579804 64806 579856 64812
rect 579816 64569 579844 64806
rect 579802 64560 579858 64569
rect 579802 64495 579858 64504
rect 580172 41268 580224 41274
rect 580172 41210 580224 41216
rect 580184 41041 580212 41210
rect 580170 41032 580226 41041
rect 580170 40967 580226 40976
rect 577504 30320 577556 30326
rect 577504 30262 577556 30268
rect 579620 30320 579672 30326
rect 579620 30262 579672 30268
rect 579632 29345 579660 30262
rect 579618 29336 579674 29345
rect 579618 29271 579674 29280
rect 575020 17876 575072 17882
rect 575020 17818 575072 17824
rect 580172 17876 580224 17882
rect 580172 17818 580224 17824
rect 575032 17762 575060 17818
rect 574756 17734 575060 17762
rect 580184 17649 580212 17818
rect 580170 17640 580226 17649
rect 580170 17575 580226 17584
rect 3148 7200 3200 7206
rect 3146 7168 3148 7177
rect 6184 7200 6236 7206
rect 3200 7168 3202 7177
rect 6184 7142 6236 7148
rect 3146 7103 3202 7112
rect 5540 6180 5592 6186
rect 5540 6122 5592 6128
rect 572 4072 624 4078
rect 572 4014 624 4020
rect 584 480 612 4014
rect 5264 3596 5316 3602
rect 5264 3538 5316 3544
rect 4068 3460 4120 3466
rect 4068 3402 4120 3408
rect 2872 3120 2924 3126
rect 2872 3062 2924 3068
rect 1676 2916 1728 2922
rect 1676 2858 1728 2864
rect 1688 480 1716 2858
rect 2884 480 2912 3062
rect 4080 480 4108 3402
rect 5276 480 5304 3538
rect 5552 3126 5580 6122
rect 8588 4078 8616 8092
rect 9692 5658 9720 8092
rect 10796 6186 10824 8092
rect 11624 8078 11914 8106
rect 12452 8078 13110 8106
rect 10784 6180 10836 6186
rect 10784 6122 10836 6128
rect 9600 5630 9720 5658
rect 8576 4072 8628 4078
rect 8576 4014 8628 4020
rect 6460 3936 6512 3942
rect 6460 3878 6512 3884
rect 5540 3120 5592 3126
rect 5540 3062 5592 3068
rect 6472 480 6500 3878
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 7668 480 7696 3470
rect 8852 3392 8904 3398
rect 8852 3334 8904 3340
rect 8864 480 8892 3334
rect 9600 2922 9628 5630
rect 11060 5568 11112 5574
rect 11060 5510 11112 5516
rect 11072 3942 11100 5510
rect 11244 4072 11296 4078
rect 11244 4014 11296 4020
rect 11060 3936 11112 3942
rect 11060 3878 11112 3884
rect 9588 2916 9640 2922
rect 9588 2858 9640 2864
rect 10048 2916 10100 2922
rect 10048 2858 10100 2864
rect 10060 480 10088 2858
rect 11256 480 11284 4014
rect 11624 3466 11652 8078
rect 12452 5658 12480 8078
rect 12268 5630 12480 5658
rect 13820 5636 13872 5642
rect 12268 3602 12296 5630
rect 13820 5578 13872 5584
rect 12256 3596 12308 3602
rect 12256 3538 12308 3544
rect 11612 3460 11664 3466
rect 11612 3402 11664 3408
rect 13832 3398 13860 5578
rect 14200 5574 14228 8092
rect 15212 8078 15318 8106
rect 15212 5794 15240 8078
rect 15028 5766 15240 5794
rect 14188 5568 14240 5574
rect 14188 5510 14240 5516
rect 15028 3534 15056 5766
rect 15200 5704 15252 5710
rect 15200 5646 15252 5652
rect 15016 3528 15068 3534
rect 15016 3470 15068 3476
rect 14832 3460 14884 3466
rect 14832 3402 14884 3408
rect 13820 3392 13872 3398
rect 13820 3334 13872 3340
rect 13636 3188 13688 3194
rect 13636 3130 13688 3136
rect 12440 3052 12492 3058
rect 12440 2994 12492 3000
rect 12452 480 12480 2994
rect 13648 480 13676 3130
rect 14844 480 14872 3402
rect 15212 2922 15240 5646
rect 16500 5642 16528 8092
rect 17604 5710 17632 8092
rect 17592 5704 17644 5710
rect 17592 5646 17644 5652
rect 18604 5704 18656 5710
rect 18604 5646 18656 5652
rect 16488 5636 16540 5642
rect 16488 5578 16540 5584
rect 18052 5636 18104 5642
rect 18052 5578 18104 5584
rect 16948 5568 17000 5574
rect 16948 5510 17000 5516
rect 16960 4078 16988 5510
rect 16948 4072 17000 4078
rect 16948 4014 17000 4020
rect 16028 3596 16080 3602
rect 16028 3538 16080 3544
rect 15200 2916 15252 2922
rect 15200 2858 15252 2864
rect 16040 480 16068 3538
rect 17224 3528 17276 3534
rect 17224 3470 17276 3476
rect 17236 480 17264 3470
rect 18064 3058 18092 5578
rect 18328 3392 18380 3398
rect 18328 3334 18380 3340
rect 18052 3052 18104 3058
rect 18052 2994 18104 3000
rect 18340 480 18368 3334
rect 18616 3194 18644 5646
rect 18708 5574 18736 8092
rect 18822 6012 19386 6032
rect 18822 6010 18836 6012
rect 18892 6010 18916 6012
rect 18972 6010 18996 6012
rect 19052 6010 19076 6012
rect 19132 6010 19156 6012
rect 19212 6010 19236 6012
rect 19292 6010 19316 6012
rect 19372 6010 19386 6012
rect 19066 5958 19076 6010
rect 19132 5958 19142 6010
rect 18822 5956 18836 5958
rect 18892 5956 18916 5958
rect 18972 5956 18996 5958
rect 19052 5956 19076 5958
rect 19132 5956 19156 5958
rect 19212 5956 19236 5958
rect 19292 5956 19316 5958
rect 19372 5956 19386 5958
rect 18822 5936 19386 5956
rect 19904 5642 19932 8092
rect 21008 5710 21036 8092
rect 20996 5704 21048 5710
rect 20996 5646 21048 5652
rect 19892 5636 19944 5642
rect 19892 5578 19944 5584
rect 20720 5636 20772 5642
rect 20720 5578 20772 5584
rect 18696 5568 18748 5574
rect 18696 5510 18748 5516
rect 19432 5568 19484 5574
rect 19432 5510 19484 5516
rect 18822 4924 19386 4944
rect 18822 4922 18836 4924
rect 18892 4922 18916 4924
rect 18972 4922 18996 4924
rect 19052 4922 19076 4924
rect 19132 4922 19156 4924
rect 19212 4922 19236 4924
rect 19292 4922 19316 4924
rect 19372 4922 19386 4924
rect 19066 4870 19076 4922
rect 19132 4870 19142 4922
rect 18822 4868 18836 4870
rect 18892 4868 18916 4870
rect 18972 4868 18996 4870
rect 19052 4868 19076 4870
rect 19132 4868 19156 4870
rect 19212 4868 19236 4870
rect 19292 4868 19316 4870
rect 19372 4868 19386 4870
rect 18822 4848 19386 4868
rect 18822 3836 19386 3856
rect 18822 3834 18836 3836
rect 18892 3834 18916 3836
rect 18972 3834 18996 3836
rect 19052 3834 19076 3836
rect 19132 3834 19156 3836
rect 19212 3834 19236 3836
rect 19292 3834 19316 3836
rect 19372 3834 19386 3836
rect 19066 3782 19076 3834
rect 19132 3782 19142 3834
rect 18822 3780 18836 3782
rect 18892 3780 18916 3782
rect 18972 3780 18996 3782
rect 19052 3780 19076 3782
rect 19132 3780 19156 3782
rect 19212 3780 19236 3782
rect 19292 3780 19316 3782
rect 19372 3780 19386 3782
rect 18822 3760 19386 3780
rect 19444 3466 19472 5510
rect 20732 3602 20760 5578
rect 22112 5574 22140 8092
rect 23112 5704 23164 5710
rect 23112 5646 23164 5652
rect 22100 5568 22152 5574
rect 22100 5510 22152 5516
rect 20812 4140 20864 4146
rect 20812 4082 20864 4088
rect 20720 3596 20772 3602
rect 20720 3538 20772 3544
rect 19432 3460 19484 3466
rect 19432 3402 19484 3408
rect 18604 3188 18656 3194
rect 18604 3130 18656 3136
rect 19524 2848 19576 2854
rect 19524 2790 19576 2796
rect 18822 2748 19386 2768
rect 18822 2746 18836 2748
rect 18892 2746 18916 2748
rect 18972 2746 18996 2748
rect 19052 2746 19076 2748
rect 19132 2746 19156 2748
rect 19212 2746 19236 2748
rect 19292 2746 19316 2748
rect 19372 2746 19386 2748
rect 19066 2694 19076 2746
rect 19132 2694 19142 2746
rect 18822 2692 18836 2694
rect 18892 2692 18916 2694
rect 18972 2692 18996 2694
rect 19052 2692 19076 2694
rect 19132 2692 19156 2694
rect 19212 2692 19236 2694
rect 19292 2692 19316 2694
rect 19372 2692 19386 2694
rect 18822 2672 19386 2692
rect 19536 480 19564 2790
rect 20824 2122 20852 4082
rect 21916 4072 21968 4078
rect 21916 4014 21968 4020
rect 20732 2094 20852 2122
rect 20732 480 20760 2094
rect 21928 480 21956 4014
rect 23124 3534 23152 5646
rect 23308 5642 23336 8092
rect 23848 5772 23900 5778
rect 23848 5714 23900 5720
rect 23296 5636 23348 5642
rect 23296 5578 23348 5584
rect 23112 3528 23164 3534
rect 23112 3470 23164 3476
rect 23860 3398 23888 5714
rect 24412 5710 24440 8092
rect 25516 5778 25544 8092
rect 26252 8078 26726 8106
rect 27632 8078 27830 8106
rect 26252 5794 26280 8078
rect 25504 5772 25556 5778
rect 25504 5714 25556 5720
rect 26160 5766 26280 5794
rect 24400 5704 24452 5710
rect 24400 5646 24452 5652
rect 25504 4004 25556 4010
rect 25504 3946 25556 3952
rect 24308 3936 24360 3942
rect 24308 3878 24360 3884
rect 23848 3392 23900 3398
rect 23848 3334 23900 3340
rect 23112 3188 23164 3194
rect 23112 3130 23164 3136
rect 23124 480 23152 3130
rect 24320 480 24348 3878
rect 25516 480 25544 3946
rect 26160 2854 26188 5766
rect 26240 5704 26292 5710
rect 26240 5646 26292 5652
rect 26252 4078 26280 5646
rect 27632 5556 27660 8078
rect 28920 5710 28948 8092
rect 28908 5704 28960 5710
rect 28908 5646 28960 5652
rect 30116 5642 30144 8092
rect 27712 5636 27764 5642
rect 27712 5578 27764 5584
rect 30104 5636 30156 5642
rect 30104 5578 30156 5584
rect 27540 5528 27660 5556
rect 27540 4146 27568 5528
rect 27528 4140 27580 4146
rect 27528 4082 27580 4088
rect 26240 4072 26292 4078
rect 26240 4014 26292 4020
rect 26700 3528 26752 3534
rect 26700 3470 26752 3476
rect 26148 2848 26200 2854
rect 26148 2790 26200 2796
rect 26712 480 26740 3470
rect 27724 3194 27752 5578
rect 31220 5574 31248 8092
rect 31772 8078 32338 8106
rect 33152 8078 33534 8106
rect 34532 8078 34638 8106
rect 31772 5658 31800 8078
rect 31680 5630 31800 5658
rect 29000 5568 29052 5574
rect 29000 5510 29052 5516
rect 31208 5568 31260 5574
rect 31208 5510 31260 5516
rect 29012 3942 29040 5510
rect 31484 4072 31536 4078
rect 31484 4014 31536 4020
rect 29000 3936 29052 3942
rect 29000 3878 29052 3884
rect 29092 3664 29144 3670
rect 29092 3606 29144 3612
rect 27896 3460 27948 3466
rect 27896 3402 27948 3408
rect 27712 3188 27764 3194
rect 27712 3130 27764 3136
rect 27908 480 27936 3402
rect 29104 480 29132 3606
rect 30288 2848 30340 2854
rect 30288 2790 30340 2796
rect 30300 480 30328 2790
rect 31496 480 31524 4014
rect 31680 4010 31708 5630
rect 33152 5574 33180 8078
rect 34532 5794 34560 8078
rect 34348 5766 34560 5794
rect 31760 5568 31812 5574
rect 31760 5510 31812 5516
rect 33140 5568 33192 5574
rect 33140 5510 33192 5516
rect 31668 4004 31720 4010
rect 31668 3946 31720 3952
rect 31772 3534 31800 5510
rect 31760 3528 31812 3534
rect 31760 3470 31812 3476
rect 33876 3528 33928 3534
rect 33876 3470 33928 3476
rect 32680 3120 32732 3126
rect 32680 3062 32732 3068
rect 32692 480 32720 3062
rect 33888 480 33916 3470
rect 34348 3466 34376 5766
rect 34520 5636 34572 5642
rect 34520 5578 34572 5584
rect 34336 3460 34388 3466
rect 34336 3402 34388 3408
rect 34532 2854 34560 5578
rect 35728 3670 35756 8092
rect 36924 5642 36952 8092
rect 36912 5636 36964 5642
rect 36912 5578 36964 5584
rect 37464 5636 37516 5642
rect 37464 5578 37516 5584
rect 36452 5568 36504 5574
rect 36452 5510 36504 5516
rect 36464 4078 36492 5510
rect 36822 5468 37386 5488
rect 36822 5466 36836 5468
rect 36892 5466 36916 5468
rect 36972 5466 36996 5468
rect 37052 5466 37076 5468
rect 37132 5466 37156 5468
rect 37212 5466 37236 5468
rect 37292 5466 37316 5468
rect 37372 5466 37386 5468
rect 37066 5414 37076 5466
rect 37132 5414 37142 5466
rect 36822 5412 36836 5414
rect 36892 5412 36916 5414
rect 36972 5412 36996 5414
rect 37052 5412 37076 5414
rect 37132 5412 37156 5414
rect 37212 5412 37236 5414
rect 37292 5412 37316 5414
rect 37372 5412 37386 5414
rect 36822 5392 37386 5412
rect 36822 4380 37386 4400
rect 36822 4378 36836 4380
rect 36892 4378 36916 4380
rect 36972 4378 36996 4380
rect 37052 4378 37076 4380
rect 37132 4378 37156 4380
rect 37212 4378 37236 4380
rect 37292 4378 37316 4380
rect 37372 4378 37386 4380
rect 37066 4326 37076 4378
rect 37132 4326 37142 4378
rect 36822 4324 36836 4326
rect 36892 4324 36916 4326
rect 36972 4324 36996 4326
rect 37052 4324 37076 4326
rect 37132 4324 37156 4326
rect 37212 4324 37236 4326
rect 37292 4324 37316 4326
rect 37372 4324 37386 4326
rect 36822 4304 37386 4324
rect 36452 4072 36504 4078
rect 36452 4014 36504 4020
rect 35716 3664 35768 3670
rect 35716 3606 35768 3612
rect 34980 3596 35032 3602
rect 34980 3538 35032 3544
rect 34520 2848 34572 2854
rect 34520 2790 34572 2796
rect 34992 480 35020 3538
rect 36176 3392 36228 3398
rect 36176 3334 36228 3340
rect 36188 480 36216 3334
rect 36822 3292 37386 3312
rect 36822 3290 36836 3292
rect 36892 3290 36916 3292
rect 36972 3290 36996 3292
rect 37052 3290 37076 3292
rect 37132 3290 37156 3292
rect 37212 3290 37236 3292
rect 37292 3290 37316 3292
rect 37372 3290 37386 3292
rect 37066 3238 37076 3290
rect 37132 3238 37142 3290
rect 36822 3236 36836 3238
rect 36892 3236 36916 3238
rect 36972 3236 36996 3238
rect 37052 3236 37076 3238
rect 37132 3236 37156 3238
rect 37212 3236 37236 3238
rect 37292 3236 37316 3238
rect 37372 3236 37386 3238
rect 36822 3216 37386 3236
rect 37476 3126 37504 5578
rect 38028 5574 38056 8092
rect 39132 5642 39160 8092
rect 40052 8078 40342 8106
rect 40052 5658 40080 8078
rect 41432 5658 41460 8092
rect 39120 5636 39172 5642
rect 39120 5578 39172 5584
rect 39960 5630 40080 5658
rect 41340 5630 41460 5658
rect 38016 5568 38068 5574
rect 38016 5510 38068 5516
rect 39960 3534 39988 5630
rect 40960 4072 41012 4078
rect 40960 4014 41012 4020
rect 39948 3528 40000 3534
rect 39948 3470 40000 3476
rect 38568 3460 38620 3466
rect 38568 3402 38620 3408
rect 37464 3120 37516 3126
rect 37464 3062 37516 3068
rect 37464 2984 37516 2990
rect 37464 2926 37516 2932
rect 36822 2204 37386 2224
rect 36822 2202 36836 2204
rect 36892 2202 36916 2204
rect 36972 2202 36996 2204
rect 37052 2202 37076 2204
rect 37132 2202 37156 2204
rect 37212 2202 37236 2204
rect 37292 2202 37316 2204
rect 37372 2202 37386 2204
rect 37066 2150 37076 2202
rect 37132 2150 37142 2202
rect 36822 2148 36836 2150
rect 36892 2148 36916 2150
rect 36972 2148 36996 2150
rect 37052 2148 37076 2150
rect 37132 2148 37156 2150
rect 37212 2148 37236 2150
rect 37292 2148 37316 2150
rect 37372 2148 37386 2150
rect 36822 2128 37386 2148
rect 37476 1986 37504 2926
rect 37384 1958 37504 1986
rect 37384 480 37412 1958
rect 38580 480 38608 3402
rect 39764 2848 39816 2854
rect 39764 2790 39816 2796
rect 39776 480 39804 2790
rect 40972 480 41000 4014
rect 41340 3602 41368 5630
rect 42156 4140 42208 4146
rect 42156 4082 42208 4088
rect 41328 3596 41380 3602
rect 41328 3538 41380 3544
rect 42168 480 42196 4082
rect 42536 3398 42564 8092
rect 42800 5568 42852 5574
rect 42800 5510 42852 5516
rect 42812 3466 42840 5510
rect 43352 3936 43404 3942
rect 43352 3878 43404 3884
rect 42800 3460 42852 3466
rect 42800 3402 42852 3408
rect 42524 3392 42576 3398
rect 42524 3334 42576 3340
rect 43364 480 43392 3878
rect 43732 2990 43760 8092
rect 44836 5574 44864 8092
rect 45572 8078 45954 8106
rect 46952 8078 47058 8106
rect 45572 5658 45600 8078
rect 45480 5630 45600 5658
rect 44824 5568 44876 5574
rect 44824 5510 44876 5516
rect 44548 3596 44600 3602
rect 44548 3538 44600 3544
rect 43720 2984 43772 2990
rect 43720 2926 43772 2932
rect 44560 480 44588 3538
rect 45480 2854 45508 5630
rect 46952 5556 46980 8078
rect 46860 5528 46980 5556
rect 46860 4078 46888 5528
rect 48240 4146 48268 8092
rect 48228 4140 48280 4146
rect 48228 4082 48280 4088
rect 46848 4072 46900 4078
rect 46848 4014 46900 4020
rect 49344 3942 49372 8092
rect 49332 3936 49384 3942
rect 49332 3878 49384 3884
rect 45744 3664 45796 3670
rect 45744 3606 45796 3612
rect 45468 2848 45520 2854
rect 45468 2790 45520 2796
rect 45756 480 45784 3606
rect 50448 3602 50476 8092
rect 50528 4072 50580 4078
rect 50528 4014 50580 4020
rect 50436 3596 50488 3602
rect 50436 3538 50488 3544
rect 48136 3460 48188 3466
rect 48136 3402 48188 3408
rect 46940 3120 46992 3126
rect 46940 3062 46992 3068
rect 46952 480 46980 3062
rect 48148 480 48176 3402
rect 49332 3188 49384 3194
rect 49332 3130 49384 3136
rect 49344 480 49372 3130
rect 50540 480 50568 4014
rect 51644 3670 51672 8092
rect 51632 3664 51684 3670
rect 51632 3606 51684 3612
rect 51632 3528 51684 3534
rect 51632 3470 51684 3476
rect 51644 480 51672 3470
rect 52748 3126 52776 8092
rect 53852 5556 53880 8092
rect 53668 5528 53880 5556
rect 54680 8078 55062 8106
rect 52828 3596 52880 3602
rect 52828 3538 52880 3544
rect 52736 3120 52788 3126
rect 52736 3062 52788 3068
rect 52840 480 52868 3538
rect 53668 3466 53696 5528
rect 53656 3460 53708 3466
rect 53656 3402 53708 3408
rect 54024 3460 54076 3466
rect 54024 3402 54076 3408
rect 54036 480 54064 3402
rect 54680 3194 54708 8078
rect 54822 6012 55386 6032
rect 54822 6010 54836 6012
rect 54892 6010 54916 6012
rect 54972 6010 54996 6012
rect 55052 6010 55076 6012
rect 55132 6010 55156 6012
rect 55212 6010 55236 6012
rect 55292 6010 55316 6012
rect 55372 6010 55386 6012
rect 55066 5958 55076 6010
rect 55132 5958 55142 6010
rect 54822 5956 54836 5958
rect 54892 5956 54916 5958
rect 54972 5956 54996 5958
rect 55052 5956 55076 5958
rect 55132 5956 55156 5958
rect 55212 5956 55236 5958
rect 55292 5956 55316 5958
rect 55372 5956 55386 5958
rect 54822 5936 55386 5956
rect 55404 5568 55456 5574
rect 55404 5510 55456 5516
rect 54822 4924 55386 4944
rect 54822 4922 54836 4924
rect 54892 4922 54916 4924
rect 54972 4922 54996 4924
rect 55052 4922 55076 4924
rect 55132 4922 55156 4924
rect 55212 4922 55236 4924
rect 55292 4922 55316 4924
rect 55372 4922 55386 4924
rect 55066 4870 55076 4922
rect 55132 4870 55142 4922
rect 54822 4868 54836 4870
rect 54892 4868 54916 4870
rect 54972 4868 54996 4870
rect 55052 4868 55076 4870
rect 55132 4868 55156 4870
rect 55212 4868 55236 4870
rect 55292 4868 55316 4870
rect 55372 4868 55386 4870
rect 54822 4848 55386 4868
rect 54822 3836 55386 3856
rect 54822 3834 54836 3836
rect 54892 3834 54916 3836
rect 54972 3834 54996 3836
rect 55052 3834 55076 3836
rect 55132 3834 55156 3836
rect 55212 3834 55236 3836
rect 55292 3834 55316 3836
rect 55372 3834 55386 3836
rect 55066 3782 55076 3834
rect 55132 3782 55142 3834
rect 54822 3780 54836 3782
rect 54892 3780 54916 3782
rect 54972 3780 54996 3782
rect 55052 3780 55076 3782
rect 55132 3780 55156 3782
rect 55212 3780 55236 3782
rect 55292 3780 55316 3782
rect 55372 3780 55386 3782
rect 54822 3760 55386 3780
rect 54668 3188 54720 3194
rect 54668 3130 54720 3136
rect 54822 2748 55386 2768
rect 54822 2746 54836 2748
rect 54892 2746 54916 2748
rect 54972 2746 54996 2748
rect 55052 2746 55076 2748
rect 55132 2746 55156 2748
rect 55212 2746 55236 2748
rect 55292 2746 55316 2748
rect 55372 2746 55386 2748
rect 55066 2694 55076 2746
rect 55132 2694 55142 2746
rect 54822 2692 54836 2694
rect 54892 2692 54916 2694
rect 54972 2692 54996 2694
rect 55052 2692 55076 2694
rect 55132 2692 55156 2694
rect 55212 2692 55236 2694
rect 55292 2692 55316 2694
rect 55372 2692 55386 2694
rect 54822 2672 55386 2692
rect 55416 2530 55444 5510
rect 56152 4078 56180 8092
rect 56140 4072 56192 4078
rect 56140 4014 56192 4020
rect 57256 3534 57284 8092
rect 58452 3602 58480 8092
rect 58440 3596 58492 3602
rect 58440 3538 58492 3544
rect 57244 3528 57296 3534
rect 57244 3470 57296 3476
rect 57612 3528 57664 3534
rect 57612 3470 57664 3476
rect 56416 3188 56468 3194
rect 56416 3130 56468 3136
rect 55232 2502 55444 2530
rect 55232 480 55260 2502
rect 56428 480 56456 3130
rect 57624 480 57652 3470
rect 59556 3466 59584 8092
rect 60660 5574 60688 8092
rect 60648 5568 60700 5574
rect 60648 5510 60700 5516
rect 61200 4140 61252 4146
rect 61200 4082 61252 4088
rect 60004 4004 60056 4010
rect 60004 3946 60056 3952
rect 59544 3460 59596 3466
rect 59544 3402 59596 3408
rect 58808 3392 58860 3398
rect 58808 3334 58860 3340
rect 58820 480 58848 3334
rect 60016 480 60044 3946
rect 61212 480 61240 4082
rect 61856 3194 61884 8092
rect 62396 5568 62448 5574
rect 62396 5510 62448 5516
rect 61844 3188 61896 3194
rect 61844 3130 61896 3136
rect 62408 480 62436 5510
rect 62960 3534 62988 8092
rect 63592 6180 63644 6186
rect 63592 6122 63644 6128
rect 62948 3528 63000 3534
rect 62948 3470 63000 3476
rect 63604 480 63632 6122
rect 64064 3398 64092 8092
rect 65260 4010 65288 8092
rect 66364 4146 66392 8092
rect 67468 5574 67496 8092
rect 68664 6186 68692 8092
rect 68652 6180 68704 6186
rect 68652 6122 68704 6128
rect 69480 5636 69532 5642
rect 69480 5578 69532 5584
rect 67456 5568 67508 5574
rect 67456 5510 67508 5516
rect 66352 4140 66404 4146
rect 66352 4082 66404 4088
rect 65248 4004 65300 4010
rect 65248 3946 65300 3952
rect 64788 3664 64840 3670
rect 64788 3606 64840 3612
rect 64052 3392 64104 3398
rect 64052 3334 64104 3340
rect 64800 480 64828 3606
rect 65984 3528 66036 3534
rect 65984 3470 66036 3476
rect 65996 480 66024 3470
rect 68284 3460 68336 3466
rect 68284 3402 68336 3408
rect 67180 3188 67232 3194
rect 67180 3130 67232 3136
rect 67192 480 67220 3130
rect 68296 480 68324 3402
rect 69492 480 69520 5578
rect 69768 3670 69796 8092
rect 70676 6520 70728 6526
rect 70676 6462 70728 6468
rect 69756 3664 69808 3670
rect 69756 3606 69808 3612
rect 70688 480 70716 6462
rect 70872 3534 70900 8092
rect 71872 5568 71924 5574
rect 71872 5510 71924 5516
rect 70860 3528 70912 3534
rect 70860 3470 70912 3476
rect 71884 480 71912 5510
rect 72068 3194 72096 8092
rect 73186 8078 73476 8106
rect 72822 5468 73386 5488
rect 72822 5466 72836 5468
rect 72892 5466 72916 5468
rect 72972 5466 72996 5468
rect 73052 5466 73076 5468
rect 73132 5466 73156 5468
rect 73212 5466 73236 5468
rect 73292 5466 73316 5468
rect 73372 5466 73386 5468
rect 73066 5414 73076 5466
rect 73132 5414 73142 5466
rect 72822 5412 72836 5414
rect 72892 5412 72916 5414
rect 72972 5412 72996 5414
rect 73052 5412 73076 5414
rect 73132 5412 73156 5414
rect 73212 5412 73236 5414
rect 73292 5412 73316 5414
rect 73372 5412 73386 5414
rect 72822 5392 73386 5412
rect 72822 4380 73386 4400
rect 72822 4378 72836 4380
rect 72892 4378 72916 4380
rect 72972 4378 72996 4380
rect 73052 4378 73076 4380
rect 73132 4378 73156 4380
rect 73212 4378 73236 4380
rect 73292 4378 73316 4380
rect 73372 4378 73386 4380
rect 73066 4326 73076 4378
rect 73132 4326 73142 4378
rect 72822 4324 72836 4326
rect 72892 4324 72916 4326
rect 72972 4324 72996 4326
rect 73052 4324 73076 4326
rect 73132 4324 73156 4326
rect 73212 4324 73236 4326
rect 73292 4324 73316 4326
rect 73372 4324 73386 4326
rect 72822 4304 73386 4324
rect 72700 3528 72752 3534
rect 72700 3470 72752 3476
rect 72056 3188 72108 3194
rect 72056 3130 72108 3136
rect 72712 1850 72740 3470
rect 73448 3466 73476 8078
rect 74276 5642 74304 8092
rect 75472 6526 75500 8092
rect 75460 6520 75512 6526
rect 75460 6462 75512 6468
rect 75460 5704 75512 5710
rect 75460 5646 75512 5652
rect 74264 5636 74316 5642
rect 74264 5578 74316 5584
rect 74264 3596 74316 3602
rect 74264 3538 74316 3544
rect 73436 3460 73488 3466
rect 73436 3402 73488 3408
rect 72822 3292 73386 3312
rect 72822 3290 72836 3292
rect 72892 3290 72916 3292
rect 72972 3290 72996 3292
rect 73052 3290 73076 3292
rect 73132 3290 73156 3292
rect 73212 3290 73236 3292
rect 73292 3290 73316 3292
rect 73372 3290 73386 3292
rect 73066 3238 73076 3290
rect 73132 3238 73142 3290
rect 72822 3236 72836 3238
rect 72892 3236 72916 3238
rect 72972 3236 72996 3238
rect 73052 3236 73076 3238
rect 73132 3236 73156 3238
rect 73212 3236 73236 3238
rect 73292 3236 73316 3238
rect 73372 3236 73386 3238
rect 72822 3216 73386 3236
rect 72822 2204 73386 2224
rect 72822 2202 72836 2204
rect 72892 2202 72916 2204
rect 72972 2202 72996 2204
rect 73052 2202 73076 2204
rect 73132 2202 73156 2204
rect 73212 2202 73236 2204
rect 73292 2202 73316 2204
rect 73372 2202 73386 2204
rect 73066 2150 73076 2202
rect 73132 2150 73142 2202
rect 72822 2148 72836 2150
rect 72892 2148 72916 2150
rect 72972 2148 72996 2150
rect 73052 2148 73076 2150
rect 73132 2148 73156 2150
rect 73212 2148 73236 2150
rect 73292 2148 73316 2150
rect 73372 2148 73386 2150
rect 72822 2128 73386 2148
rect 72712 1822 73108 1850
rect 73080 480 73108 1822
rect 74276 480 74304 3538
rect 75472 480 75500 5646
rect 76576 5574 76604 8092
rect 76564 5568 76616 5574
rect 76564 5510 76616 5516
rect 76656 5568 76708 5574
rect 76656 5510 76708 5516
rect 76668 480 76696 5510
rect 77680 3534 77708 8092
rect 77852 5636 77904 5642
rect 77852 5578 77904 5584
rect 77668 3528 77720 3534
rect 77668 3470 77720 3476
rect 77864 480 77892 5578
rect 78876 3602 78904 8092
rect 79048 5772 79100 5778
rect 79048 5714 79100 5720
rect 78864 3596 78916 3602
rect 78864 3538 78916 3544
rect 79060 480 79088 5714
rect 79980 5710 80008 8092
rect 79968 5704 80020 5710
rect 79968 5646 80020 5652
rect 80244 5704 80296 5710
rect 80244 5646 80296 5652
rect 80256 480 80284 5646
rect 81084 5574 81112 8092
rect 82280 5642 82308 8092
rect 83384 5778 83412 8092
rect 83832 6248 83884 6254
rect 83832 6190 83884 6196
rect 83372 5772 83424 5778
rect 83372 5714 83424 5720
rect 82268 5636 82320 5642
rect 82268 5578 82320 5584
rect 82636 5636 82688 5642
rect 82636 5578 82688 5584
rect 81072 5568 81124 5574
rect 81072 5510 81124 5516
rect 81440 5568 81492 5574
rect 81440 5510 81492 5516
rect 81452 480 81480 5510
rect 82648 480 82676 5578
rect 83844 480 83872 6190
rect 84488 5710 84516 8092
rect 84936 5772 84988 5778
rect 84936 5714 84988 5720
rect 84476 5704 84528 5710
rect 84476 5646 84528 5652
rect 84948 480 84976 5714
rect 85592 5574 85620 8092
rect 86788 5642 86816 8092
rect 87892 6254 87920 8092
rect 87880 6248 87932 6254
rect 87880 6190 87932 6196
rect 87328 6180 87380 6186
rect 87328 6122 87380 6128
rect 86776 5636 86828 5642
rect 86776 5578 86828 5584
rect 85580 5568 85632 5574
rect 85580 5510 85632 5516
rect 86132 5568 86184 5574
rect 86132 5510 86184 5516
rect 86144 480 86172 5510
rect 87340 480 87368 6122
rect 88996 5778 89024 8092
rect 88984 5772 89036 5778
rect 88984 5714 89036 5720
rect 89720 5772 89772 5778
rect 89720 5714 89772 5720
rect 88524 5704 88576 5710
rect 88524 5646 88576 5652
rect 88536 480 88564 5646
rect 89732 480 89760 5714
rect 90192 5574 90220 8092
rect 91296 6186 91324 8092
rect 91284 6180 91336 6186
rect 91284 6122 91336 6128
rect 90822 6012 91386 6032
rect 90822 6010 90836 6012
rect 90892 6010 90916 6012
rect 90972 6010 90996 6012
rect 91052 6010 91076 6012
rect 91132 6010 91156 6012
rect 91212 6010 91236 6012
rect 91292 6010 91316 6012
rect 91372 6010 91386 6012
rect 91066 5958 91076 6010
rect 91132 5958 91142 6010
rect 90822 5956 90836 5958
rect 90892 5956 90916 5958
rect 90972 5956 90996 5958
rect 91052 5956 91076 5958
rect 91132 5956 91156 5958
rect 91212 5956 91236 5958
rect 91292 5956 91316 5958
rect 91372 5956 91386 5958
rect 90822 5936 91386 5956
rect 92400 5710 92428 8092
rect 93308 6384 93360 6390
rect 93308 6326 93360 6332
rect 92388 5704 92440 5710
rect 92388 5646 92440 5652
rect 90732 5636 90784 5642
rect 90732 5578 90784 5584
rect 90180 5568 90232 5574
rect 90180 5510 90232 5516
rect 90744 2530 90772 5578
rect 92112 5568 92164 5574
rect 92112 5510 92164 5516
rect 90822 4924 91386 4944
rect 90822 4922 90836 4924
rect 90892 4922 90916 4924
rect 90972 4922 90996 4924
rect 91052 4922 91076 4924
rect 91132 4922 91156 4924
rect 91212 4922 91236 4924
rect 91292 4922 91316 4924
rect 91372 4922 91386 4924
rect 91066 4870 91076 4922
rect 91132 4870 91142 4922
rect 90822 4868 90836 4870
rect 90892 4868 90916 4870
rect 90972 4868 90996 4870
rect 91052 4868 91076 4870
rect 91132 4868 91156 4870
rect 91212 4868 91236 4870
rect 91292 4868 91316 4870
rect 91372 4868 91386 4870
rect 90822 4848 91386 4868
rect 90822 3836 91386 3856
rect 90822 3834 90836 3836
rect 90892 3834 90916 3836
rect 90972 3834 90996 3836
rect 91052 3834 91076 3836
rect 91132 3834 91156 3836
rect 91212 3834 91236 3836
rect 91292 3834 91316 3836
rect 91372 3834 91386 3836
rect 91066 3782 91076 3834
rect 91132 3782 91142 3834
rect 90822 3780 90836 3782
rect 90892 3780 90916 3782
rect 90972 3780 90996 3782
rect 91052 3780 91076 3782
rect 91132 3780 91156 3782
rect 91212 3780 91236 3782
rect 91292 3780 91316 3782
rect 91372 3780 91386 3782
rect 90822 3760 91386 3780
rect 90822 2748 91386 2768
rect 90822 2746 90836 2748
rect 90892 2746 90916 2748
rect 90972 2746 90996 2748
rect 91052 2746 91076 2748
rect 91132 2746 91156 2748
rect 91212 2746 91236 2748
rect 91292 2746 91316 2748
rect 91372 2746 91386 2748
rect 91066 2694 91076 2746
rect 91132 2694 91142 2746
rect 90822 2692 90836 2694
rect 90892 2692 90916 2694
rect 90972 2692 90996 2694
rect 91052 2692 91076 2694
rect 91132 2692 91156 2694
rect 91212 2692 91236 2694
rect 91292 2692 91316 2694
rect 91372 2692 91386 2694
rect 90822 2672 91386 2692
rect 90744 2502 90956 2530
rect 90928 480 90956 2502
rect 92124 480 92152 5510
rect 93320 480 93348 6326
rect 93596 5778 93624 8092
rect 94504 5840 94556 5846
rect 94504 5782 94556 5788
rect 93584 5772 93636 5778
rect 93584 5714 93636 5720
rect 94516 480 94544 5782
rect 94700 5642 94728 8092
rect 95700 5704 95752 5710
rect 95700 5646 95752 5652
rect 94688 5636 94740 5642
rect 94688 5578 94740 5584
rect 95712 480 95740 5646
rect 95804 5574 95832 8092
rect 97000 6390 97028 8092
rect 96988 6384 97040 6390
rect 96988 6326 97040 6332
rect 98104 5846 98132 8092
rect 98092 5840 98144 5846
rect 98092 5782 98144 5788
rect 96896 5772 96948 5778
rect 96896 5714 96948 5720
rect 95792 5568 95844 5574
rect 95792 5510 95844 5516
rect 96908 480 96936 5714
rect 99208 5710 99236 8092
rect 100404 5778 100432 8092
rect 100392 5772 100444 5778
rect 100392 5714 100444 5720
rect 99196 5704 99248 5710
rect 99196 5646 99248 5652
rect 100484 5704 100536 5710
rect 100484 5646 100536 5652
rect 98092 5636 98144 5642
rect 98092 5578 98144 5584
rect 98104 480 98132 5578
rect 99288 5568 99340 5574
rect 99288 5510 99340 5516
rect 99300 480 99328 5510
rect 100496 480 100524 5646
rect 101508 5642 101536 8092
rect 101496 5636 101548 5642
rect 101496 5578 101548 5584
rect 101588 5636 101640 5642
rect 101588 5578 101640 5584
rect 101600 480 101628 5578
rect 102612 5574 102640 8092
rect 103808 5710 103836 8092
rect 103796 5704 103848 5710
rect 103796 5646 103848 5652
rect 103980 5704 104032 5710
rect 103980 5646 104032 5652
rect 102600 5568 102652 5574
rect 102600 5510 102652 5516
rect 102784 5568 102836 5574
rect 102784 5510 102836 5516
rect 102796 480 102824 5510
rect 103992 480 104020 5646
rect 104912 5642 104940 8092
rect 105176 5772 105228 5778
rect 105176 5714 105228 5720
rect 104900 5636 104952 5642
rect 104900 5578 104952 5584
rect 105188 480 105216 5714
rect 106016 5574 106044 8092
rect 107212 5710 107240 8092
rect 108316 5778 108344 8092
rect 108304 5772 108356 5778
rect 108304 5714 108356 5720
rect 107200 5704 107252 5710
rect 107200 5646 107252 5652
rect 107568 5704 107620 5710
rect 107568 5646 107620 5652
rect 106372 5636 106424 5642
rect 106372 5578 106424 5584
rect 106004 5568 106056 5574
rect 106004 5510 106056 5516
rect 106384 480 106412 5578
rect 107580 480 107608 5646
rect 109420 5642 109448 8092
rect 110616 5710 110644 8092
rect 110604 5704 110656 5710
rect 110604 5646 110656 5652
rect 111156 5704 111208 5710
rect 111156 5646 111208 5652
rect 109408 5636 109460 5642
rect 109408 5578 109460 5584
rect 109960 5636 110012 5642
rect 109960 5578 110012 5584
rect 108672 5568 108724 5574
rect 108672 5510 108724 5516
rect 108684 1986 108712 5510
rect 108822 5468 109386 5488
rect 108822 5466 108836 5468
rect 108892 5466 108916 5468
rect 108972 5466 108996 5468
rect 109052 5466 109076 5468
rect 109132 5466 109156 5468
rect 109212 5466 109236 5468
rect 109292 5466 109316 5468
rect 109372 5466 109386 5468
rect 109066 5414 109076 5466
rect 109132 5414 109142 5466
rect 108822 5412 108836 5414
rect 108892 5412 108916 5414
rect 108972 5412 108996 5414
rect 109052 5412 109076 5414
rect 109132 5412 109156 5414
rect 109212 5412 109236 5414
rect 109292 5412 109316 5414
rect 109372 5412 109386 5414
rect 108822 5392 109386 5412
rect 108822 4380 109386 4400
rect 108822 4378 108836 4380
rect 108892 4378 108916 4380
rect 108972 4378 108996 4380
rect 109052 4378 109076 4380
rect 109132 4378 109156 4380
rect 109212 4378 109236 4380
rect 109292 4378 109316 4380
rect 109372 4378 109386 4380
rect 109066 4326 109076 4378
rect 109132 4326 109142 4378
rect 108822 4324 108836 4326
rect 108892 4324 108916 4326
rect 108972 4324 108996 4326
rect 109052 4324 109076 4326
rect 109132 4324 109156 4326
rect 109212 4324 109236 4326
rect 109292 4324 109316 4326
rect 109372 4324 109386 4326
rect 108822 4304 109386 4324
rect 108822 3292 109386 3312
rect 108822 3290 108836 3292
rect 108892 3290 108916 3292
rect 108972 3290 108996 3292
rect 109052 3290 109076 3292
rect 109132 3290 109156 3292
rect 109212 3290 109236 3292
rect 109292 3290 109316 3292
rect 109372 3290 109386 3292
rect 109066 3238 109076 3290
rect 109132 3238 109142 3290
rect 108822 3236 108836 3238
rect 108892 3236 108916 3238
rect 108972 3236 108996 3238
rect 109052 3236 109076 3238
rect 109132 3236 109156 3238
rect 109212 3236 109236 3238
rect 109292 3236 109316 3238
rect 109372 3236 109386 3238
rect 108822 3216 109386 3236
rect 108822 2204 109386 2224
rect 108822 2202 108836 2204
rect 108892 2202 108916 2204
rect 108972 2202 108996 2204
rect 109052 2202 109076 2204
rect 109132 2202 109156 2204
rect 109212 2202 109236 2204
rect 109292 2202 109316 2204
rect 109372 2202 109386 2204
rect 109066 2150 109076 2202
rect 109132 2150 109142 2202
rect 108822 2148 108836 2150
rect 108892 2148 108916 2150
rect 108972 2148 108996 2150
rect 109052 2148 109076 2150
rect 109132 2148 109156 2150
rect 109212 2148 109236 2150
rect 109292 2148 109316 2150
rect 109372 2148 109386 2150
rect 108822 2128 109386 2148
rect 108684 1958 108804 1986
rect 108776 480 108804 1958
rect 109972 480 110000 5578
rect 111168 480 111196 5646
rect 111720 5574 111748 8092
rect 112824 5642 112852 8092
rect 114020 5710 114048 8092
rect 114008 5704 114060 5710
rect 114008 5646 114060 5652
rect 114744 5704 114796 5710
rect 114744 5646 114796 5652
rect 112812 5636 112864 5642
rect 112812 5578 112864 5584
rect 113548 5636 113600 5642
rect 113548 5578 113600 5584
rect 111708 5568 111760 5574
rect 111708 5510 111760 5516
rect 112352 5568 112404 5574
rect 112352 5510 112404 5516
rect 112364 480 112392 5510
rect 113560 480 113588 5578
rect 114756 480 114784 5646
rect 115124 5574 115152 8092
rect 116228 5642 116256 8092
rect 117424 5710 117452 8092
rect 118240 5772 118292 5778
rect 118240 5714 118292 5720
rect 117412 5704 117464 5710
rect 117412 5646 117464 5652
rect 116216 5636 116268 5642
rect 116216 5578 116268 5584
rect 117136 5636 117188 5642
rect 117136 5578 117188 5584
rect 115112 5568 115164 5574
rect 115112 5510 115164 5516
rect 115940 5568 115992 5574
rect 115940 5510 115992 5516
rect 115952 480 115980 5510
rect 117148 480 117176 5578
rect 118252 480 118280 5714
rect 118528 5574 118556 8092
rect 119632 5642 119660 8092
rect 120828 5778 120856 8092
rect 120816 5772 120868 5778
rect 120816 5714 120868 5720
rect 120632 5704 120684 5710
rect 120632 5646 120684 5652
rect 119620 5636 119672 5642
rect 119620 5578 119672 5584
rect 118516 5568 118568 5574
rect 118516 5510 118568 5516
rect 119436 5568 119488 5574
rect 119436 5510 119488 5516
rect 119448 480 119476 5510
rect 120644 480 120672 5646
rect 121828 5636 121880 5642
rect 121828 5578 121880 5584
rect 121840 480 121868 5578
rect 121932 5574 121960 8092
rect 123036 5710 123064 8092
rect 123024 5704 123076 5710
rect 123024 5646 123076 5652
rect 124140 5642 124168 8092
rect 124128 5636 124180 5642
rect 124128 5578 124180 5584
rect 124220 5636 124272 5642
rect 124220 5578 124272 5584
rect 121920 5568 121972 5574
rect 121920 5510 121972 5516
rect 123024 5568 123076 5574
rect 123024 5510 123076 5516
rect 123036 480 123064 5510
rect 124232 480 124260 5578
rect 125336 5574 125364 8092
rect 126440 5642 126468 8092
rect 126822 6012 127386 6032
rect 126822 6010 126836 6012
rect 126892 6010 126916 6012
rect 126972 6010 126996 6012
rect 127052 6010 127076 6012
rect 127132 6010 127156 6012
rect 127212 6010 127236 6012
rect 127292 6010 127316 6012
rect 127372 6010 127386 6012
rect 127066 5958 127076 6010
rect 127132 5958 127142 6010
rect 126822 5956 126836 5958
rect 126892 5956 126916 5958
rect 126972 5956 126996 5958
rect 127052 5956 127076 5958
rect 127132 5956 127156 5958
rect 127212 5956 127236 5958
rect 127292 5956 127316 5958
rect 127372 5956 127386 5958
rect 126822 5936 127386 5956
rect 126428 5636 126480 5642
rect 126428 5578 126480 5584
rect 126612 5636 126664 5642
rect 126612 5578 126664 5584
rect 125324 5568 125376 5574
rect 125324 5510 125376 5516
rect 125416 5568 125468 5574
rect 125416 5510 125468 5516
rect 125428 480 125456 5510
rect 126624 480 126652 5578
rect 127544 5574 127572 8092
rect 128740 5642 128768 8092
rect 128728 5636 128780 5642
rect 128728 5578 128780 5584
rect 129004 5636 129056 5642
rect 129004 5578 129056 5584
rect 127532 5568 127584 5574
rect 127532 5510 127584 5516
rect 127808 5568 127860 5574
rect 127808 5510 127860 5516
rect 126822 4924 127386 4944
rect 126822 4922 126836 4924
rect 126892 4922 126916 4924
rect 126972 4922 126996 4924
rect 127052 4922 127076 4924
rect 127132 4922 127156 4924
rect 127212 4922 127236 4924
rect 127292 4922 127316 4924
rect 127372 4922 127386 4924
rect 127066 4870 127076 4922
rect 127132 4870 127142 4922
rect 126822 4868 126836 4870
rect 126892 4868 126916 4870
rect 126972 4868 126996 4870
rect 127052 4868 127076 4870
rect 127132 4868 127156 4870
rect 127212 4868 127236 4870
rect 127292 4868 127316 4870
rect 127372 4868 127386 4870
rect 126822 4848 127386 4868
rect 126822 3836 127386 3856
rect 126822 3834 126836 3836
rect 126892 3834 126916 3836
rect 126972 3834 126996 3836
rect 127052 3834 127076 3836
rect 127132 3834 127156 3836
rect 127212 3834 127236 3836
rect 127292 3834 127316 3836
rect 127372 3834 127386 3836
rect 127066 3782 127076 3834
rect 127132 3782 127142 3834
rect 126822 3780 126836 3782
rect 126892 3780 126916 3782
rect 126972 3780 126996 3782
rect 127052 3780 127076 3782
rect 127132 3780 127156 3782
rect 127212 3780 127236 3782
rect 127292 3780 127316 3782
rect 127372 3780 127386 3782
rect 126822 3760 127386 3780
rect 126822 2748 127386 2768
rect 126822 2746 126836 2748
rect 126892 2746 126916 2748
rect 126972 2746 126996 2748
rect 127052 2746 127076 2748
rect 127132 2746 127156 2748
rect 127212 2746 127236 2748
rect 127292 2746 127316 2748
rect 127372 2746 127386 2748
rect 127066 2694 127076 2746
rect 127132 2694 127142 2746
rect 126822 2692 126836 2694
rect 126892 2692 126916 2694
rect 126972 2692 126996 2694
rect 127052 2692 127076 2694
rect 127132 2692 127156 2694
rect 127212 2692 127236 2694
rect 127292 2692 127316 2694
rect 127372 2692 127386 2694
rect 126822 2672 127386 2692
rect 127820 480 127848 5510
rect 129016 480 129044 5578
rect 129844 5574 129872 8092
rect 130948 5642 130976 8092
rect 130936 5636 130988 5642
rect 130936 5578 130988 5584
rect 131396 5636 131448 5642
rect 131396 5578 131448 5584
rect 129832 5568 129884 5574
rect 129832 5510 129884 5516
rect 130200 5568 130252 5574
rect 130200 5510 130252 5516
rect 130212 480 130240 5510
rect 131408 480 131436 5578
rect 132144 5574 132172 8092
rect 132592 5704 132644 5710
rect 132592 5646 132644 5652
rect 132132 5568 132184 5574
rect 132132 5510 132184 5516
rect 132604 480 132632 5646
rect 133248 5642 133276 8092
rect 134352 5710 134380 8092
rect 134340 5704 134392 5710
rect 134340 5646 134392 5652
rect 133236 5636 133288 5642
rect 133236 5578 133288 5584
rect 134892 5636 134944 5642
rect 134892 5578 134944 5584
rect 133788 5568 133840 5574
rect 133788 5510 133840 5516
rect 133800 480 133828 5510
rect 134904 480 134932 5578
rect 135548 5574 135576 8092
rect 136652 5642 136680 8092
rect 136640 5636 136692 5642
rect 136640 5578 136692 5584
rect 137284 5636 137336 5642
rect 137284 5578 137336 5584
rect 135536 5568 135588 5574
rect 135536 5510 135588 5516
rect 136088 5568 136140 5574
rect 136088 5510 136140 5516
rect 136100 480 136128 5510
rect 137296 480 137324 5578
rect 137756 5574 137784 8092
rect 138952 5642 138980 8092
rect 138940 5636 138992 5642
rect 138940 5578 138992 5584
rect 139676 5636 139728 5642
rect 139676 5578 139728 5584
rect 137744 5568 137796 5574
rect 137744 5510 137796 5516
rect 138480 5568 138532 5574
rect 138480 5510 138532 5516
rect 138492 480 138520 5510
rect 139688 480 139716 5578
rect 140056 5574 140084 8092
rect 141160 5642 141188 8092
rect 141148 5636 141200 5642
rect 141148 5578 141200 5584
rect 142068 5636 142120 5642
rect 142068 5578 142120 5584
rect 140044 5568 140096 5574
rect 140044 5510 140096 5516
rect 140872 5568 140924 5574
rect 140872 5510 140924 5516
rect 140884 480 140912 5510
rect 142080 480 142108 5578
rect 142356 5574 142384 8092
rect 143264 5704 143316 5710
rect 143264 5646 143316 5652
rect 142344 5568 142396 5574
rect 142344 5510 142396 5516
rect 143276 480 143304 5646
rect 143460 5642 143488 8092
rect 144564 5710 144592 8092
rect 144552 5704 144604 5710
rect 144552 5646 144604 5652
rect 145656 5704 145708 5710
rect 145656 5646 145708 5652
rect 143448 5636 143500 5642
rect 143448 5578 143500 5584
rect 144460 5568 144512 5574
rect 144460 5510 144512 5516
rect 144472 480 144500 5510
rect 144822 5468 145386 5488
rect 144822 5466 144836 5468
rect 144892 5466 144916 5468
rect 144972 5466 144996 5468
rect 145052 5466 145076 5468
rect 145132 5466 145156 5468
rect 145212 5466 145236 5468
rect 145292 5466 145316 5468
rect 145372 5466 145386 5468
rect 145066 5414 145076 5466
rect 145132 5414 145142 5466
rect 144822 5412 144836 5414
rect 144892 5412 144916 5414
rect 144972 5412 144996 5414
rect 145052 5412 145076 5414
rect 145132 5412 145156 5414
rect 145212 5412 145236 5414
rect 145292 5412 145316 5414
rect 145372 5412 145386 5414
rect 144822 5392 145386 5412
rect 144822 4380 145386 4400
rect 144822 4378 144836 4380
rect 144892 4378 144916 4380
rect 144972 4378 144996 4380
rect 145052 4378 145076 4380
rect 145132 4378 145156 4380
rect 145212 4378 145236 4380
rect 145292 4378 145316 4380
rect 145372 4378 145386 4380
rect 145066 4326 145076 4378
rect 145132 4326 145142 4378
rect 144822 4324 144836 4326
rect 144892 4324 144916 4326
rect 144972 4324 144996 4326
rect 145052 4324 145076 4326
rect 145132 4324 145156 4326
rect 145212 4324 145236 4326
rect 145292 4324 145316 4326
rect 145372 4324 145386 4326
rect 144822 4304 145386 4324
rect 144822 3292 145386 3312
rect 144822 3290 144836 3292
rect 144892 3290 144916 3292
rect 144972 3290 144996 3292
rect 145052 3290 145076 3292
rect 145132 3290 145156 3292
rect 145212 3290 145236 3292
rect 145292 3290 145316 3292
rect 145372 3290 145386 3292
rect 145066 3238 145076 3290
rect 145132 3238 145142 3290
rect 144822 3236 144836 3238
rect 144892 3236 144916 3238
rect 144972 3236 144996 3238
rect 145052 3236 145076 3238
rect 145132 3236 145156 3238
rect 145212 3236 145236 3238
rect 145292 3236 145316 3238
rect 145372 3236 145386 3238
rect 144822 3216 145386 3236
rect 144822 2204 145386 2224
rect 144822 2202 144836 2204
rect 144892 2202 144916 2204
rect 144972 2202 144996 2204
rect 145052 2202 145076 2204
rect 145132 2202 145156 2204
rect 145212 2202 145236 2204
rect 145292 2202 145316 2204
rect 145372 2202 145386 2204
rect 145066 2150 145076 2202
rect 145132 2150 145142 2202
rect 144822 2148 144836 2150
rect 144892 2148 144916 2150
rect 144972 2148 144996 2150
rect 145052 2148 145076 2150
rect 145132 2148 145156 2150
rect 145212 2148 145236 2150
rect 145292 2148 145316 2150
rect 145372 2148 145386 2150
rect 144822 2128 145386 2148
rect 145668 480 145696 5646
rect 145760 5574 145788 8092
rect 146864 5710 146892 8092
rect 146852 5704 146904 5710
rect 146852 5646 146904 5652
rect 147968 5574 147996 8092
rect 149164 5574 149192 8092
rect 145748 5568 145800 5574
rect 145748 5510 145800 5516
rect 146852 5568 146904 5574
rect 146852 5510 146904 5516
rect 147956 5568 148008 5574
rect 147956 5510 148008 5516
rect 148048 5568 148100 5574
rect 148048 5510 148100 5516
rect 149152 5568 149204 5574
rect 149152 5510 149204 5516
rect 146864 480 146892 5510
rect 148060 480 148088 5510
rect 150268 3534 150296 8092
rect 151372 3534 151400 8092
rect 152568 5574 152596 8092
rect 153672 5574 153700 8092
rect 154776 5574 154804 8092
rect 155972 5574 156000 8092
rect 151544 5568 151596 5574
rect 151544 5510 151596 5516
rect 152556 5568 152608 5574
rect 152556 5510 152608 5516
rect 152740 5568 152792 5574
rect 152740 5510 152792 5516
rect 153660 5568 153712 5574
rect 153660 5510 153712 5516
rect 153936 5568 153988 5574
rect 153936 5510 153988 5516
rect 154764 5568 154816 5574
rect 154764 5510 154816 5516
rect 155132 5568 155184 5574
rect 155132 5510 155184 5516
rect 155960 5568 156012 5574
rect 155960 5510 156012 5516
rect 149244 3528 149296 3534
rect 149244 3470 149296 3476
rect 150256 3528 150308 3534
rect 150256 3470 150308 3476
rect 150440 3528 150492 3534
rect 150440 3470 150492 3476
rect 151360 3528 151412 3534
rect 151360 3470 151412 3476
rect 149256 480 149284 3470
rect 150452 480 150480 3470
rect 151556 480 151584 5510
rect 152752 480 152780 5510
rect 153948 480 153976 5510
rect 155144 480 155172 5510
rect 157076 3534 157104 8092
rect 157536 8078 158194 8106
rect 158732 8078 159390 8106
rect 160112 8078 160494 8106
rect 161492 8078 161598 8106
rect 162320 8078 162702 8106
rect 163516 8078 163898 8106
rect 164712 8078 165002 8106
rect 165908 8078 166106 8106
rect 167104 8078 167302 8106
rect 156328 3528 156380 3534
rect 156328 3470 156380 3476
rect 157064 3528 157116 3534
rect 157064 3470 157116 3476
rect 156340 480 156368 3470
rect 157536 480 157564 8078
rect 158732 480 158760 8078
rect 160112 5556 160140 8078
rect 161492 5658 161520 8078
rect 160020 5528 160140 5556
rect 161124 5630 161520 5658
rect 160020 626 160048 5528
rect 159928 598 160048 626
rect 159928 480 159956 598
rect 161124 480 161152 5630
rect 162320 480 162348 8078
rect 162822 6012 163386 6032
rect 162822 6010 162836 6012
rect 162892 6010 162916 6012
rect 162972 6010 162996 6012
rect 163052 6010 163076 6012
rect 163132 6010 163156 6012
rect 163212 6010 163236 6012
rect 163292 6010 163316 6012
rect 163372 6010 163386 6012
rect 163066 5958 163076 6010
rect 163132 5958 163142 6010
rect 162822 5956 162836 5958
rect 162892 5956 162916 5958
rect 162972 5956 162996 5958
rect 163052 5956 163076 5958
rect 163132 5956 163156 5958
rect 163212 5956 163236 5958
rect 163292 5956 163316 5958
rect 163372 5956 163386 5958
rect 162822 5936 163386 5956
rect 162822 4924 163386 4944
rect 162822 4922 162836 4924
rect 162892 4922 162916 4924
rect 162972 4922 162996 4924
rect 163052 4922 163076 4924
rect 163132 4922 163156 4924
rect 163212 4922 163236 4924
rect 163292 4922 163316 4924
rect 163372 4922 163386 4924
rect 163066 4870 163076 4922
rect 163132 4870 163142 4922
rect 162822 4868 162836 4870
rect 162892 4868 162916 4870
rect 162972 4868 162996 4870
rect 163052 4868 163076 4870
rect 163132 4868 163156 4870
rect 163212 4868 163236 4870
rect 163292 4868 163316 4870
rect 163372 4868 163386 4870
rect 162822 4848 163386 4868
rect 162822 3836 163386 3856
rect 162822 3834 162836 3836
rect 162892 3834 162916 3836
rect 162972 3834 162996 3836
rect 163052 3834 163076 3836
rect 163132 3834 163156 3836
rect 163212 3834 163236 3836
rect 163292 3834 163316 3836
rect 163372 3834 163386 3836
rect 163066 3782 163076 3834
rect 163132 3782 163142 3834
rect 162822 3780 162836 3782
rect 162892 3780 162916 3782
rect 162972 3780 162996 3782
rect 163052 3780 163076 3782
rect 163132 3780 163156 3782
rect 163212 3780 163236 3782
rect 163292 3780 163316 3782
rect 163372 3780 163386 3782
rect 162822 3760 163386 3780
rect 162822 2748 163386 2768
rect 162822 2746 162836 2748
rect 162892 2746 162916 2748
rect 162972 2746 162996 2748
rect 163052 2746 163076 2748
rect 163132 2746 163156 2748
rect 163212 2746 163236 2748
rect 163292 2746 163316 2748
rect 163372 2746 163386 2748
rect 163066 2694 163076 2746
rect 163132 2694 163142 2746
rect 162822 2692 162836 2694
rect 162892 2692 162916 2694
rect 162972 2692 162996 2694
rect 163052 2692 163076 2694
rect 163132 2692 163156 2694
rect 163212 2692 163236 2694
rect 163292 2692 163316 2694
rect 163372 2692 163386 2694
rect 162822 2672 163386 2692
rect 163516 480 163544 8078
rect 164712 480 164740 8078
rect 165908 480 165936 8078
rect 167104 480 167132 8078
rect 168392 5658 168420 8092
rect 168300 5630 168420 5658
rect 169404 8078 169510 8106
rect 170600 8078 170706 8106
rect 168300 626 168328 5630
rect 168208 598 168328 626
rect 168208 480 168236 598
rect 169404 480 169432 8078
rect 170600 480 170628 8078
rect 171796 480 171824 8092
rect 172914 8078 173020 8106
rect 174110 8078 174216 8106
rect 172992 480 173020 8078
rect 174188 480 174216 8078
rect 175200 5658 175228 8092
rect 176318 8078 176608 8106
rect 177514 8078 177804 8106
rect 178618 8078 179000 8106
rect 179722 8078 180196 8106
rect 180918 8078 181484 8106
rect 175200 5630 175320 5658
rect 175292 626 175320 5630
rect 175292 598 175412 626
rect 175384 480 175412 598
rect 176580 480 176608 8078
rect 177776 480 177804 8078
rect 178972 480 179000 8078
rect 180168 480 180196 8078
rect 180822 5468 181386 5488
rect 180822 5466 180836 5468
rect 180892 5466 180916 5468
rect 180972 5466 180996 5468
rect 181052 5466 181076 5468
rect 181132 5466 181156 5468
rect 181212 5466 181236 5468
rect 181292 5466 181316 5468
rect 181372 5466 181386 5468
rect 181066 5414 181076 5466
rect 181132 5414 181142 5466
rect 180822 5412 180836 5414
rect 180892 5412 180916 5414
rect 180972 5412 180996 5414
rect 181052 5412 181076 5414
rect 181132 5412 181156 5414
rect 181212 5412 181236 5414
rect 181292 5412 181316 5414
rect 181372 5412 181386 5414
rect 180822 5392 181386 5412
rect 180822 4380 181386 4400
rect 180822 4378 180836 4380
rect 180892 4378 180916 4380
rect 180972 4378 180996 4380
rect 181052 4378 181076 4380
rect 181132 4378 181156 4380
rect 181212 4378 181236 4380
rect 181292 4378 181316 4380
rect 181372 4378 181386 4380
rect 181066 4326 181076 4378
rect 181132 4326 181142 4378
rect 180822 4324 180836 4326
rect 180892 4324 180916 4326
rect 180972 4324 180996 4326
rect 181052 4324 181076 4326
rect 181132 4324 181156 4326
rect 181212 4324 181236 4326
rect 181292 4324 181316 4326
rect 181372 4324 181386 4326
rect 180822 4304 181386 4324
rect 180822 3292 181386 3312
rect 180822 3290 180836 3292
rect 180892 3290 180916 3292
rect 180972 3290 180996 3292
rect 181052 3290 181076 3292
rect 181132 3290 181156 3292
rect 181212 3290 181236 3292
rect 181292 3290 181316 3292
rect 181372 3290 181386 3292
rect 181066 3238 181076 3290
rect 181132 3238 181142 3290
rect 180822 3236 180836 3238
rect 180892 3236 180916 3238
rect 180972 3236 180996 3238
rect 181052 3236 181076 3238
rect 181132 3236 181156 3238
rect 181212 3236 181236 3238
rect 181292 3236 181316 3238
rect 181372 3236 181386 3238
rect 180822 3216 181386 3236
rect 180822 2204 181386 2224
rect 180822 2202 180836 2204
rect 180892 2202 180916 2204
rect 180972 2202 180996 2204
rect 181052 2202 181076 2204
rect 181132 2202 181156 2204
rect 181212 2202 181236 2204
rect 181292 2202 181316 2204
rect 181372 2202 181386 2204
rect 181066 2150 181076 2202
rect 181132 2150 181142 2202
rect 180822 2148 180836 2150
rect 180892 2148 180916 2150
rect 180972 2148 180996 2150
rect 181052 2148 181076 2150
rect 181132 2148 181156 2150
rect 181212 2148 181236 2150
rect 181292 2148 181316 2150
rect 181372 2148 181386 2150
rect 180822 2128 181386 2148
rect 181456 1986 181484 8078
rect 182008 5574 182036 8092
rect 183112 5574 183140 8092
rect 184322 8078 184888 8106
rect 185426 8078 186084 8106
rect 186530 8078 187280 8106
rect 181996 5568 182048 5574
rect 181996 5510 182048 5516
rect 182548 5568 182600 5574
rect 182548 5510 182600 5516
rect 183100 5568 183152 5574
rect 183100 5510 183152 5516
rect 183744 5568 183796 5574
rect 183744 5510 183796 5516
rect 181364 1958 181484 1986
rect 181364 480 181392 1958
rect 182560 480 182588 5510
rect 183756 480 183784 5510
rect 184860 480 184888 8078
rect 186056 480 186084 8078
rect 187252 480 187280 8078
rect 187712 3534 187740 8092
rect 188816 5574 188844 8092
rect 189920 5574 189948 8092
rect 191116 5574 191144 8092
rect 192220 5574 192248 8092
rect 188804 5568 188856 5574
rect 188804 5510 188856 5516
rect 189632 5568 189684 5574
rect 189632 5510 189684 5516
rect 189908 5568 189960 5574
rect 189908 5510 189960 5516
rect 190828 5568 190880 5574
rect 190828 5510 190880 5516
rect 191104 5568 191156 5574
rect 191104 5510 191156 5516
rect 192024 5568 192076 5574
rect 192024 5510 192076 5516
rect 192208 5568 192260 5574
rect 192208 5510 192260 5516
rect 193220 5568 193272 5574
rect 193220 5510 193272 5516
rect 187700 3528 187752 3534
rect 187700 3470 187752 3476
rect 188436 3528 188488 3534
rect 188436 3470 188488 3476
rect 188448 480 188476 3470
rect 189644 480 189672 5510
rect 190840 480 190868 5510
rect 192036 480 192064 5510
rect 193232 480 193260 5510
rect 193324 3534 193352 8092
rect 194520 5574 194548 8092
rect 195624 5710 195652 8092
rect 195612 5704 195664 5710
rect 195612 5646 195664 5652
rect 196728 5574 196756 8092
rect 196808 5704 196860 5710
rect 196808 5646 196860 5652
rect 194508 5568 194560 5574
rect 194508 5510 194560 5516
rect 195612 5568 195664 5574
rect 195612 5510 195664 5516
rect 196716 5568 196768 5574
rect 196716 5510 196768 5516
rect 193312 3528 193364 3534
rect 193312 3470 193364 3476
rect 194416 3528 194468 3534
rect 194416 3470 194468 3476
rect 194428 480 194456 3470
rect 195624 480 195652 5510
rect 196820 480 196848 5646
rect 197924 5642 197952 8092
rect 199028 6186 199056 8092
rect 199016 6180 199068 6186
rect 199016 6122 199068 6128
rect 198822 6012 199386 6032
rect 198822 6010 198836 6012
rect 198892 6010 198916 6012
rect 198972 6010 198996 6012
rect 199052 6010 199076 6012
rect 199132 6010 199156 6012
rect 199212 6010 199236 6012
rect 199292 6010 199316 6012
rect 199372 6010 199386 6012
rect 199066 5958 199076 6010
rect 199132 5958 199142 6010
rect 198822 5956 198836 5958
rect 198892 5956 198916 5958
rect 198972 5956 198996 5958
rect 199052 5956 199076 5958
rect 199132 5956 199156 5958
rect 199212 5956 199236 5958
rect 199292 5956 199316 5958
rect 199372 5956 199386 5958
rect 198822 5936 199386 5956
rect 197912 5636 197964 5642
rect 197912 5578 197964 5584
rect 198740 5636 198792 5642
rect 198740 5578 198792 5584
rect 198004 5568 198056 5574
rect 198004 5510 198056 5516
rect 198016 480 198044 5510
rect 198752 2530 198780 5578
rect 200132 5574 200160 8092
rect 200396 6180 200448 6186
rect 200396 6122 200448 6128
rect 200120 5568 200172 5574
rect 200120 5510 200172 5516
rect 198822 4924 199386 4944
rect 198822 4922 198836 4924
rect 198892 4922 198916 4924
rect 198972 4922 198996 4924
rect 199052 4922 199076 4924
rect 199132 4922 199156 4924
rect 199212 4922 199236 4924
rect 199292 4922 199316 4924
rect 199372 4922 199386 4924
rect 199066 4870 199076 4922
rect 199132 4870 199142 4922
rect 198822 4868 198836 4870
rect 198892 4868 198916 4870
rect 198972 4868 198996 4870
rect 199052 4868 199076 4870
rect 199132 4868 199156 4870
rect 199212 4868 199236 4870
rect 199292 4868 199316 4870
rect 199372 4868 199386 4870
rect 198822 4848 199386 4868
rect 198822 3836 199386 3856
rect 198822 3834 198836 3836
rect 198892 3834 198916 3836
rect 198972 3834 198996 3836
rect 199052 3834 199076 3836
rect 199132 3834 199156 3836
rect 199212 3834 199236 3836
rect 199292 3834 199316 3836
rect 199372 3834 199386 3836
rect 199066 3782 199076 3834
rect 199132 3782 199142 3834
rect 198822 3780 198836 3782
rect 198892 3780 198916 3782
rect 198972 3780 198996 3782
rect 199052 3780 199076 3782
rect 199132 3780 199156 3782
rect 199212 3780 199236 3782
rect 199292 3780 199316 3782
rect 199372 3780 199386 3782
rect 198822 3760 199386 3780
rect 198822 2748 199386 2768
rect 198822 2746 198836 2748
rect 198892 2746 198916 2748
rect 198972 2746 198996 2748
rect 199052 2746 199076 2748
rect 199132 2746 199156 2748
rect 199212 2746 199236 2748
rect 199292 2746 199316 2748
rect 199372 2746 199386 2748
rect 199066 2694 199076 2746
rect 199132 2694 199142 2746
rect 198822 2692 198836 2694
rect 198892 2692 198916 2694
rect 198972 2692 198996 2694
rect 199052 2692 199076 2694
rect 199132 2692 199156 2694
rect 199212 2692 199236 2694
rect 199292 2692 199316 2694
rect 199372 2692 199386 2694
rect 198822 2672 199386 2692
rect 198752 2502 199240 2530
rect 199212 480 199240 2502
rect 200408 480 200436 6122
rect 201236 5642 201264 8092
rect 201224 5636 201276 5642
rect 201224 5578 201276 5584
rect 202432 5574 202460 8092
rect 203536 5642 203564 8092
rect 202696 5636 202748 5642
rect 202696 5578 202748 5584
rect 203524 5636 203576 5642
rect 203524 5578 203576 5584
rect 201500 5568 201552 5574
rect 201500 5510 201552 5516
rect 202420 5568 202472 5574
rect 202420 5510 202472 5516
rect 201512 480 201540 5510
rect 202708 480 202736 5578
rect 204640 5574 204668 8092
rect 205836 5642 205864 8092
rect 206940 5710 206968 8092
rect 206928 5704 206980 5710
rect 206928 5646 206980 5652
rect 205088 5636 205140 5642
rect 205088 5578 205140 5584
rect 205824 5636 205876 5642
rect 205824 5578 205876 5584
rect 207480 5636 207532 5642
rect 207480 5578 207532 5584
rect 203892 5568 203944 5574
rect 203892 5510 203944 5516
rect 204628 5568 204680 5574
rect 204628 5510 204680 5516
rect 203904 480 203932 5510
rect 205100 480 205128 5578
rect 206284 5568 206336 5574
rect 206284 5510 206336 5516
rect 206296 480 206324 5510
rect 207492 480 207520 5578
rect 208044 5574 208072 8092
rect 208676 5704 208728 5710
rect 208676 5646 208728 5652
rect 208032 5568 208084 5574
rect 208032 5510 208084 5516
rect 208688 480 208716 5646
rect 209240 5642 209268 8092
rect 209228 5636 209280 5642
rect 209228 5578 209280 5584
rect 210344 5574 210372 8092
rect 211448 5642 211476 8092
rect 211068 5636 211120 5642
rect 211068 5578 211120 5584
rect 211436 5636 211488 5642
rect 211436 5578 211488 5584
rect 209872 5568 209924 5574
rect 209872 5510 209924 5516
rect 210332 5568 210384 5574
rect 210332 5510 210384 5516
rect 209884 480 209912 5510
rect 211080 480 211108 5578
rect 212644 5574 212672 8092
rect 213748 5642 213776 8092
rect 214852 5710 214880 8092
rect 214840 5704 214892 5710
rect 214840 5646 214892 5652
rect 213460 5636 213512 5642
rect 213460 5578 213512 5584
rect 213736 5636 213788 5642
rect 213736 5578 213788 5584
rect 215852 5636 215904 5642
rect 215852 5578 215904 5584
rect 212264 5568 212316 5574
rect 212264 5510 212316 5516
rect 212632 5568 212684 5574
rect 212632 5510 212684 5516
rect 212276 480 212304 5510
rect 213472 480 213500 5578
rect 214656 5568 214708 5574
rect 214656 5510 214708 5516
rect 214668 480 214696 5510
rect 215864 480 215892 5578
rect 216048 5574 216076 8092
rect 216680 5704 216732 5710
rect 216680 5646 216732 5652
rect 216036 5568 216088 5574
rect 216036 5510 216088 5516
rect 216692 1986 216720 5646
rect 217152 5642 217180 8092
rect 217140 5636 217192 5642
rect 217140 5578 217192 5584
rect 218256 5574 218284 8092
rect 219452 5642 219480 8092
rect 220556 5710 220584 8092
rect 220544 5704 220596 5710
rect 220544 5646 220596 5652
rect 219348 5636 219400 5642
rect 219348 5578 219400 5584
rect 219440 5636 219492 5642
rect 219440 5578 219492 5584
rect 218152 5568 218204 5574
rect 218152 5510 218204 5516
rect 218244 5568 218296 5574
rect 218244 5510 218296 5516
rect 216822 5468 217386 5488
rect 216822 5466 216836 5468
rect 216892 5466 216916 5468
rect 216972 5466 216996 5468
rect 217052 5466 217076 5468
rect 217132 5466 217156 5468
rect 217212 5466 217236 5468
rect 217292 5466 217316 5468
rect 217372 5466 217386 5468
rect 217066 5414 217076 5466
rect 217132 5414 217142 5466
rect 216822 5412 216836 5414
rect 216892 5412 216916 5414
rect 216972 5412 216996 5414
rect 217052 5412 217076 5414
rect 217132 5412 217156 5414
rect 217212 5412 217236 5414
rect 217292 5412 217316 5414
rect 217372 5412 217386 5414
rect 216822 5392 217386 5412
rect 216822 4380 217386 4400
rect 216822 4378 216836 4380
rect 216892 4378 216916 4380
rect 216972 4378 216996 4380
rect 217052 4378 217076 4380
rect 217132 4378 217156 4380
rect 217212 4378 217236 4380
rect 217292 4378 217316 4380
rect 217372 4378 217386 4380
rect 217066 4326 217076 4378
rect 217132 4326 217142 4378
rect 216822 4324 216836 4326
rect 216892 4324 216916 4326
rect 216972 4324 216996 4326
rect 217052 4324 217076 4326
rect 217132 4324 217156 4326
rect 217212 4324 217236 4326
rect 217292 4324 217316 4326
rect 217372 4324 217386 4326
rect 216822 4304 217386 4324
rect 216822 3292 217386 3312
rect 216822 3290 216836 3292
rect 216892 3290 216916 3292
rect 216972 3290 216996 3292
rect 217052 3290 217076 3292
rect 217132 3290 217156 3292
rect 217212 3290 217236 3292
rect 217292 3290 217316 3292
rect 217372 3290 217386 3292
rect 217066 3238 217076 3290
rect 217132 3238 217142 3290
rect 216822 3236 216836 3238
rect 216892 3236 216916 3238
rect 216972 3236 216996 3238
rect 217052 3236 217076 3238
rect 217132 3236 217156 3238
rect 217212 3236 217236 3238
rect 217292 3236 217316 3238
rect 217372 3236 217386 3238
rect 216822 3216 217386 3236
rect 216822 2204 217386 2224
rect 216822 2202 216836 2204
rect 216892 2202 216916 2204
rect 216972 2202 216996 2204
rect 217052 2202 217076 2204
rect 217132 2202 217156 2204
rect 217212 2202 217236 2204
rect 217292 2202 217316 2204
rect 217372 2202 217386 2204
rect 217066 2150 217076 2202
rect 217132 2150 217142 2202
rect 216822 2148 216836 2150
rect 216892 2148 216916 2150
rect 216972 2148 216996 2150
rect 217052 2148 217076 2150
rect 217132 2148 217156 2150
rect 217212 2148 217236 2150
rect 217292 2148 217316 2150
rect 217372 2148 217386 2150
rect 216822 2128 217386 2148
rect 216692 1958 217088 1986
rect 217060 480 217088 1958
rect 218164 480 218192 5510
rect 219360 480 219388 5578
rect 221660 5574 221688 8092
rect 222856 5642 222884 8092
rect 223960 5710 223988 8092
rect 222936 5704 222988 5710
rect 222936 5646 222988 5652
rect 223948 5704 224000 5710
rect 223948 5646 224000 5652
rect 221740 5636 221792 5642
rect 221740 5578 221792 5584
rect 222844 5636 222896 5642
rect 222844 5578 222896 5584
rect 220544 5568 220596 5574
rect 220544 5510 220596 5516
rect 221648 5568 221700 5574
rect 221648 5510 221700 5516
rect 220556 480 220584 5510
rect 221752 480 221780 5578
rect 222948 480 222976 5646
rect 225064 5574 225092 8092
rect 226260 5778 226288 8092
rect 226248 5772 226300 5778
rect 226248 5714 226300 5720
rect 226524 5704 226576 5710
rect 226524 5646 226576 5652
rect 225328 5636 225380 5642
rect 225328 5578 225380 5584
rect 224132 5568 224184 5574
rect 224132 5510 224184 5516
rect 225052 5568 225104 5574
rect 225052 5510 225104 5516
rect 224144 480 224172 5510
rect 225340 480 225368 5578
rect 226536 480 226564 5646
rect 227364 5642 227392 8092
rect 228468 5710 228496 8092
rect 228916 5772 228968 5778
rect 228916 5714 228968 5720
rect 228456 5704 228508 5710
rect 228456 5646 228508 5652
rect 227352 5636 227404 5642
rect 227352 5578 227404 5584
rect 227720 5568 227772 5574
rect 227720 5510 227772 5516
rect 227732 480 227760 5510
rect 228928 480 228956 5714
rect 229664 5574 229692 8092
rect 230768 5642 230796 8092
rect 231872 5710 231900 8092
rect 231308 5704 231360 5710
rect 231308 5646 231360 5652
rect 231860 5704 231912 5710
rect 231860 5646 231912 5652
rect 230112 5636 230164 5642
rect 230112 5578 230164 5584
rect 230756 5636 230808 5642
rect 230756 5578 230808 5584
rect 229652 5568 229704 5574
rect 229652 5510 229704 5516
rect 230124 480 230152 5578
rect 231320 480 231348 5646
rect 233068 5574 233096 8092
rect 234172 5778 234200 8092
rect 235276 6186 235304 8092
rect 235264 6180 235316 6186
rect 235264 6122 235316 6128
rect 234822 6012 235386 6032
rect 234822 6010 234836 6012
rect 234892 6010 234916 6012
rect 234972 6010 234996 6012
rect 235052 6010 235076 6012
rect 235132 6010 235156 6012
rect 235212 6010 235236 6012
rect 235292 6010 235316 6012
rect 235372 6010 235386 6012
rect 235066 5958 235076 6010
rect 235132 5958 235142 6010
rect 234822 5956 234836 5958
rect 234892 5956 234916 5958
rect 234972 5956 234996 5958
rect 235052 5956 235076 5958
rect 235132 5956 235156 5958
rect 235212 5956 235236 5958
rect 235292 5956 235316 5958
rect 235372 5956 235386 5958
rect 234822 5936 235386 5956
rect 234160 5772 234212 5778
rect 234160 5714 234212 5720
rect 234712 5704 234764 5710
rect 234712 5646 234764 5652
rect 233700 5636 233752 5642
rect 233700 5578 233752 5584
rect 232504 5568 232556 5574
rect 232504 5510 232556 5516
rect 233056 5568 233108 5574
rect 233056 5510 233108 5516
rect 232516 480 232544 5510
rect 233712 480 233740 5578
rect 234724 2530 234752 5646
rect 236380 5642 236408 8092
rect 237196 5772 237248 5778
rect 237196 5714 237248 5720
rect 236368 5636 236420 5642
rect 236368 5578 236420 5584
rect 235908 5568 235960 5574
rect 235908 5510 235960 5516
rect 234822 4924 235386 4944
rect 234822 4922 234836 4924
rect 234892 4922 234916 4924
rect 234972 4922 234996 4924
rect 235052 4922 235076 4924
rect 235132 4922 235156 4924
rect 235212 4922 235236 4924
rect 235292 4922 235316 4924
rect 235372 4922 235386 4924
rect 235066 4870 235076 4922
rect 235132 4870 235142 4922
rect 234822 4868 234836 4870
rect 234892 4868 234916 4870
rect 234972 4868 234996 4870
rect 235052 4868 235076 4870
rect 235132 4868 235156 4870
rect 235212 4868 235236 4870
rect 235292 4868 235316 4870
rect 235372 4868 235386 4870
rect 234822 4848 235386 4868
rect 234822 3836 235386 3856
rect 234822 3834 234836 3836
rect 234892 3834 234916 3836
rect 234972 3834 234996 3836
rect 235052 3834 235076 3836
rect 235132 3834 235156 3836
rect 235212 3834 235236 3836
rect 235292 3834 235316 3836
rect 235372 3834 235386 3836
rect 235066 3782 235076 3834
rect 235132 3782 235142 3834
rect 234822 3780 234836 3782
rect 234892 3780 234916 3782
rect 234972 3780 234996 3782
rect 235052 3780 235076 3782
rect 235132 3780 235156 3782
rect 235212 3780 235236 3782
rect 235292 3780 235316 3782
rect 235372 3780 235386 3782
rect 234822 3760 235386 3780
rect 235920 3482 235948 5510
rect 235920 3454 236040 3482
rect 234822 2748 235386 2768
rect 234822 2746 234836 2748
rect 234892 2746 234916 2748
rect 234972 2746 234996 2748
rect 235052 2746 235076 2748
rect 235132 2746 235156 2748
rect 235212 2746 235236 2748
rect 235292 2746 235316 2748
rect 235372 2746 235386 2748
rect 235066 2694 235076 2746
rect 235132 2694 235142 2746
rect 234822 2692 234836 2694
rect 234892 2692 234916 2694
rect 234972 2692 234996 2694
rect 235052 2692 235076 2694
rect 235132 2692 235156 2694
rect 235212 2692 235236 2694
rect 235292 2692 235316 2694
rect 235372 2692 235386 2694
rect 234822 2672 235386 2692
rect 234724 2502 234844 2530
rect 234816 480 234844 2502
rect 236012 480 236040 3454
rect 237208 480 237236 5714
rect 237576 5574 237604 8092
rect 238392 6180 238444 6186
rect 238392 6122 238444 6128
rect 237564 5568 237616 5574
rect 237564 5510 237616 5516
rect 238404 480 238432 6122
rect 238680 5846 238708 8092
rect 238668 5840 238720 5846
rect 238668 5782 238720 5788
rect 239784 5642 239812 8092
rect 240140 5840 240192 5846
rect 240140 5782 240192 5788
rect 239588 5636 239640 5642
rect 239588 5578 239640 5584
rect 239772 5636 239824 5642
rect 239772 5578 239824 5584
rect 239600 480 239628 5578
rect 240152 2922 240180 5782
rect 240980 5574 241008 8092
rect 242084 5710 242112 8092
rect 243188 5778 243216 8092
rect 243176 5772 243228 5778
rect 243176 5714 243228 5720
rect 242072 5704 242124 5710
rect 242072 5646 242124 5652
rect 244384 5642 244412 8092
rect 245488 6118 245516 8092
rect 245476 6112 245528 6118
rect 245476 6054 245528 6060
rect 245568 5704 245620 5710
rect 245568 5646 245620 5652
rect 242808 5636 242860 5642
rect 242808 5578 242860 5584
rect 244372 5636 244424 5642
rect 244372 5578 244424 5584
rect 240784 5568 240836 5574
rect 240784 5510 240836 5516
rect 240968 5568 241020 5574
rect 240968 5510 241020 5516
rect 240140 2916 240192 2922
rect 240140 2858 240192 2864
rect 240796 480 240824 5510
rect 242820 3482 242848 5578
rect 244188 5568 244240 5574
rect 244188 5510 244240 5516
rect 244200 3482 244228 5510
rect 242820 3454 243216 3482
rect 244200 3454 244412 3482
rect 241980 2916 242032 2922
rect 241980 2858 242032 2864
rect 241992 480 242020 2858
rect 243188 480 243216 3454
rect 244384 480 244412 3454
rect 245580 480 245608 5646
rect 246592 5574 246620 8092
rect 247040 6112 247092 6118
rect 247040 6054 247092 6060
rect 246764 5772 246816 5778
rect 246764 5714 246816 5720
rect 246580 5568 246632 5574
rect 246580 5510 246632 5516
rect 246776 480 246804 5714
rect 247052 4078 247080 6054
rect 247788 5778 247816 8092
rect 247776 5772 247828 5778
rect 247776 5714 247828 5720
rect 248892 5642 248920 8092
rect 249996 5710 250024 8092
rect 251088 5772 251140 5778
rect 251088 5714 251140 5720
rect 249984 5704 250036 5710
rect 249984 5646 250036 5652
rect 247960 5636 248012 5642
rect 247960 5578 248012 5584
rect 248880 5636 248932 5642
rect 248880 5578 248932 5584
rect 247040 4072 247092 4078
rect 247040 4014 247092 4020
rect 247972 480 248000 5578
rect 249248 5568 249300 5574
rect 249248 5510 249300 5516
rect 249156 4072 249208 4078
rect 249156 4014 249208 4020
rect 249168 480 249196 4014
rect 249260 2922 249288 5510
rect 251100 3210 251128 5714
rect 251192 5574 251220 8092
rect 252296 5778 252324 8092
rect 252284 5772 252336 5778
rect 252284 5714 252336 5720
rect 253400 5642 253428 8092
rect 254596 6118 254624 8092
rect 254584 6112 254636 6118
rect 254584 6054 254636 6060
rect 254216 5772 254268 5778
rect 254216 5714 254268 5720
rect 253848 5704 253900 5710
rect 253848 5646 253900 5652
rect 252468 5636 252520 5642
rect 252468 5578 252520 5584
rect 253388 5636 253440 5642
rect 253388 5578 253440 5584
rect 251180 5568 251232 5574
rect 251180 5510 251232 5516
rect 252480 3482 252508 5578
rect 252822 5468 253386 5488
rect 252822 5466 252836 5468
rect 252892 5466 252916 5468
rect 252972 5466 252996 5468
rect 253052 5466 253076 5468
rect 253132 5466 253156 5468
rect 253212 5466 253236 5468
rect 253292 5466 253316 5468
rect 253372 5466 253386 5468
rect 253066 5414 253076 5466
rect 253132 5414 253142 5466
rect 252822 5412 252836 5414
rect 252892 5412 252916 5414
rect 252972 5412 252996 5414
rect 253052 5412 253076 5414
rect 253132 5412 253156 5414
rect 253212 5412 253236 5414
rect 253292 5412 253316 5414
rect 253372 5412 253386 5414
rect 252822 5392 253386 5412
rect 252822 4380 253386 4400
rect 252822 4378 252836 4380
rect 252892 4378 252916 4380
rect 252972 4378 252996 4380
rect 253052 4378 253076 4380
rect 253132 4378 253156 4380
rect 253212 4378 253236 4380
rect 253292 4378 253316 4380
rect 253372 4378 253386 4380
rect 253066 4326 253076 4378
rect 253132 4326 253142 4378
rect 252822 4324 252836 4326
rect 252892 4324 252916 4326
rect 252972 4324 252996 4326
rect 253052 4324 253076 4326
rect 253132 4324 253156 4326
rect 253212 4324 253236 4326
rect 253292 4324 253316 4326
rect 253372 4324 253386 4326
rect 252822 4304 253386 4324
rect 252480 3454 252692 3482
rect 251100 3182 251496 3210
rect 249248 2916 249300 2922
rect 249248 2858 249300 2864
rect 250352 2916 250404 2922
rect 250352 2858 250404 2864
rect 250364 480 250392 2858
rect 251468 480 251496 3182
rect 252664 480 252692 3454
rect 252822 3292 253386 3312
rect 252822 3290 252836 3292
rect 252892 3290 252916 3292
rect 252972 3290 252996 3292
rect 253052 3290 253076 3292
rect 253132 3290 253156 3292
rect 253212 3290 253236 3292
rect 253292 3290 253316 3292
rect 253372 3290 253386 3292
rect 253066 3238 253076 3290
rect 253132 3238 253142 3290
rect 252822 3236 252836 3238
rect 252892 3236 252916 3238
rect 252972 3236 252996 3238
rect 253052 3236 253076 3238
rect 253132 3236 253156 3238
rect 253212 3236 253236 3238
rect 253292 3236 253316 3238
rect 253372 3236 253386 3238
rect 252822 3216 253386 3236
rect 252822 2204 253386 2224
rect 252822 2202 252836 2204
rect 252892 2202 252916 2204
rect 252972 2202 252996 2204
rect 253052 2202 253076 2204
rect 253132 2202 253156 2204
rect 253212 2202 253236 2204
rect 253292 2202 253316 2204
rect 253372 2202 253386 2204
rect 253066 2150 253076 2202
rect 253132 2150 253142 2202
rect 252822 2148 252836 2150
rect 252892 2148 252916 2150
rect 252972 2148 252996 2150
rect 253052 2148 253076 2150
rect 253132 2148 253156 2150
rect 253212 2148 253236 2150
rect 253292 2148 253316 2150
rect 253372 2148 253386 2150
rect 252822 2128 253386 2148
rect 253860 480 253888 5646
rect 254228 3466 254256 5714
rect 255412 5636 255464 5642
rect 255412 5578 255464 5584
rect 255044 5568 255096 5574
rect 255044 5510 255096 5516
rect 254216 3460 254268 3466
rect 254216 3402 254268 3408
rect 255056 480 255084 5510
rect 255424 3534 255452 5578
rect 255700 5574 255728 8092
rect 256700 6112 256752 6118
rect 256700 6054 256752 6060
rect 255688 5568 255740 5574
rect 255688 5510 255740 5516
rect 256712 4078 256740 6054
rect 256804 5642 256832 8092
rect 258000 5846 258028 8092
rect 257988 5840 258040 5846
rect 257988 5782 258040 5788
rect 256792 5636 256844 5642
rect 256792 5578 256844 5584
rect 259104 5574 259132 8092
rect 260104 5840 260156 5846
rect 260104 5782 260156 5788
rect 259000 5568 259052 5574
rect 259000 5510 259052 5516
rect 259092 5568 259144 5574
rect 259092 5510 259144 5516
rect 256700 4072 256752 4078
rect 256700 4014 256752 4020
rect 258632 4072 258684 4078
rect 258632 4014 258684 4020
rect 255412 3528 255464 3534
rect 255412 3470 255464 3476
rect 257436 3528 257488 3534
rect 257436 3470 257488 3476
rect 256240 3460 256292 3466
rect 256240 3402 256292 3408
rect 256252 480 256280 3402
rect 257448 480 257476 3470
rect 258644 480 258672 4014
rect 259012 2922 259040 5510
rect 260116 2990 260144 5782
rect 260208 5710 260236 8092
rect 260196 5704 260248 5710
rect 260196 5646 260248 5652
rect 261404 5642 261432 8092
rect 262508 5710 262536 8092
rect 262404 5704 262456 5710
rect 262404 5646 262456 5652
rect 262496 5704 262548 5710
rect 262496 5646 262548 5652
rect 260748 5636 260800 5642
rect 260748 5578 260800 5584
rect 261392 5636 261444 5642
rect 261392 5578 261444 5584
rect 260760 3074 260788 5578
rect 261208 5568 261260 5574
rect 261208 5510 261260 5516
rect 261220 3466 261248 5510
rect 262416 3534 262444 5646
rect 263612 5574 263640 8092
rect 264808 6254 264836 8092
rect 264796 6248 264848 6254
rect 264796 6190 264848 6196
rect 265912 5846 265940 8092
rect 266360 6248 266412 6254
rect 266360 6190 266412 6196
rect 265900 5840 265952 5846
rect 265900 5782 265952 5788
rect 264980 5704 265032 5710
rect 264980 5646 265032 5652
rect 263692 5636 263744 5642
rect 263692 5578 263744 5584
rect 263600 5568 263652 5574
rect 263600 5510 263652 5516
rect 262404 3528 262456 3534
rect 262404 3470 262456 3476
rect 263704 3466 263732 5578
rect 264992 3534 265020 5646
rect 266372 3738 266400 6190
rect 267016 5914 267044 8092
rect 267004 5908 267056 5914
rect 267004 5850 267056 5856
rect 268212 5574 268240 8092
rect 269028 5840 269080 5846
rect 269028 5782 269080 5788
rect 266452 5568 266504 5574
rect 266452 5510 266504 5516
rect 268200 5568 268252 5574
rect 268200 5510 268252 5516
rect 266464 4010 266492 5510
rect 266452 4004 266504 4010
rect 266452 3946 266504 3952
rect 268108 4004 268160 4010
rect 268108 3946 268160 3952
rect 266360 3732 266412 3738
rect 266360 3674 266412 3680
rect 264612 3528 264664 3534
rect 264612 3470 264664 3476
rect 264980 3528 265032 3534
rect 264980 3470 265032 3476
rect 267004 3528 267056 3534
rect 267004 3470 267056 3476
rect 261208 3460 261260 3466
rect 261208 3402 261260 3408
rect 263416 3460 263468 3466
rect 263416 3402 263468 3408
rect 263692 3460 263744 3466
rect 263692 3402 263744 3408
rect 260760 3046 261064 3074
rect 260104 2984 260156 2990
rect 260104 2926 260156 2932
rect 259000 2916 259052 2922
rect 259000 2858 259052 2864
rect 259828 2916 259880 2922
rect 259828 2858 259880 2864
rect 259840 480 259868 2858
rect 261036 480 261064 3046
rect 262220 2984 262272 2990
rect 262220 2926 262272 2932
rect 262232 480 262260 2926
rect 263428 480 263456 3402
rect 264624 480 264652 3470
rect 265808 3460 265860 3466
rect 265808 3402 265860 3408
rect 265820 480 265848 3402
rect 267016 480 267044 3470
rect 268120 480 268148 3946
rect 269040 2922 269068 5782
rect 269316 5642 269344 8092
rect 269672 5908 269724 5914
rect 269672 5850 269724 5856
rect 269304 5636 269356 5642
rect 269304 5578 269356 5584
rect 269304 3732 269356 3738
rect 269304 3674 269356 3680
rect 269028 2916 269080 2922
rect 269028 2858 269080 2864
rect 269316 480 269344 3674
rect 269684 3058 269712 5850
rect 270420 5710 270448 8092
rect 270822 6012 271386 6032
rect 270822 6010 270836 6012
rect 270892 6010 270916 6012
rect 270972 6010 270996 6012
rect 271052 6010 271076 6012
rect 271132 6010 271156 6012
rect 271212 6010 271236 6012
rect 271292 6010 271316 6012
rect 271372 6010 271386 6012
rect 271066 5958 271076 6010
rect 271132 5958 271142 6010
rect 270822 5956 270836 5958
rect 270892 5956 270916 5958
rect 270972 5956 270996 5958
rect 271052 5956 271076 5958
rect 271132 5956 271156 5958
rect 271212 5956 271236 5958
rect 271292 5956 271316 5958
rect 271372 5956 271386 5958
rect 270822 5936 271386 5956
rect 270408 5704 270460 5710
rect 270408 5646 270460 5652
rect 271616 5574 271644 8092
rect 272720 6390 272748 8092
rect 272708 6384 272760 6390
rect 272708 6326 272760 6332
rect 273824 6254 273852 8092
rect 273812 6248 273864 6254
rect 273812 6190 273864 6196
rect 272984 5704 273036 5710
rect 272984 5646 273036 5652
rect 271880 5636 271932 5642
rect 271880 5578 271932 5584
rect 270500 5568 270552 5574
rect 270500 5510 270552 5516
rect 271604 5568 271656 5574
rect 271604 5510 271656 5516
rect 270512 3466 270540 5510
rect 270822 4924 271386 4944
rect 270822 4922 270836 4924
rect 270892 4922 270916 4924
rect 270972 4922 270996 4924
rect 271052 4922 271076 4924
rect 271132 4922 271156 4924
rect 271212 4922 271236 4924
rect 271292 4922 271316 4924
rect 271372 4922 271386 4924
rect 271066 4870 271076 4922
rect 271132 4870 271142 4922
rect 270822 4868 270836 4870
rect 270892 4868 270916 4870
rect 270972 4868 270996 4870
rect 271052 4868 271076 4870
rect 271132 4868 271156 4870
rect 271212 4868 271236 4870
rect 271292 4868 271316 4870
rect 271372 4868 271386 4870
rect 270822 4848 271386 4868
rect 270822 3836 271386 3856
rect 270822 3834 270836 3836
rect 270892 3834 270916 3836
rect 270972 3834 270996 3836
rect 271052 3834 271076 3836
rect 271132 3834 271156 3836
rect 271212 3834 271236 3836
rect 271292 3834 271316 3836
rect 271372 3834 271386 3836
rect 271066 3782 271076 3834
rect 271132 3782 271142 3834
rect 270822 3780 270836 3782
rect 270892 3780 270916 3782
rect 270972 3780 270996 3782
rect 271052 3780 271076 3782
rect 271132 3780 271156 3782
rect 271212 3780 271236 3782
rect 271292 3780 271316 3782
rect 271372 3780 271386 3782
rect 270822 3760 271386 3780
rect 270500 3460 270552 3466
rect 270500 3402 270552 3408
rect 271892 3058 271920 5578
rect 272996 3466 273024 5646
rect 274928 5574 274956 8092
rect 275100 6384 275152 6390
rect 275100 6326 275152 6332
rect 273996 5568 274048 5574
rect 273996 5510 274048 5516
rect 274916 5568 274968 5574
rect 274916 5510 274968 5516
rect 272892 3460 272944 3466
rect 272892 3402 272944 3408
rect 272984 3460 273036 3466
rect 272984 3402 273036 3408
rect 269672 3052 269724 3058
rect 269672 2994 269724 3000
rect 271696 3052 271748 3058
rect 271696 2994 271748 3000
rect 271880 3052 271932 3058
rect 271880 2994 271932 3000
rect 270500 2916 270552 2922
rect 270500 2858 270552 2864
rect 270512 480 270540 2858
rect 270822 2748 271386 2768
rect 270822 2746 270836 2748
rect 270892 2746 270916 2748
rect 270972 2746 270996 2748
rect 271052 2746 271076 2748
rect 271132 2746 271156 2748
rect 271212 2746 271236 2748
rect 271292 2746 271316 2748
rect 271372 2746 271386 2748
rect 271066 2694 271076 2746
rect 271132 2694 271142 2746
rect 270822 2692 270836 2694
rect 270892 2692 270916 2694
rect 270972 2692 270996 2694
rect 271052 2692 271076 2694
rect 271132 2692 271156 2694
rect 271212 2692 271236 2694
rect 271292 2692 271316 2694
rect 271372 2692 271386 2694
rect 270822 2672 271386 2692
rect 271708 480 271736 2994
rect 272904 480 272932 3402
rect 274008 3194 274036 5510
rect 275112 3738 275140 6326
rect 276020 6248 276072 6254
rect 276020 6190 276072 6196
rect 276032 4078 276060 6190
rect 276124 5710 276152 8092
rect 277228 5778 277256 8092
rect 277216 5772 277268 5778
rect 277216 5714 277268 5720
rect 276112 5704 276164 5710
rect 276112 5646 276164 5652
rect 278332 5642 278360 8092
rect 279332 5704 279384 5710
rect 279332 5646 279384 5652
rect 278320 5636 278372 5642
rect 278320 5578 278372 5584
rect 278412 5568 278464 5574
rect 278412 5510 278464 5516
rect 276020 4072 276072 4078
rect 276020 4014 276072 4020
rect 275100 3732 275152 3738
rect 275100 3674 275152 3680
rect 277676 3732 277728 3738
rect 277676 3674 277728 3680
rect 275284 3460 275336 3466
rect 275284 3402 275336 3408
rect 273996 3188 274048 3194
rect 273996 3130 274048 3136
rect 274088 3052 274140 3058
rect 274088 2994 274140 3000
rect 274100 480 274128 2994
rect 275296 480 275324 3402
rect 276480 3188 276532 3194
rect 276480 3130 276532 3136
rect 276492 480 276520 3130
rect 277688 480 277716 3674
rect 278424 2854 278452 5510
rect 278872 4072 278924 4078
rect 278872 4014 278924 4020
rect 278412 2848 278464 2854
rect 278412 2790 278464 2796
rect 278884 480 278912 4014
rect 279344 3058 279372 5646
rect 279528 5574 279556 8092
rect 280632 5778 280660 8092
rect 279792 5772 279844 5778
rect 279792 5714 279844 5720
rect 280620 5772 280672 5778
rect 280620 5714 280672 5720
rect 279516 5568 279568 5574
rect 279516 5510 279568 5516
rect 279804 4146 279832 5714
rect 281736 5710 281764 8092
rect 282932 5846 282960 8092
rect 284036 6390 284064 8092
rect 284024 6384 284076 6390
rect 284024 6326 284076 6332
rect 282920 5840 282972 5846
rect 282920 5782 282972 5788
rect 283196 5772 283248 5778
rect 283196 5714 283248 5720
rect 281724 5704 281776 5710
rect 281724 5646 281776 5652
rect 280896 5636 280948 5642
rect 280896 5578 280948 5584
rect 279792 4140 279844 4146
rect 279792 4082 279844 4088
rect 280908 3398 280936 5578
rect 282092 5568 282144 5574
rect 282092 5510 282144 5516
rect 282104 3534 282132 5510
rect 282460 4140 282512 4146
rect 282460 4082 282512 4088
rect 282092 3528 282144 3534
rect 282092 3470 282144 3476
rect 280896 3392 280948 3398
rect 280896 3334 280948 3340
rect 279332 3052 279384 3058
rect 279332 2994 279384 3000
rect 281264 3052 281316 3058
rect 281264 2994 281316 3000
rect 280068 2848 280120 2854
rect 280068 2790 280120 2796
rect 280080 480 280108 2790
rect 281276 480 281304 2994
rect 282472 480 282500 4082
rect 283208 3194 283236 5714
rect 284392 5704 284444 5710
rect 284392 5646 284444 5652
rect 284404 4010 284432 5646
rect 285140 5574 285168 8092
rect 285680 6384 285732 6390
rect 285680 6326 285732 6332
rect 285128 5568 285180 5574
rect 285128 5510 285180 5516
rect 285692 4146 285720 6326
rect 286336 5846 286364 8092
rect 285772 5840 285824 5846
rect 285772 5782 285824 5788
rect 286324 5840 286376 5846
rect 286324 5782 286376 5788
rect 285680 4140 285732 4146
rect 285680 4082 285732 4088
rect 285784 4078 285812 5782
rect 287440 5642 287468 8092
rect 287428 5636 287480 5642
rect 287428 5578 287480 5584
rect 288544 5574 288572 8092
rect 289452 5840 289504 5846
rect 289452 5782 289504 5788
rect 288256 5568 288308 5574
rect 288256 5510 288308 5516
rect 288532 5568 288584 5574
rect 288532 5510 288584 5516
rect 285772 4072 285824 4078
rect 285772 4014 285824 4020
rect 284392 4004 284444 4010
rect 284392 3946 284444 3952
rect 287152 4004 287204 4010
rect 287152 3946 287204 3952
rect 284760 3528 284812 3534
rect 284760 3470 284812 3476
rect 283656 3392 283708 3398
rect 283656 3334 283708 3340
rect 283196 3188 283248 3194
rect 283196 3130 283248 3136
rect 283668 480 283696 3334
rect 284772 480 284800 3470
rect 285956 3188 286008 3194
rect 285956 3130 286008 3136
rect 285968 480 285996 3130
rect 287164 480 287192 3946
rect 288268 2922 288296 5510
rect 288822 5468 289386 5488
rect 288822 5466 288836 5468
rect 288892 5466 288916 5468
rect 288972 5466 288996 5468
rect 289052 5466 289076 5468
rect 289132 5466 289156 5468
rect 289212 5466 289236 5468
rect 289292 5466 289316 5468
rect 289372 5466 289386 5468
rect 289066 5414 289076 5466
rect 289132 5414 289142 5466
rect 288822 5412 288836 5414
rect 288892 5412 288916 5414
rect 288972 5412 288996 5414
rect 289052 5412 289076 5414
rect 289132 5412 289156 5414
rect 289212 5412 289236 5414
rect 289292 5412 289316 5414
rect 289372 5412 289386 5414
rect 288822 5392 289386 5412
rect 288822 4380 289386 4400
rect 288822 4378 288836 4380
rect 288892 4378 288916 4380
rect 288972 4378 288996 4380
rect 289052 4378 289076 4380
rect 289132 4378 289156 4380
rect 289212 4378 289236 4380
rect 289292 4378 289316 4380
rect 289372 4378 289386 4380
rect 289066 4326 289076 4378
rect 289132 4326 289142 4378
rect 288822 4324 288836 4326
rect 288892 4324 288916 4326
rect 288972 4324 288996 4326
rect 289052 4324 289076 4326
rect 289132 4324 289156 4326
rect 289212 4324 289236 4326
rect 289292 4324 289316 4326
rect 289372 4324 289386 4326
rect 288822 4304 289386 4324
rect 289464 4078 289492 5782
rect 289740 5778 289768 8092
rect 290844 6118 290872 8092
rect 290832 6112 290884 6118
rect 290832 6054 290884 6060
rect 289728 5772 289780 5778
rect 289728 5714 289780 5720
rect 291948 5710 291976 8092
rect 293144 6118 293172 8092
rect 292580 6112 292632 6118
rect 292580 6054 292632 6060
rect 293132 6112 293184 6118
rect 293132 6054 293184 6060
rect 292488 5772 292540 5778
rect 292488 5714 292540 5720
rect 291936 5704 291988 5710
rect 291936 5646 291988 5652
rect 290188 5636 290240 5642
rect 290188 5578 290240 5584
rect 289544 4140 289596 4146
rect 289544 4082 289596 4088
rect 288348 4072 288400 4078
rect 288348 4014 288400 4020
rect 289452 4072 289504 4078
rect 289452 4014 289504 4020
rect 288256 2916 288308 2922
rect 288256 2858 288308 2864
rect 288360 480 288388 4014
rect 288822 3292 289386 3312
rect 288822 3290 288836 3292
rect 288892 3290 288916 3292
rect 288972 3290 288996 3292
rect 289052 3290 289076 3292
rect 289132 3290 289156 3292
rect 289212 3290 289236 3292
rect 289292 3290 289316 3292
rect 289372 3290 289386 3292
rect 289066 3238 289076 3290
rect 289132 3238 289142 3290
rect 288822 3236 288836 3238
rect 288892 3236 288916 3238
rect 288972 3236 288996 3238
rect 289052 3236 289076 3238
rect 289132 3236 289156 3238
rect 289212 3236 289236 3238
rect 289292 3236 289316 3238
rect 289372 3236 289386 3238
rect 288822 3216 289386 3236
rect 288822 2204 289386 2224
rect 288822 2202 288836 2204
rect 288892 2202 288916 2204
rect 288972 2202 288996 2204
rect 289052 2202 289076 2204
rect 289132 2202 289156 2204
rect 289212 2202 289236 2204
rect 289292 2202 289316 2204
rect 289372 2202 289386 2204
rect 289066 2150 289076 2202
rect 289132 2150 289142 2202
rect 288822 2148 288836 2150
rect 288892 2148 288916 2150
rect 288972 2148 288996 2150
rect 289052 2148 289076 2150
rect 289132 2148 289156 2150
rect 289212 2148 289236 2150
rect 289292 2148 289316 2150
rect 289372 2148 289386 2150
rect 288822 2128 289386 2148
rect 289556 480 289584 4082
rect 290200 3534 290228 5578
rect 291384 5568 291436 5574
rect 291384 5510 291436 5516
rect 290188 3528 290240 3534
rect 290188 3470 290240 3476
rect 291396 3398 291424 5510
rect 291936 4072 291988 4078
rect 291936 4014 291988 4020
rect 291384 3392 291436 3398
rect 291384 3334 291436 3340
rect 290740 2916 290792 2922
rect 290740 2858 290792 2864
rect 290752 480 290780 2858
rect 291948 480 291976 4014
rect 292500 3602 292528 5714
rect 292592 3738 292620 6054
rect 294248 5574 294276 8092
rect 295352 5846 295380 8092
rect 295432 6112 295484 6118
rect 295432 6054 295484 6060
rect 295340 5840 295392 5846
rect 295340 5782 295392 5788
rect 294328 5704 294380 5710
rect 294328 5646 294380 5652
rect 294236 5568 294288 5574
rect 294236 5510 294288 5516
rect 294340 4078 294368 5646
rect 295444 4146 295472 6054
rect 296548 5710 296576 8092
rect 296536 5704 296588 5710
rect 296536 5646 296588 5652
rect 297652 5642 297680 8092
rect 297640 5636 297692 5642
rect 297640 5578 297692 5584
rect 298756 5574 298784 8092
rect 298928 5840 298980 5846
rect 298928 5782 298980 5788
rect 297824 5568 297876 5574
rect 297824 5510 297876 5516
rect 298744 5568 298796 5574
rect 298744 5510 298796 5516
rect 295432 4140 295484 4146
rect 295432 4082 295484 4088
rect 294328 4072 294380 4078
rect 294328 4014 294380 4020
rect 292580 3732 292632 3738
rect 292580 3674 292632 3680
rect 296720 3732 296772 3738
rect 296720 3674 296772 3680
rect 292488 3596 292540 3602
rect 292488 3538 292540 3544
rect 295524 3596 295576 3602
rect 295524 3538 295576 3544
rect 293132 3528 293184 3534
rect 293132 3470 293184 3476
rect 293144 480 293172 3470
rect 294328 3392 294380 3398
rect 294328 3334 294380 3340
rect 294340 480 294368 3334
rect 295536 480 295564 3538
rect 296732 480 296760 3674
rect 297836 2922 297864 5510
rect 297916 4072 297968 4078
rect 297916 4014 297968 4020
rect 297824 2916 297876 2922
rect 297824 2858 297876 2864
rect 297928 480 297956 4014
rect 298940 3058 298968 5782
rect 299952 5710 299980 8092
rect 301056 5846 301084 8092
rect 302160 6118 302188 8092
rect 302148 6112 302200 6118
rect 302148 6054 302200 6060
rect 301044 5840 301096 5846
rect 301044 5782 301096 5788
rect 303356 5710 303384 8092
rect 304264 6112 304316 6118
rect 304264 6054 304316 6060
rect 303712 5840 303764 5846
rect 303712 5782 303764 5788
rect 299204 5704 299256 5710
rect 299204 5646 299256 5652
rect 299940 5704 299992 5710
rect 299940 5646 299992 5652
rect 303068 5704 303120 5710
rect 303068 5646 303120 5652
rect 303344 5704 303396 5710
rect 303344 5646 303396 5652
rect 299112 4140 299164 4146
rect 299112 4082 299164 4088
rect 298928 3052 298980 3058
rect 298928 2994 298980 3000
rect 299124 480 299152 4082
rect 299216 3466 299244 5646
rect 300676 5636 300728 5642
rect 300676 5578 300728 5584
rect 300688 3534 300716 5578
rect 301780 5568 301832 5574
rect 301780 5510 301832 5516
rect 300676 3528 300728 3534
rect 300676 3470 300728 3476
rect 299204 3460 299256 3466
rect 299204 3402 299256 3408
rect 301792 3398 301820 5510
rect 303080 3466 303108 5646
rect 303724 4146 303752 5782
rect 303712 4140 303764 4146
rect 303712 4082 303764 4088
rect 304276 4010 304304 6054
rect 304460 5846 304488 8092
rect 304448 5840 304500 5846
rect 304448 5782 304500 5788
rect 305564 5710 305592 8092
rect 305000 5704 305052 5710
rect 305000 5646 305052 5652
rect 305552 5704 305604 5710
rect 305552 5646 305604 5652
rect 304264 4004 304316 4010
rect 304264 3946 304316 3952
rect 305012 3602 305040 5646
rect 306760 5574 306788 8092
rect 306822 6012 307386 6032
rect 306822 6010 306836 6012
rect 306892 6010 306916 6012
rect 306972 6010 306996 6012
rect 307052 6010 307076 6012
rect 307132 6010 307156 6012
rect 307212 6010 307236 6012
rect 307292 6010 307316 6012
rect 307372 6010 307386 6012
rect 307066 5958 307076 6010
rect 307132 5958 307142 6010
rect 306822 5956 306836 5958
rect 306892 5956 306916 5958
rect 306972 5956 306996 5958
rect 307052 5956 307076 5958
rect 307132 5956 307156 5958
rect 307212 5956 307236 5958
rect 307292 5956 307316 5958
rect 307372 5956 307386 5958
rect 306822 5936 307386 5956
rect 307668 5840 307720 5846
rect 307668 5782 307720 5788
rect 306748 5568 306800 5574
rect 306748 5510 306800 5516
rect 306822 4924 307386 4944
rect 306822 4922 306836 4924
rect 306892 4922 306916 4924
rect 306972 4922 306996 4924
rect 307052 4922 307076 4924
rect 307132 4922 307156 4924
rect 307212 4922 307236 4924
rect 307292 4922 307316 4924
rect 307372 4922 307386 4924
rect 307066 4870 307076 4922
rect 307132 4870 307142 4922
rect 306822 4868 306836 4870
rect 306892 4868 306916 4870
rect 306972 4868 306996 4870
rect 307052 4868 307076 4870
rect 307132 4868 307156 4870
rect 307212 4868 307236 4870
rect 307292 4868 307316 4870
rect 307372 4868 307386 4870
rect 306822 4848 307386 4868
rect 307484 4140 307536 4146
rect 307484 4082 307536 4088
rect 306822 3836 307386 3856
rect 306822 3834 306836 3836
rect 306892 3834 306916 3836
rect 306972 3834 306996 3836
rect 307052 3834 307076 3836
rect 307132 3834 307156 3836
rect 307212 3834 307236 3836
rect 307292 3834 307316 3836
rect 307372 3834 307386 3836
rect 307066 3782 307076 3834
rect 307132 3782 307142 3834
rect 306822 3780 306836 3782
rect 306892 3780 306916 3782
rect 306972 3780 306996 3782
rect 307052 3780 307076 3782
rect 307132 3780 307156 3782
rect 307212 3780 307236 3782
rect 307292 3780 307316 3782
rect 307372 3780 307386 3782
rect 306822 3760 307386 3780
rect 305000 3596 305052 3602
rect 305000 3538 305052 3544
rect 303804 3528 303856 3534
rect 303804 3470 303856 3476
rect 302608 3460 302660 3466
rect 302608 3402 302660 3408
rect 303068 3460 303120 3466
rect 303068 3402 303120 3408
rect 301780 3392 301832 3398
rect 301780 3334 301832 3340
rect 301412 3052 301464 3058
rect 301412 2994 301464 3000
rect 300308 2916 300360 2922
rect 300308 2858 300360 2864
rect 300320 480 300348 2858
rect 301424 480 301452 2994
rect 302620 480 302648 3402
rect 303816 480 303844 3470
rect 306196 3460 306248 3466
rect 306196 3402 306248 3408
rect 305000 3392 305052 3398
rect 305000 3334 305052 3340
rect 305012 480 305040 3334
rect 306208 480 306236 3402
rect 306822 2748 307386 2768
rect 306822 2746 306836 2748
rect 306892 2746 306916 2748
rect 306972 2746 306996 2748
rect 307052 2746 307076 2748
rect 307132 2746 307156 2748
rect 307212 2746 307236 2748
rect 307292 2746 307316 2748
rect 307372 2746 307386 2748
rect 307066 2694 307076 2746
rect 307132 2694 307142 2746
rect 306822 2692 306836 2694
rect 306892 2692 306916 2694
rect 306972 2692 306996 2694
rect 307052 2692 307076 2694
rect 307132 2692 307156 2694
rect 307212 2692 307236 2694
rect 307292 2692 307316 2694
rect 307372 2692 307386 2694
rect 306822 2672 307386 2692
rect 307496 2530 307524 4082
rect 307680 3194 307708 5782
rect 307864 5642 307892 8092
rect 308968 5778 308996 8092
rect 308956 5772 309008 5778
rect 308956 5714 309008 5720
rect 310164 5710 310192 8092
rect 308220 5704 308272 5710
rect 308220 5646 308272 5652
rect 310152 5704 310204 5710
rect 310152 5646 310204 5652
rect 307852 5636 307904 5642
rect 307852 5578 307904 5584
rect 307668 3188 307720 3194
rect 307668 3130 307720 3136
rect 308232 2854 308260 5646
rect 311164 5636 311216 5642
rect 311164 5578 311216 5584
rect 309968 5568 310020 5574
rect 309968 5510 310020 5516
rect 308588 4004 308640 4010
rect 308588 3946 308640 3952
rect 308220 2848 308272 2854
rect 308220 2790 308272 2796
rect 307404 2502 307524 2530
rect 307404 480 307432 2502
rect 308600 480 308628 3946
rect 309784 3596 309836 3602
rect 309784 3538 309836 3544
rect 309796 480 309824 3538
rect 309980 3466 310008 5510
rect 311176 3534 311204 5578
rect 311268 5574 311296 8092
rect 311808 5772 311860 5778
rect 311808 5714 311860 5720
rect 311256 5568 311308 5574
rect 311256 5510 311308 5516
rect 311820 3602 311848 5714
rect 312372 5642 312400 8092
rect 313096 5704 313148 5710
rect 313096 5646 313148 5652
rect 312360 5636 312412 5642
rect 312360 5578 312412 5584
rect 313108 4078 313136 5646
rect 313476 5574 313504 8092
rect 314672 6118 314700 8092
rect 314660 6112 314712 6118
rect 314660 6054 314712 6060
rect 315776 5914 315804 8092
rect 315764 5908 315816 5914
rect 315764 5850 315816 5856
rect 316880 5642 316908 8092
rect 318076 5710 318104 8092
rect 319180 6390 319208 8092
rect 319168 6384 319220 6390
rect 319168 6326 319220 6332
rect 318248 6112 318300 6118
rect 318248 6054 318300 6060
rect 318064 5704 318116 5710
rect 318064 5646 318116 5652
rect 314660 5636 314712 5642
rect 314660 5578 314712 5584
rect 316868 5636 316920 5642
rect 316868 5578 316920 5584
rect 313372 5568 313424 5574
rect 313372 5510 313424 5516
rect 313464 5568 313516 5574
rect 313464 5510 313516 5516
rect 313384 4146 313412 5510
rect 313372 4140 313424 4146
rect 313372 4082 313424 4088
rect 313096 4072 313148 4078
rect 313096 4014 313148 4020
rect 311808 3596 311860 3602
rect 311808 3538 311860 3544
rect 311164 3528 311216 3534
rect 311164 3470 311216 3476
rect 314568 3528 314620 3534
rect 314568 3470 314620 3476
rect 309968 3460 310020 3466
rect 309968 3402 310020 3408
rect 313372 3460 313424 3466
rect 313372 3402 313424 3408
rect 310980 3188 311032 3194
rect 310980 3130 311032 3136
rect 310992 480 311020 3130
rect 312176 2848 312228 2854
rect 312176 2790 312228 2796
rect 312188 480 312216 2790
rect 313384 480 313412 3402
rect 314580 480 314608 3470
rect 314672 3466 314700 5578
rect 317236 5568 317288 5574
rect 317236 5510 317288 5516
rect 316960 4072 317012 4078
rect 316960 4014 317012 4020
rect 315764 3596 315816 3602
rect 315764 3538 315816 3544
rect 314660 3460 314712 3466
rect 314660 3402 314712 3408
rect 315776 480 315804 3538
rect 316972 480 317000 4014
rect 317248 3194 317276 5510
rect 318064 4140 318116 4146
rect 318064 4082 318116 4088
rect 317236 3188 317288 3194
rect 317236 3130 317288 3136
rect 318076 480 318104 4082
rect 318260 3126 318288 6054
rect 318708 5908 318760 5914
rect 318708 5850 318760 5856
rect 318248 3120 318300 3126
rect 318248 3062 318300 3068
rect 318720 3058 318748 5850
rect 320088 5636 320140 5642
rect 320088 5578 320140 5584
rect 320100 3466 320128 5578
rect 320284 5574 320312 8092
rect 321480 5846 321508 8092
rect 322480 6384 322532 6390
rect 322480 6326 322532 6332
rect 321468 5840 321520 5846
rect 321468 5782 321520 5788
rect 321468 5704 321520 5710
rect 321468 5646 321520 5652
rect 320272 5568 320324 5574
rect 320272 5510 320324 5516
rect 319260 3460 319312 3466
rect 319260 3402 319312 3408
rect 320088 3460 320140 3466
rect 320088 3402 320140 3408
rect 318708 3052 318760 3058
rect 318708 2994 318760 3000
rect 319272 480 319300 3402
rect 321480 3398 321508 5646
rect 322492 4146 322520 6326
rect 322584 5914 322612 8092
rect 322572 5908 322624 5914
rect 322572 5850 322624 5856
rect 323584 5840 323636 5846
rect 323584 5782 323636 5788
rect 323032 5568 323084 5574
rect 323032 5510 323084 5516
rect 322480 4140 322532 4146
rect 322480 4082 322532 4088
rect 323044 4010 323072 5510
rect 323032 4004 323084 4010
rect 323032 3946 323084 3952
rect 323596 3534 323624 5782
rect 323688 5778 323716 8092
rect 324884 5914 324912 8092
rect 324320 5908 324372 5914
rect 324320 5850 324372 5856
rect 324872 5908 324924 5914
rect 324872 5850 324924 5856
rect 323676 5772 323728 5778
rect 323676 5714 323728 5720
rect 324332 3602 324360 5850
rect 325988 5574 326016 8092
rect 326988 5772 327040 5778
rect 326988 5714 327040 5720
rect 325976 5568 326028 5574
rect 325976 5510 326028 5516
rect 324822 5468 325386 5488
rect 324822 5466 324836 5468
rect 324892 5466 324916 5468
rect 324972 5466 324996 5468
rect 325052 5466 325076 5468
rect 325132 5466 325156 5468
rect 325212 5466 325236 5468
rect 325292 5466 325316 5468
rect 325372 5466 325386 5468
rect 325066 5414 325076 5466
rect 325132 5414 325142 5466
rect 324822 5412 324836 5414
rect 324892 5412 324916 5414
rect 324972 5412 324996 5414
rect 325052 5412 325076 5414
rect 325132 5412 325156 5414
rect 325212 5412 325236 5414
rect 325292 5412 325316 5414
rect 325372 5412 325386 5414
rect 324822 5392 325386 5412
rect 324822 4380 325386 4400
rect 324822 4378 324836 4380
rect 324892 4378 324916 4380
rect 324972 4378 324996 4380
rect 325052 4378 325076 4380
rect 325132 4378 325156 4380
rect 325212 4378 325236 4380
rect 325292 4378 325316 4380
rect 325372 4378 325386 4380
rect 325066 4326 325076 4378
rect 325132 4326 325142 4378
rect 324822 4324 324836 4326
rect 324892 4324 324916 4326
rect 324972 4324 324996 4326
rect 325052 4324 325076 4326
rect 325132 4324 325156 4326
rect 325212 4324 325236 4326
rect 325292 4324 325316 4326
rect 325372 4324 325386 4326
rect 324822 4304 325386 4324
rect 326436 4140 326488 4146
rect 326436 4082 326488 4088
rect 324320 3596 324372 3602
rect 324320 3538 324372 3544
rect 323584 3528 323636 3534
rect 323584 3470 323636 3476
rect 324044 3460 324096 3466
rect 324044 3402 324096 3408
rect 321468 3392 321520 3398
rect 321468 3334 321520 3340
rect 320456 3188 320508 3194
rect 320456 3130 320508 3136
rect 320468 480 320496 3130
rect 321652 3120 321704 3126
rect 321652 3062 321704 3068
rect 321664 480 321692 3062
rect 322848 3052 322900 3058
rect 322848 2994 322900 3000
rect 322860 480 322888 2994
rect 324056 480 324084 3402
rect 325424 3392 325476 3398
rect 325424 3334 325476 3340
rect 324822 3292 325386 3312
rect 324822 3290 324836 3292
rect 324892 3290 324916 3292
rect 324972 3290 324996 3292
rect 325052 3290 325076 3292
rect 325132 3290 325156 3292
rect 325212 3290 325236 3292
rect 325292 3290 325316 3292
rect 325372 3290 325386 3292
rect 325066 3238 325076 3290
rect 325132 3238 325142 3290
rect 324822 3236 324836 3238
rect 324892 3236 324916 3238
rect 324972 3236 324996 3238
rect 325052 3236 325076 3238
rect 325132 3236 325156 3238
rect 325212 3236 325236 3238
rect 325292 3236 325316 3238
rect 325372 3236 325386 3238
rect 324822 3216 325386 3236
rect 324822 2204 325386 2224
rect 324822 2202 324836 2204
rect 324892 2202 324916 2204
rect 324972 2202 324996 2204
rect 325052 2202 325076 2204
rect 325132 2202 325156 2204
rect 325212 2202 325236 2204
rect 325292 2202 325316 2204
rect 325372 2202 325386 2204
rect 325066 2150 325076 2202
rect 325132 2150 325142 2202
rect 324822 2148 324836 2150
rect 324892 2148 324916 2150
rect 324972 2148 324996 2150
rect 325052 2148 325076 2150
rect 325132 2148 325156 2150
rect 325212 2148 325236 2150
rect 325292 2148 325316 2150
rect 325372 2148 325386 2150
rect 324822 2128 325386 2148
rect 325436 1986 325464 3334
rect 325252 1958 325464 1986
rect 325252 480 325280 1958
rect 326448 480 326476 4082
rect 327000 3194 327028 5714
rect 327092 5642 327120 8092
rect 328288 6390 328316 8092
rect 328276 6384 328328 6390
rect 328276 6326 328328 6332
rect 328276 5908 328328 5914
rect 328276 5850 328328 5856
rect 327080 5636 327132 5642
rect 327080 5578 327132 5584
rect 327632 4004 327684 4010
rect 327632 3946 327684 3952
rect 326988 3188 327040 3194
rect 326988 3130 327040 3136
rect 327644 480 327672 3946
rect 328288 3058 328316 5850
rect 329392 5710 329420 8092
rect 330496 5846 330524 8092
rect 331692 6662 331720 8092
rect 331680 6656 331732 6662
rect 331680 6598 331732 6604
rect 330576 6384 330628 6390
rect 330576 6326 330628 6332
rect 330484 5840 330536 5846
rect 330484 5782 330536 5788
rect 329380 5704 329432 5710
rect 329380 5646 329432 5652
rect 329748 5568 329800 5574
rect 329748 5510 329800 5516
rect 329760 3534 329788 5510
rect 330024 3596 330076 3602
rect 330024 3538 330076 3544
rect 328828 3528 328880 3534
rect 328828 3470 328880 3476
rect 329748 3528 329800 3534
rect 329748 3470 329800 3476
rect 328276 3052 328328 3058
rect 328276 2994 328328 3000
rect 328840 480 328868 3470
rect 330036 480 330064 3538
rect 330588 3126 330616 6326
rect 332796 6118 332824 8092
rect 332784 6112 332836 6118
rect 332784 6054 332836 6060
rect 332968 5840 333020 5846
rect 332968 5782 333020 5788
rect 332416 5704 332468 5710
rect 332416 5646 332468 5652
rect 330852 5636 330904 5642
rect 330852 5578 330904 5584
rect 330864 3466 330892 5578
rect 332428 4078 332456 5646
rect 332416 4072 332468 4078
rect 332416 4014 332468 4020
rect 332980 3670 333008 5782
rect 333900 5642 333928 8092
rect 333980 6656 334032 6662
rect 333980 6598 334032 6604
rect 333888 5636 333940 5642
rect 333888 5578 333940 5584
rect 332968 3664 333020 3670
rect 332968 3606 333020 3612
rect 333992 3602 334020 6598
rect 335096 5914 335124 8092
rect 335084 5908 335136 5914
rect 335084 5850 335136 5856
rect 336200 5574 336228 8092
rect 337304 6254 337332 8092
rect 337292 6248 337344 6254
rect 337292 6190 337344 6196
rect 336280 6112 336332 6118
rect 336280 6054 336332 6060
rect 336188 5568 336240 5574
rect 336188 5510 336240 5516
rect 336292 4010 336320 6054
rect 337384 5908 337436 5914
rect 337384 5850 337436 5856
rect 336648 5636 336700 5642
rect 336648 5578 336700 5584
rect 336280 4004 336332 4010
rect 336280 3946 336332 3952
rect 333980 3596 334032 3602
rect 333980 3538 334032 3544
rect 333612 3528 333664 3534
rect 333612 3470 333664 3476
rect 330852 3460 330904 3466
rect 330852 3402 330904 3408
rect 331220 3188 331272 3194
rect 331220 3130 331272 3136
rect 330576 3120 330628 3126
rect 330576 3062 330628 3068
rect 331232 480 331260 3130
rect 332416 3052 332468 3058
rect 332416 2994 332468 3000
rect 332428 480 332456 2994
rect 333624 480 333652 3470
rect 334716 3460 334768 3466
rect 334716 3402 334768 3408
rect 334728 480 334756 3402
rect 336660 3194 336688 5578
rect 337108 4072 337160 4078
rect 337108 4014 337160 4020
rect 336648 3188 336700 3194
rect 336648 3130 336700 3136
rect 335912 3120 335964 3126
rect 335912 3062 335964 3068
rect 335924 480 335952 3062
rect 337120 480 337148 4014
rect 337396 2990 337424 5850
rect 338500 5710 338528 8092
rect 338488 5704 338540 5710
rect 338488 5646 338540 5652
rect 339604 5574 339632 8092
rect 340708 6390 340736 8092
rect 340696 6384 340748 6390
rect 340696 6326 340748 6332
rect 339684 6248 339736 6254
rect 339684 6190 339736 6196
rect 339408 5568 339460 5574
rect 339408 5510 339460 5516
rect 339592 5568 339644 5574
rect 339592 5510 339644 5516
rect 338304 3664 338356 3670
rect 338304 3606 338356 3612
rect 337384 2984 337436 2990
rect 337384 2926 337436 2932
rect 338316 480 338344 3606
rect 339420 3534 339448 5510
rect 339500 3596 339552 3602
rect 339500 3538 339552 3544
rect 339408 3528 339460 3534
rect 339408 3470 339460 3476
rect 339512 480 339540 3538
rect 339696 3126 339724 6190
rect 341904 5710 341932 8092
rect 342720 6384 342772 6390
rect 342720 6326 342772 6332
rect 341800 5704 341852 5710
rect 341800 5646 341852 5652
rect 341892 5704 341944 5710
rect 341892 5646 341944 5652
rect 341812 4078 341840 5646
rect 342260 5568 342312 5574
rect 342260 5510 342312 5516
rect 341800 4072 341852 4078
rect 341800 4014 341852 4020
rect 340696 4004 340748 4010
rect 340696 3946 340748 3952
rect 339684 3120 339736 3126
rect 339684 3062 339736 3068
rect 340708 480 340736 3946
rect 342272 3670 342300 5510
rect 342732 3942 342760 6326
rect 343008 6186 343036 8092
rect 342996 6180 343048 6186
rect 342996 6122 343048 6128
rect 342822 6012 343386 6032
rect 342822 6010 342836 6012
rect 342892 6010 342916 6012
rect 342972 6010 342996 6012
rect 343052 6010 343076 6012
rect 343132 6010 343156 6012
rect 343212 6010 343236 6012
rect 343292 6010 343316 6012
rect 343372 6010 343386 6012
rect 343066 5958 343076 6010
rect 343132 5958 343142 6010
rect 342822 5956 342836 5958
rect 342892 5956 342916 5958
rect 342972 5956 342996 5958
rect 343052 5956 343076 5958
rect 343132 5956 343156 5958
rect 343212 5956 343236 5958
rect 343292 5956 343316 5958
rect 343372 5956 343386 5958
rect 342822 5936 343386 5956
rect 344112 5846 344140 8092
rect 344100 5840 344152 5846
rect 344100 5782 344152 5788
rect 343640 5704 343692 5710
rect 343640 5646 343692 5652
rect 342822 4924 343386 4944
rect 342822 4922 342836 4924
rect 342892 4922 342916 4924
rect 342972 4922 342996 4924
rect 343052 4922 343076 4924
rect 343132 4922 343156 4924
rect 343212 4922 343236 4924
rect 343292 4922 343316 4924
rect 343372 4922 343386 4924
rect 343066 4870 343076 4922
rect 343132 4870 343142 4922
rect 342822 4868 342836 4870
rect 342892 4868 342916 4870
rect 342972 4868 342996 4870
rect 343052 4868 343076 4870
rect 343132 4868 343156 4870
rect 343212 4868 343236 4870
rect 343292 4868 343316 4870
rect 343372 4868 343386 4870
rect 342822 4848 343386 4868
rect 342720 3936 342772 3942
rect 342720 3878 342772 3884
rect 342822 3836 343386 3856
rect 342822 3834 342836 3836
rect 342892 3834 342916 3836
rect 342972 3834 342996 3836
rect 343052 3834 343076 3836
rect 343132 3834 343156 3836
rect 343212 3834 343236 3836
rect 343292 3834 343316 3836
rect 343372 3834 343386 3836
rect 343066 3782 343076 3834
rect 343132 3782 343142 3834
rect 342822 3780 342836 3782
rect 342892 3780 342916 3782
rect 342972 3780 342996 3782
rect 343052 3780 343076 3782
rect 343132 3780 343156 3782
rect 343212 3780 343236 3782
rect 343292 3780 343316 3782
rect 343372 3780 343386 3782
rect 342822 3760 343386 3780
rect 342260 3664 342312 3670
rect 342260 3606 342312 3612
rect 343652 3466 343680 5646
rect 345308 5642 345336 8092
rect 345940 6180 345992 6186
rect 345940 6122 345992 6128
rect 345296 5636 345348 5642
rect 345296 5578 345348 5584
rect 344284 3528 344336 3534
rect 344284 3470 344336 3476
rect 343640 3460 343692 3466
rect 343640 3402 343692 3408
rect 341892 3188 341944 3194
rect 341892 3130 341944 3136
rect 341904 480 341932 3130
rect 342720 2984 342772 2990
rect 342720 2926 342772 2932
rect 342732 2530 342760 2926
rect 342822 2748 343386 2768
rect 342822 2746 342836 2748
rect 342892 2746 342916 2748
rect 342972 2746 342996 2748
rect 343052 2746 343076 2748
rect 343132 2746 343156 2748
rect 343212 2746 343236 2748
rect 343292 2746 343316 2748
rect 343372 2746 343386 2748
rect 343066 2694 343076 2746
rect 343132 2694 343142 2746
rect 342822 2692 342836 2694
rect 342892 2692 342916 2694
rect 342972 2692 342996 2694
rect 343052 2692 343076 2694
rect 343132 2692 343156 2694
rect 343212 2692 343236 2694
rect 343292 2692 343316 2694
rect 343372 2692 343386 2694
rect 342822 2672 343386 2692
rect 342732 2502 343128 2530
rect 343100 480 343128 2502
rect 344296 480 344324 3470
rect 345952 3194 345980 6122
rect 346412 5574 346440 8092
rect 347516 6390 347544 8092
rect 347504 6384 347556 6390
rect 347504 6326 347556 6332
rect 348712 5846 348740 8092
rect 347412 5840 347464 5846
rect 347412 5782 347464 5788
rect 348700 5840 348752 5846
rect 348700 5782 348752 5788
rect 346400 5568 346452 5574
rect 346400 5510 346452 5516
rect 346676 4072 346728 4078
rect 346676 4014 346728 4020
rect 345940 3188 345992 3194
rect 345940 3130 345992 3136
rect 345480 3120 345532 3126
rect 345480 3062 345532 3068
rect 345492 480 345520 3062
rect 346688 480 346716 4014
rect 347424 3058 347452 5782
rect 349816 5710 349844 8092
rect 349804 5704 349856 5710
rect 349804 5646 349856 5652
rect 350920 5642 350948 8092
rect 351736 5840 351788 5846
rect 351736 5782 351788 5788
rect 348976 5636 349028 5642
rect 348976 5578 349028 5584
rect 350908 5636 350960 5642
rect 350908 5578 350960 5584
rect 347872 3664 347924 3670
rect 347872 3606 347924 3612
rect 347412 3052 347464 3058
rect 347412 2994 347464 3000
rect 347884 480 347912 3606
rect 348988 3398 349016 5578
rect 350356 5568 350408 5574
rect 350356 5510 350408 5516
rect 349068 3936 349120 3942
rect 349068 3878 349120 3884
rect 348976 3392 349028 3398
rect 348976 3334 349028 3340
rect 349080 480 349108 3878
rect 350368 3466 350396 5510
rect 351748 4146 351776 5782
rect 352024 5574 352052 8092
rect 353220 6322 353248 8092
rect 353208 6316 353260 6322
rect 353208 6258 353260 6264
rect 354324 6254 354352 8092
rect 354312 6248 354364 6254
rect 354312 6190 354364 6196
rect 355428 6186 355456 8092
rect 356624 6526 356652 8092
rect 356612 6520 356664 6526
rect 356612 6462 356664 6468
rect 356152 6384 356204 6390
rect 356152 6326 356204 6332
rect 355416 6180 355468 6186
rect 355416 6122 355468 6128
rect 352288 5704 352340 5710
rect 352288 5646 352340 5652
rect 352012 5568 352064 5574
rect 352012 5510 352064 5516
rect 351736 4140 351788 4146
rect 351736 4082 351788 4088
rect 352300 3602 352328 5646
rect 353300 5636 353352 5642
rect 353300 5578 353352 5584
rect 352288 3596 352340 3602
rect 352288 3538 352340 3544
rect 353312 3534 353340 5578
rect 355508 5568 355560 5574
rect 355508 5510 355560 5516
rect 353300 3528 353352 3534
rect 353300 3470 353352 3476
rect 350264 3460 350316 3466
rect 350264 3402 350316 3408
rect 350356 3460 350408 3466
rect 350356 3402 350408 3408
rect 354956 3460 355008 3466
rect 354956 3402 355008 3408
rect 350276 480 350304 3402
rect 353760 3392 353812 3398
rect 353760 3334 353812 3340
rect 351368 3188 351420 3194
rect 351368 3130 351420 3136
rect 351380 480 351408 3130
rect 352564 3052 352616 3058
rect 352564 2994 352616 3000
rect 352576 480 352604 2994
rect 353772 480 353800 3334
rect 354968 480 354996 3402
rect 355520 2854 355548 5510
rect 355508 2848 355560 2854
rect 355508 2790 355560 2796
rect 356164 480 356192 6326
rect 357728 5710 357756 8092
rect 357716 5704 357768 5710
rect 357716 5646 357768 5652
rect 358832 5574 358860 8092
rect 360028 6594 360056 8092
rect 360016 6588 360068 6594
rect 360016 6530 360068 6536
rect 361132 6390 361160 8092
rect 362236 6458 362264 8092
rect 362224 6452 362276 6458
rect 362224 6394 362276 6400
rect 361120 6384 361172 6390
rect 361120 6326 361172 6332
rect 362132 6316 362184 6322
rect 362132 6258 362184 6264
rect 360752 5704 360804 5710
rect 360752 5646 360804 5652
rect 358820 5568 358872 5574
rect 358820 5510 358872 5516
rect 357348 4140 357400 4146
rect 357348 4082 357400 4088
rect 357360 480 357388 4082
rect 360764 4078 360792 5646
rect 361580 5568 361632 5574
rect 361580 5510 361632 5516
rect 360822 5468 361386 5488
rect 360822 5466 360836 5468
rect 360892 5466 360916 5468
rect 360972 5466 360996 5468
rect 361052 5466 361076 5468
rect 361132 5466 361156 5468
rect 361212 5466 361236 5468
rect 361292 5466 361316 5468
rect 361372 5466 361386 5468
rect 361066 5414 361076 5466
rect 361132 5414 361142 5466
rect 360822 5412 360836 5414
rect 360892 5412 360916 5414
rect 360972 5412 360996 5414
rect 361052 5412 361076 5414
rect 361132 5412 361156 5414
rect 361212 5412 361236 5414
rect 361292 5412 361316 5414
rect 361372 5412 361386 5414
rect 360822 5392 361386 5412
rect 360822 4380 361386 4400
rect 360822 4378 360836 4380
rect 360892 4378 360916 4380
rect 360972 4378 360996 4380
rect 361052 4378 361076 4380
rect 361132 4378 361156 4380
rect 361212 4378 361236 4380
rect 361292 4378 361316 4380
rect 361372 4378 361386 4380
rect 361066 4326 361076 4378
rect 361132 4326 361142 4378
rect 360822 4324 360836 4326
rect 360892 4324 360916 4326
rect 360972 4324 360996 4326
rect 361052 4324 361076 4326
rect 361132 4324 361156 4326
rect 361212 4324 361236 4326
rect 361292 4324 361316 4326
rect 361372 4324 361386 4326
rect 360822 4304 361386 4324
rect 360752 4072 360804 4078
rect 360752 4014 360804 4020
rect 358544 3596 358596 3602
rect 358544 3538 358596 3544
rect 358556 480 358584 3538
rect 359740 3528 359792 3534
rect 359740 3470 359792 3476
rect 359752 480 359780 3470
rect 361592 3466 361620 5510
rect 361580 3460 361632 3466
rect 361580 3402 361632 3408
rect 360822 3292 361386 3312
rect 360822 3290 360836 3292
rect 360892 3290 360916 3292
rect 360972 3290 360996 3292
rect 361052 3290 361076 3292
rect 361132 3290 361156 3292
rect 361212 3290 361236 3292
rect 361292 3290 361316 3292
rect 361372 3290 361386 3292
rect 361066 3238 361076 3290
rect 361132 3238 361142 3290
rect 360822 3236 360836 3238
rect 360892 3236 360916 3238
rect 360972 3236 360996 3238
rect 361052 3236 361076 3238
rect 361132 3236 361156 3238
rect 361212 3236 361236 3238
rect 361292 3236 361316 3238
rect 361372 3236 361386 3238
rect 360822 3216 361386 3236
rect 360752 2848 360804 2854
rect 360752 2790 360804 2796
rect 360764 1986 360792 2790
rect 360822 2204 361386 2224
rect 360822 2202 360836 2204
rect 360892 2202 360916 2204
rect 360972 2202 360996 2204
rect 361052 2202 361076 2204
rect 361132 2202 361156 2204
rect 361212 2202 361236 2204
rect 361292 2202 361316 2204
rect 361372 2202 361386 2204
rect 361066 2150 361076 2202
rect 361132 2150 361142 2202
rect 360822 2148 360836 2150
rect 360892 2148 360916 2150
rect 360972 2148 360996 2150
rect 361052 2148 361076 2150
rect 361132 2148 361156 2150
rect 361212 2148 361236 2150
rect 361292 2148 361316 2150
rect 361372 2148 361386 2150
rect 360822 2128 361386 2148
rect 360764 1958 360976 1986
rect 360948 480 360976 1958
rect 362144 480 362172 6258
rect 363432 6254 363460 8092
rect 364536 6322 364564 8092
rect 364524 6316 364576 6322
rect 364524 6258 364576 6264
rect 363328 6248 363380 6254
rect 363328 6190 363380 6196
rect 363420 6248 363472 6254
rect 363420 6190 363472 6196
rect 363340 480 363368 6190
rect 364524 6180 364576 6186
rect 364524 6122 364576 6128
rect 364536 480 364564 6122
rect 365640 5642 365668 8092
rect 365720 6520 365772 6526
rect 365720 6462 365772 6468
rect 365628 5636 365680 5642
rect 365628 5578 365680 5584
rect 365732 480 365760 6462
rect 366836 5574 366864 8092
rect 367940 6322 367968 8092
rect 369044 6526 369072 8092
rect 370240 6594 370268 8092
rect 371344 6730 371372 8092
rect 371332 6724 371384 6730
rect 371332 6666 371384 6672
rect 369216 6588 369268 6594
rect 369216 6530 369268 6536
rect 370228 6588 370280 6594
rect 370228 6530 370280 6536
rect 369032 6520 369084 6526
rect 369032 6462 369084 6468
rect 367468 6316 367520 6322
rect 367468 6258 367520 6264
rect 367928 6316 367980 6322
rect 367928 6258 367980 6264
rect 367100 5636 367152 5642
rect 367100 5578 367152 5584
rect 366824 5568 366876 5574
rect 366824 5510 366876 5516
rect 366916 4072 366968 4078
rect 366916 4014 366968 4020
rect 366928 480 366956 4014
rect 367112 3194 367140 5578
rect 367480 3602 367508 6258
rect 368480 5568 368532 5574
rect 368480 5510 368532 5516
rect 367468 3596 367520 3602
rect 367468 3538 367520 3544
rect 368020 3460 368072 3466
rect 368020 3402 368072 3408
rect 367100 3188 367152 3194
rect 367100 3130 367152 3136
rect 368032 480 368060 3402
rect 368492 3398 368520 5510
rect 368480 3392 368532 3398
rect 368480 3334 368532 3340
rect 369228 480 369256 6530
rect 371608 6452 371660 6458
rect 371608 6394 371660 6400
rect 370412 6384 370464 6390
rect 370412 6326 370464 6332
rect 370424 480 370452 6326
rect 371620 480 371648 6394
rect 372448 6186 372476 8092
rect 373644 6798 373672 8092
rect 373632 6792 373684 6798
rect 373632 6734 373684 6740
rect 374748 6458 374776 8092
rect 374736 6452 374788 6458
rect 374736 6394 374788 6400
rect 375852 6254 375880 8092
rect 377048 6662 377076 8092
rect 378152 6866 378180 8092
rect 378140 6860 378192 6866
rect 378140 6802 378192 6808
rect 377036 6656 377088 6662
rect 377036 6598 377088 6604
rect 378692 6520 378744 6526
rect 378692 6462 378744 6468
rect 377588 6316 377640 6322
rect 377588 6258 377640 6264
rect 372804 6248 372856 6254
rect 372804 6190 372856 6196
rect 375840 6248 375892 6254
rect 375840 6190 375892 6196
rect 372436 6180 372488 6186
rect 372436 6122 372488 6128
rect 372816 480 372844 6190
rect 374000 3596 374052 3602
rect 374000 3538 374052 3544
rect 374012 480 374040 3538
rect 376392 3392 376444 3398
rect 376392 3334 376444 3340
rect 375196 3188 375248 3194
rect 375196 3130 375248 3136
rect 375208 480 375236 3130
rect 376404 480 376432 3334
rect 377600 480 377628 6258
rect 378704 2530 378732 6462
rect 379256 6390 379284 8092
rect 379980 6588 380032 6594
rect 379980 6530 380032 6536
rect 379244 6384 379296 6390
rect 379244 6326 379296 6332
rect 378822 6012 379386 6032
rect 378822 6010 378836 6012
rect 378892 6010 378916 6012
rect 378972 6010 378996 6012
rect 379052 6010 379076 6012
rect 379132 6010 379156 6012
rect 379212 6010 379236 6012
rect 379292 6010 379316 6012
rect 379372 6010 379386 6012
rect 379066 5958 379076 6010
rect 379132 5958 379142 6010
rect 378822 5956 378836 5958
rect 378892 5956 378916 5958
rect 378972 5956 378996 5958
rect 379052 5956 379076 5958
rect 379132 5956 379156 5958
rect 379212 5956 379236 5958
rect 379292 5956 379316 5958
rect 379372 5956 379386 5958
rect 378822 5936 379386 5956
rect 378822 4924 379386 4944
rect 378822 4922 378836 4924
rect 378892 4922 378916 4924
rect 378972 4922 378996 4924
rect 379052 4922 379076 4924
rect 379132 4922 379156 4924
rect 379212 4922 379236 4924
rect 379292 4922 379316 4924
rect 379372 4922 379386 4924
rect 379066 4870 379076 4922
rect 379132 4870 379142 4922
rect 378822 4868 378836 4870
rect 378892 4868 378916 4870
rect 378972 4868 378996 4870
rect 379052 4868 379076 4870
rect 379132 4868 379156 4870
rect 379212 4868 379236 4870
rect 379292 4868 379316 4870
rect 379372 4868 379386 4870
rect 378822 4848 379386 4868
rect 378822 3836 379386 3856
rect 378822 3834 378836 3836
rect 378892 3834 378916 3836
rect 378972 3834 378996 3836
rect 379052 3834 379076 3836
rect 379132 3834 379156 3836
rect 379212 3834 379236 3836
rect 379292 3834 379316 3836
rect 379372 3834 379386 3836
rect 379066 3782 379076 3834
rect 379132 3782 379142 3834
rect 378822 3780 378836 3782
rect 378892 3780 378916 3782
rect 378972 3780 378996 3782
rect 379052 3780 379076 3782
rect 379132 3780 379156 3782
rect 379212 3780 379236 3782
rect 379292 3780 379316 3782
rect 379372 3780 379386 3782
rect 378822 3760 379386 3780
rect 378822 2748 379386 2768
rect 378822 2746 378836 2748
rect 378892 2746 378916 2748
rect 378972 2746 378996 2748
rect 379052 2746 379076 2748
rect 379132 2746 379156 2748
rect 379212 2746 379236 2748
rect 379292 2746 379316 2748
rect 379372 2746 379386 2748
rect 379066 2694 379076 2746
rect 379132 2694 379142 2746
rect 378822 2692 378836 2694
rect 378892 2692 378916 2694
rect 378972 2692 378996 2694
rect 379052 2692 379076 2694
rect 379132 2692 379156 2694
rect 379212 2692 379236 2694
rect 379292 2692 379316 2694
rect 379372 2692 379386 2694
rect 378822 2672 379386 2692
rect 378704 2502 378824 2530
rect 378796 480 378824 2502
rect 379992 480 380020 6530
rect 380452 5846 380480 8092
rect 381176 6724 381228 6730
rect 381176 6666 381228 6672
rect 380440 5840 380492 5846
rect 380440 5782 380492 5788
rect 381188 480 381216 6666
rect 381556 5710 381584 8092
rect 382660 6526 382688 8092
rect 383856 6798 383884 8092
rect 383568 6792 383620 6798
rect 383568 6734 383620 6740
rect 383844 6792 383896 6798
rect 383844 6734 383896 6740
rect 382648 6520 382700 6526
rect 382648 6462 382700 6468
rect 382372 6180 382424 6186
rect 382372 6122 382424 6128
rect 382280 5840 382332 5846
rect 382280 5782 382332 5788
rect 381544 5704 381596 5710
rect 381544 5646 381596 5652
rect 382292 3466 382320 5782
rect 382280 3460 382332 3466
rect 382280 3402 382332 3408
rect 382384 480 382412 6122
rect 383580 480 383608 6734
rect 384960 6730 384988 8092
rect 384948 6724 385000 6730
rect 384948 6666 385000 6672
rect 384672 6452 384724 6458
rect 384672 6394 384724 6400
rect 384684 480 384712 6394
rect 386064 6322 386092 8092
rect 387064 6656 387116 6662
rect 387064 6598 387116 6604
rect 386052 6316 386104 6322
rect 386052 6258 386104 6264
rect 385868 6248 385920 6254
rect 385868 6190 385920 6196
rect 384948 5704 385000 5710
rect 384948 5646 385000 5652
rect 384960 2922 384988 5646
rect 384948 2916 385000 2922
rect 384948 2858 385000 2864
rect 385880 480 385908 6190
rect 387076 480 387104 6598
rect 387260 6458 387288 8092
rect 388260 6860 388312 6866
rect 388260 6802 388312 6808
rect 387248 6452 387300 6458
rect 387248 6394 387300 6400
rect 388272 480 388300 6802
rect 388364 6254 388392 8092
rect 389088 6384 389140 6390
rect 389088 6326 389140 6332
rect 388352 6248 388404 6254
rect 388352 6190 388404 6196
rect 389100 3210 389128 6326
rect 389468 6186 389496 8092
rect 390572 6730 390600 8092
rect 390560 6724 390612 6730
rect 390560 6666 390612 6672
rect 391768 6390 391796 8092
rect 392872 6526 392900 8092
rect 392768 6520 392820 6526
rect 392768 6462 392820 6468
rect 392860 6520 392912 6526
rect 392860 6462 392912 6468
rect 391756 6384 391808 6390
rect 391756 6326 391808 6332
rect 392780 6338 392808 6462
rect 392780 6310 393084 6338
rect 389456 6180 389508 6186
rect 389456 6122 389508 6128
rect 390652 3460 390704 3466
rect 390652 3402 390704 3408
rect 389100 3182 389496 3210
rect 389468 480 389496 3182
rect 390664 480 390692 3402
rect 391848 2916 391900 2922
rect 391848 2858 391900 2864
rect 391860 480 391888 2858
rect 393056 480 393084 6310
rect 393976 6118 394004 8092
rect 394240 6792 394292 6798
rect 394240 6734 394292 6740
rect 394056 6656 394108 6662
rect 394056 6598 394108 6604
rect 393964 6112 394016 6118
rect 393964 6054 394016 6060
rect 394068 3398 394096 6598
rect 394056 3392 394108 3398
rect 394056 3334 394108 3340
rect 394252 480 394280 6734
rect 395172 5574 395200 8092
rect 396276 6662 396304 8092
rect 396264 6656 396316 6662
rect 396264 6598 396316 6604
rect 397380 6322 397408 8092
rect 398576 6458 398604 8092
rect 399680 6866 399708 8092
rect 399668 6860 399720 6866
rect 399668 6802 399720 6808
rect 400784 6798 400812 8092
rect 400772 6792 400824 6798
rect 400772 6734 400824 6740
rect 401324 6724 401376 6730
rect 401324 6666 401376 6672
rect 397828 6452 397880 6458
rect 397828 6394 397880 6400
rect 398564 6452 398616 6458
rect 398564 6394 398616 6400
rect 396632 6316 396684 6322
rect 396632 6258 396684 6264
rect 397368 6316 397420 6322
rect 397368 6258 397420 6264
rect 395160 5568 395212 5574
rect 395160 5510 395212 5516
rect 395436 3392 395488 3398
rect 395436 3334 395488 3340
rect 395448 480 395476 3334
rect 396644 480 396672 6258
rect 396822 5468 397386 5488
rect 396822 5466 396836 5468
rect 396892 5466 396916 5468
rect 396972 5466 396996 5468
rect 397052 5466 397076 5468
rect 397132 5466 397156 5468
rect 397212 5466 397236 5468
rect 397292 5466 397316 5468
rect 397372 5466 397386 5468
rect 397066 5414 397076 5466
rect 397132 5414 397142 5466
rect 396822 5412 396836 5414
rect 396892 5412 396916 5414
rect 396972 5412 396996 5414
rect 397052 5412 397076 5414
rect 397132 5412 397156 5414
rect 397212 5412 397236 5414
rect 397292 5412 397316 5414
rect 397372 5412 397386 5414
rect 396822 5392 397386 5412
rect 396822 4380 397386 4400
rect 396822 4378 396836 4380
rect 396892 4378 396916 4380
rect 396972 4378 396996 4380
rect 397052 4378 397076 4380
rect 397132 4378 397156 4380
rect 397212 4378 397236 4380
rect 397292 4378 397316 4380
rect 397372 4378 397386 4380
rect 397066 4326 397076 4378
rect 397132 4326 397142 4378
rect 396822 4324 396836 4326
rect 396892 4324 396916 4326
rect 396972 4324 396996 4326
rect 397052 4324 397076 4326
rect 397132 4324 397156 4326
rect 397212 4324 397236 4326
rect 397292 4324 397316 4326
rect 397372 4324 397386 4326
rect 396822 4304 397386 4324
rect 396822 3292 397386 3312
rect 396822 3290 396836 3292
rect 396892 3290 396916 3292
rect 396972 3290 396996 3292
rect 397052 3290 397076 3292
rect 397132 3290 397156 3292
rect 397212 3290 397236 3292
rect 397292 3290 397316 3292
rect 397372 3290 397386 3292
rect 397066 3238 397076 3290
rect 397132 3238 397142 3290
rect 396822 3236 396836 3238
rect 396892 3236 396916 3238
rect 396972 3236 396996 3238
rect 397052 3236 397076 3238
rect 397132 3236 397156 3238
rect 397212 3236 397236 3238
rect 397292 3236 397316 3238
rect 397372 3236 397386 3238
rect 396822 3216 397386 3236
rect 396822 2204 397386 2224
rect 396822 2202 396836 2204
rect 396892 2202 396916 2204
rect 396972 2202 396996 2204
rect 397052 2202 397076 2204
rect 397132 2202 397156 2204
rect 397212 2202 397236 2204
rect 397292 2202 397316 2204
rect 397372 2202 397386 2204
rect 397066 2150 397076 2202
rect 397132 2150 397142 2202
rect 396822 2148 396836 2150
rect 396892 2148 396916 2150
rect 396972 2148 396996 2150
rect 397052 2148 397076 2150
rect 397132 2148 397156 2150
rect 397212 2148 397236 2150
rect 397292 2148 397316 2150
rect 397372 2148 397386 2150
rect 396822 2128 397386 2148
rect 397840 480 397868 6394
rect 399024 6248 399076 6254
rect 399024 6190 399076 6196
rect 398656 5568 398708 5574
rect 398656 5510 398708 5516
rect 398668 3466 398696 5510
rect 398656 3460 398708 3466
rect 398656 3402 398708 3408
rect 399036 480 399064 6190
rect 400220 6180 400272 6186
rect 400220 6122 400272 6128
rect 400232 480 400260 6122
rect 401336 480 401364 6666
rect 401980 6594 402008 8092
rect 403084 6730 403112 8092
rect 403072 6724 403124 6730
rect 403072 6666 403124 6672
rect 401968 6588 402020 6594
rect 401968 6530 402020 6536
rect 403716 6520 403768 6526
rect 403716 6462 403768 6468
rect 402520 6384 402572 6390
rect 402520 6326 402572 6332
rect 402532 480 402560 6326
rect 403728 480 403756 6462
rect 404188 6254 404216 8092
rect 404176 6248 404228 6254
rect 404176 6190 404228 6196
rect 405384 6186 405412 8092
rect 406488 6390 406516 8092
rect 407304 6656 407356 6662
rect 407304 6598 407356 6604
rect 406476 6384 406528 6390
rect 406476 6326 406528 6332
rect 405372 6180 405424 6186
rect 405372 6122 405424 6128
rect 403808 6112 403860 6118
rect 403808 6054 403860 6060
rect 403820 3058 403848 6054
rect 406108 3460 406160 3466
rect 406108 3402 406160 3408
rect 403808 3052 403860 3058
rect 403808 2994 403860 3000
rect 404912 3052 404964 3058
rect 404912 2994 404964 3000
rect 404924 480 404952 2994
rect 406120 480 406148 3402
rect 407316 480 407344 6598
rect 407592 6526 407620 8092
rect 408500 6860 408552 6866
rect 408500 6802 408552 6808
rect 407580 6520 407632 6526
rect 407580 6462 407632 6468
rect 408408 6316 408460 6322
rect 408408 6258 408460 6264
rect 408420 4026 408448 6258
rect 408512 4146 408540 6802
rect 408788 5914 408816 8092
rect 409696 6452 409748 6458
rect 409696 6394 409748 6400
rect 408776 5908 408828 5914
rect 408776 5850 408828 5856
rect 408500 4140 408552 4146
rect 408500 4082 408552 4088
rect 408420 3998 408540 4026
rect 408512 480 408540 3998
rect 409708 480 409736 6394
rect 409892 5710 409920 8092
rect 410996 5778 411024 8092
rect 412088 6792 412140 6798
rect 412088 6734 412140 6740
rect 410984 5772 411036 5778
rect 410984 5714 411036 5720
rect 409880 5704 409932 5710
rect 409880 5646 409932 5652
rect 410892 4140 410944 4146
rect 410892 4082 410944 4088
rect 410904 480 410932 4082
rect 412100 480 412128 6734
rect 412192 6526 412220 8092
rect 413296 6882 413324 8092
rect 413204 6854 413324 6882
rect 412180 6520 412232 6526
rect 412180 6462 412232 6468
rect 413204 6322 413232 6854
rect 413284 6588 413336 6594
rect 413284 6530 413336 6536
rect 413192 6316 413244 6322
rect 413192 6258 413244 6264
rect 413296 480 413324 6530
rect 414112 6248 414164 6254
rect 414112 6190 414164 6196
rect 413928 5772 413980 5778
rect 413928 5714 413980 5720
rect 413376 5704 413428 5710
rect 413376 5646 413428 5652
rect 413388 3670 413416 5646
rect 413376 3664 413428 3670
rect 413376 3606 413428 3612
rect 413940 3466 413968 5714
rect 413928 3460 413980 3466
rect 413928 3402 413980 3408
rect 414124 3194 414152 6190
rect 414400 6118 414428 8092
rect 415596 6798 415624 8092
rect 415584 6792 415636 6798
rect 415584 6734 415636 6740
rect 414480 6724 414532 6730
rect 414480 6666 414532 6672
rect 414388 6112 414440 6118
rect 414388 6054 414440 6060
rect 414112 3188 414164 3194
rect 414112 3130 414164 3136
rect 414492 480 414520 6666
rect 416700 6594 416728 8092
rect 416688 6588 416740 6594
rect 416688 6530 416740 6536
rect 417804 6458 417832 8092
rect 419000 6662 419028 8092
rect 419172 6724 419224 6730
rect 419172 6666 419224 6672
rect 418988 6656 419040 6662
rect 418988 6598 419040 6604
rect 417792 6452 417844 6458
rect 417792 6394 417844 6400
rect 417976 6384 418028 6390
rect 417976 6326 418028 6332
rect 416688 6180 416740 6186
rect 416688 6122 416740 6128
rect 414822 6012 415386 6032
rect 414822 6010 414836 6012
rect 414892 6010 414916 6012
rect 414972 6010 414996 6012
rect 415052 6010 415076 6012
rect 415132 6010 415156 6012
rect 415212 6010 415236 6012
rect 415292 6010 415316 6012
rect 415372 6010 415386 6012
rect 415066 5958 415076 6010
rect 415132 5958 415142 6010
rect 414822 5956 414836 5958
rect 414892 5956 414916 5958
rect 414972 5956 414996 5958
rect 415052 5956 415076 5958
rect 415132 5956 415156 5958
rect 415212 5956 415236 5958
rect 415292 5956 415316 5958
rect 415372 5956 415386 5958
rect 414822 5936 415386 5956
rect 414822 4924 415386 4944
rect 414822 4922 414836 4924
rect 414892 4922 414916 4924
rect 414972 4922 414996 4924
rect 415052 4922 415076 4924
rect 415132 4922 415156 4924
rect 415212 4922 415236 4924
rect 415292 4922 415316 4924
rect 415372 4922 415386 4924
rect 415066 4870 415076 4922
rect 415132 4870 415142 4922
rect 414822 4868 414836 4870
rect 414892 4868 414916 4870
rect 414972 4868 414996 4870
rect 415052 4868 415076 4870
rect 415132 4868 415156 4870
rect 415212 4868 415236 4870
rect 415292 4868 415316 4870
rect 415372 4868 415386 4870
rect 414822 4848 415386 4868
rect 416700 4026 416728 6122
rect 416700 3998 416912 4026
rect 414822 3836 415386 3856
rect 414822 3834 414836 3836
rect 414892 3834 414916 3836
rect 414972 3834 414996 3836
rect 415052 3834 415076 3836
rect 415132 3834 415156 3836
rect 415212 3834 415236 3836
rect 415292 3834 415316 3836
rect 415372 3834 415386 3836
rect 415066 3782 415076 3834
rect 415132 3782 415142 3834
rect 414822 3780 414836 3782
rect 414892 3780 414916 3782
rect 414972 3780 414996 3782
rect 415052 3780 415076 3782
rect 415132 3780 415156 3782
rect 415212 3780 415236 3782
rect 415292 3780 415316 3782
rect 415372 3780 415386 3782
rect 414822 3760 415386 3780
rect 415676 3188 415728 3194
rect 415676 3130 415728 3136
rect 414822 2748 415386 2768
rect 414822 2746 414836 2748
rect 414892 2746 414916 2748
rect 414972 2746 414996 2748
rect 415052 2746 415076 2748
rect 415132 2746 415156 2748
rect 415212 2746 415236 2748
rect 415292 2746 415316 2748
rect 415372 2746 415386 2748
rect 415066 2694 415076 2746
rect 415132 2694 415142 2746
rect 414822 2692 414836 2694
rect 414892 2692 414916 2694
rect 414972 2692 414996 2694
rect 415052 2692 415076 2694
rect 415132 2692 415156 2694
rect 415212 2692 415236 2694
rect 415292 2692 415316 2694
rect 415372 2692 415386 2694
rect 414822 2672 415386 2692
rect 415688 480 415716 3130
rect 416884 480 416912 3998
rect 417988 480 418016 6326
rect 418160 5908 418212 5914
rect 418160 5850 418212 5856
rect 418172 3194 418200 5850
rect 418160 3188 418212 3194
rect 418160 3130 418212 3136
rect 419184 480 419212 6666
rect 420104 6254 420132 8092
rect 421208 6390 421236 8092
rect 421196 6384 421248 6390
rect 421196 6326 421248 6332
rect 420092 6248 420144 6254
rect 420092 6190 420144 6196
rect 422404 6186 422432 8092
rect 423508 6866 423536 8092
rect 423496 6860 423548 6866
rect 423496 6802 423548 6808
rect 424612 6526 424640 8092
rect 423588 6520 423640 6526
rect 423588 6462 423640 6468
rect 424600 6520 424652 6526
rect 424600 6462 424652 6468
rect 422392 6180 422444 6186
rect 422392 6122 422444 6128
rect 421564 3664 421616 3670
rect 421564 3606 421616 3612
rect 420368 3188 420420 3194
rect 420368 3130 420420 3136
rect 420380 480 420408 3130
rect 421576 480 421604 3606
rect 423600 3482 423628 6462
rect 424968 6316 425020 6322
rect 424968 6258 425020 6264
rect 424324 6112 424376 6118
rect 424324 6054 424376 6060
rect 422760 3460 422812 3466
rect 423600 3454 423996 3482
rect 422760 3402 422812 3408
rect 422772 480 422800 3402
rect 423968 480 423996 3454
rect 424336 3126 424364 6054
rect 424980 3346 425008 6258
rect 425716 5574 425744 8092
rect 426912 6798 426940 8092
rect 426532 6792 426584 6798
rect 426532 6734 426584 6740
rect 426900 6792 426952 6798
rect 426900 6734 426952 6740
rect 426544 6594 426572 6734
rect 426440 6588 426492 6594
rect 426440 6530 426492 6536
rect 426532 6588 426584 6594
rect 426532 6530 426584 6536
rect 427544 6588 427596 6594
rect 427544 6530 427596 6536
rect 425704 5568 425756 5574
rect 425704 5510 425756 5516
rect 426452 3466 426480 6530
rect 426440 3460 426492 3466
rect 426440 3402 426492 3408
rect 424980 3318 425192 3346
rect 424324 3120 424376 3126
rect 424324 3062 424376 3068
rect 425164 480 425192 3318
rect 426348 3120 426400 3126
rect 426348 3062 426400 3068
rect 426360 480 426388 3062
rect 427556 480 427584 6530
rect 427820 6452 427872 6458
rect 427820 6394 427872 6400
rect 427832 3194 427860 6394
rect 428016 6186 428044 8092
rect 429120 6322 429148 8092
rect 429200 6656 429252 6662
rect 429200 6598 429252 6604
rect 429108 6316 429160 6322
rect 429108 6258 429160 6264
rect 428004 6180 428056 6186
rect 428004 6122 428056 6128
rect 428832 5568 428884 5574
rect 428832 5510 428884 5516
rect 428844 3466 428872 5510
rect 428740 3460 428792 3466
rect 428740 3402 428792 3408
rect 428832 3460 428884 3466
rect 428832 3402 428884 3408
rect 427820 3188 427872 3194
rect 427820 3130 427872 3136
rect 428752 480 428780 3402
rect 429212 3398 429240 6598
rect 430316 6594 430344 8092
rect 431420 6662 431448 8092
rect 431408 6656 431460 6662
rect 431408 6598 431460 6604
rect 430304 6588 430356 6594
rect 430304 6530 430356 6536
rect 432524 6254 432552 8092
rect 432696 6384 432748 6390
rect 432696 6326 432748 6332
rect 430580 6248 430632 6254
rect 430580 6190 430632 6196
rect 432512 6248 432564 6254
rect 432512 6190 432564 6196
rect 429200 3392 429252 3398
rect 429200 3334 429252 3340
rect 430592 3194 430620 6190
rect 432708 4078 432736 6326
rect 433720 5846 433748 8092
rect 433892 6860 433944 6866
rect 433892 6802 433944 6808
rect 433708 5840 433760 5846
rect 433708 5782 433760 5788
rect 432822 5468 433386 5488
rect 432822 5466 432836 5468
rect 432892 5466 432916 5468
rect 432972 5466 432996 5468
rect 433052 5466 433076 5468
rect 433132 5466 433156 5468
rect 433212 5466 433236 5468
rect 433292 5466 433316 5468
rect 433372 5466 433386 5468
rect 433066 5414 433076 5466
rect 433132 5414 433142 5466
rect 432822 5412 432836 5414
rect 432892 5412 432916 5414
rect 432972 5412 432996 5414
rect 433052 5412 433076 5414
rect 433132 5412 433156 5414
rect 433212 5412 433236 5414
rect 433292 5412 433316 5414
rect 433372 5412 433386 5414
rect 432822 5392 433386 5412
rect 432822 4380 433386 4400
rect 432822 4378 432836 4380
rect 432892 4378 432916 4380
rect 432972 4378 432996 4380
rect 433052 4378 433076 4380
rect 433132 4378 433156 4380
rect 433212 4378 433236 4380
rect 433292 4378 433316 4380
rect 433372 4378 433386 4380
rect 433066 4326 433076 4378
rect 433132 4326 433142 4378
rect 432822 4324 432836 4326
rect 432892 4324 432916 4326
rect 432972 4324 432996 4326
rect 433052 4324 433076 4326
rect 433132 4324 433156 4326
rect 433212 4324 433236 4326
rect 433292 4324 433316 4326
rect 433372 4324 433386 4326
rect 432822 4304 433386 4324
rect 432696 4072 432748 4078
rect 432696 4014 432748 4020
rect 433524 4072 433576 4078
rect 433524 4014 433576 4020
rect 431132 3392 431184 3398
rect 431132 3334 431184 3340
rect 429936 3188 429988 3194
rect 429936 3130 429988 3136
rect 430580 3188 430632 3194
rect 430580 3130 430632 3136
rect 429948 480 429976 3130
rect 431144 480 431172 3334
rect 432822 3292 433386 3312
rect 432822 3290 432836 3292
rect 432892 3290 432916 3292
rect 432972 3290 432996 3292
rect 433052 3290 433076 3292
rect 433132 3290 433156 3292
rect 433212 3290 433236 3292
rect 433292 3290 433316 3292
rect 433372 3290 433386 3292
rect 433066 3238 433076 3290
rect 433132 3238 433142 3290
rect 432822 3236 432836 3238
rect 432892 3236 432916 3238
rect 432972 3236 432996 3238
rect 433052 3236 433076 3238
rect 433132 3236 433156 3238
rect 433212 3236 433236 3238
rect 433292 3236 433316 3238
rect 433372 3236 433386 3238
rect 432822 3216 433386 3236
rect 432328 3188 432380 3194
rect 432328 3130 432380 3136
rect 432340 480 432368 3130
rect 432822 2204 433386 2224
rect 432822 2202 432836 2204
rect 432892 2202 432916 2204
rect 432972 2202 432996 2204
rect 433052 2202 433076 2204
rect 433132 2202 433156 2204
rect 433212 2202 433236 2204
rect 433292 2202 433316 2204
rect 433372 2202 433386 2204
rect 433066 2150 433076 2202
rect 433132 2150 433142 2202
rect 432822 2148 432836 2150
rect 432892 2148 432916 2150
rect 432972 2148 432996 2150
rect 433052 2148 433076 2150
rect 433132 2148 433156 2150
rect 433212 2148 433236 2150
rect 433292 2148 433316 2150
rect 433372 2148 433386 2150
rect 432822 2128 433386 2148
rect 433536 480 433564 4014
rect 433904 3602 433932 6802
rect 434824 6730 434852 8092
rect 434812 6724 434864 6730
rect 434812 6666 434864 6672
rect 434536 6520 434588 6526
rect 434536 6462 434588 6468
rect 434548 4146 434576 6462
rect 435928 6458 435956 8092
rect 437124 6526 437152 8092
rect 437480 6792 437532 6798
rect 437480 6734 437532 6740
rect 437112 6520 437164 6526
rect 437112 6462 437164 6468
rect 435916 6452 435968 6458
rect 435916 6394 435968 6400
rect 434628 6112 434680 6118
rect 434628 6054 434680 6060
rect 434536 4140 434588 4146
rect 434536 4082 434588 4088
rect 433892 3596 433944 3602
rect 433892 3538 433944 3544
rect 434640 480 434668 6054
rect 437020 4140 437072 4146
rect 437020 4082 437072 4088
rect 435824 3596 435876 3602
rect 435824 3538 435876 3544
rect 435836 480 435864 3538
rect 437032 480 437060 4082
rect 437492 3398 437520 6734
rect 438228 6390 438256 8092
rect 439044 6588 439096 6594
rect 439044 6530 439096 6536
rect 438216 6384 438268 6390
rect 438216 6326 438268 6332
rect 438860 6316 438912 6322
rect 438860 6258 438912 6264
rect 438216 3460 438268 3466
rect 438216 3402 438268 3408
rect 437480 3392 437532 3398
rect 437480 3334 437532 3340
rect 438228 480 438256 3402
rect 438872 3126 438900 6258
rect 438952 6180 439004 6186
rect 438952 6122 439004 6128
rect 438964 3194 438992 6122
rect 438952 3188 439004 3194
rect 438952 3130 439004 3136
rect 438860 3120 438912 3126
rect 438860 3062 438912 3068
rect 439056 3058 439084 6530
rect 439332 6118 439360 8092
rect 439320 6112 439372 6118
rect 439320 6054 439372 6060
rect 440528 5710 440556 8092
rect 441632 6798 441660 8092
rect 441620 6792 441672 6798
rect 441620 6734 441672 6740
rect 442356 6656 442408 6662
rect 442356 6598 442408 6604
rect 440516 5704 440568 5710
rect 440516 5646 440568 5652
rect 442368 3398 442396 6598
rect 442736 6594 442764 8092
rect 442724 6588 442776 6594
rect 442724 6530 442776 6536
rect 443932 6322 443960 8092
rect 443920 6316 443972 6322
rect 443920 6258 443972 6264
rect 443552 6248 443604 6254
rect 443552 6190 443604 6196
rect 439412 3392 439464 3398
rect 439412 3334 439464 3340
rect 442356 3392 442408 3398
rect 442356 3334 442408 3340
rect 439044 3052 439096 3058
rect 439044 2994 439096 3000
rect 439424 480 439452 3334
rect 443564 3194 443592 6190
rect 445036 5914 445064 8092
rect 445852 6724 445904 6730
rect 445852 6666 445904 6672
rect 445760 6452 445812 6458
rect 445760 6394 445812 6400
rect 445024 5908 445076 5914
rect 445024 5850 445076 5856
rect 444380 5840 444432 5846
rect 444380 5782 444432 5788
rect 444288 5704 444340 5710
rect 444288 5646 444340 5652
rect 444300 3466 444328 5646
rect 444288 3460 444340 3466
rect 444288 3402 444340 3408
rect 444196 3392 444248 3398
rect 444196 3334 444248 3340
rect 440608 3188 440660 3194
rect 440608 3130 440660 3136
rect 443552 3188 443604 3194
rect 443552 3130 443604 3136
rect 440620 480 440648 3130
rect 441804 3120 441856 3126
rect 441804 3062 441856 3068
rect 441816 480 441844 3062
rect 443000 3052 443052 3058
rect 443000 2994 443052 3000
rect 443012 480 443040 2994
rect 444208 480 444236 3334
rect 444392 3058 444420 5782
rect 445772 4078 445800 6394
rect 445760 4072 445812 4078
rect 445760 4014 445812 4020
rect 445864 3398 445892 6666
rect 446140 6662 446168 8092
rect 446128 6656 446180 6662
rect 446128 6598 446180 6604
rect 447140 6520 447192 6526
rect 447140 6462 447192 6468
rect 445852 3392 445904 3398
rect 445852 3334 445904 3340
rect 445392 3188 445444 3194
rect 445392 3130 445444 3136
rect 444380 3052 444432 3058
rect 444380 2994 444432 3000
rect 445404 480 445432 3130
rect 447152 3126 447180 6462
rect 447336 6254 447364 8092
rect 448440 6458 448468 8092
rect 449544 6730 449572 8092
rect 449532 6724 449584 6730
rect 449532 6666 449584 6672
rect 448428 6452 448480 6458
rect 448428 6394 448480 6400
rect 450740 6390 450768 8092
rect 451844 6866 451872 8092
rect 451832 6860 451884 6866
rect 451832 6802 451884 6808
rect 448612 6384 448664 6390
rect 448612 6326 448664 6332
rect 450728 6384 450780 6390
rect 450728 6326 450780 6332
rect 447324 6248 447376 6254
rect 447324 6190 447376 6196
rect 448520 6112 448572 6118
rect 448520 6054 448572 6060
rect 448532 4146 448560 6054
rect 448520 4140 448572 4146
rect 448520 4082 448572 4088
rect 447784 3392 447836 3398
rect 447784 3334 447836 3340
rect 447140 3120 447192 3126
rect 447140 3062 447192 3068
rect 446588 3052 446640 3058
rect 446588 2994 446640 3000
rect 446600 480 446628 2994
rect 447796 480 447824 3334
rect 448624 3194 448652 6326
rect 452948 6186 452976 8092
rect 453120 6792 453172 6798
rect 453120 6734 453172 6740
rect 452936 6180 452988 6186
rect 452936 6122 452988 6128
rect 450822 6012 451386 6032
rect 450822 6010 450836 6012
rect 450892 6010 450916 6012
rect 450972 6010 450996 6012
rect 451052 6010 451076 6012
rect 451132 6010 451156 6012
rect 451212 6010 451236 6012
rect 451292 6010 451316 6012
rect 451372 6010 451386 6012
rect 451066 5958 451076 6010
rect 451132 5958 451142 6010
rect 450822 5956 450836 5958
rect 450892 5956 450916 5958
rect 450972 5956 450996 5958
rect 451052 5956 451076 5958
rect 451132 5956 451156 5958
rect 451212 5956 451236 5958
rect 451292 5956 451316 5958
rect 451372 5956 451386 5958
rect 450822 5936 451386 5956
rect 450822 4924 451386 4944
rect 450822 4922 450836 4924
rect 450892 4922 450916 4924
rect 450972 4922 450996 4924
rect 451052 4922 451076 4924
rect 451132 4922 451156 4924
rect 451212 4922 451236 4924
rect 451292 4922 451316 4924
rect 451372 4922 451386 4924
rect 451066 4870 451076 4922
rect 451132 4870 451142 4922
rect 450822 4868 450836 4870
rect 450892 4868 450916 4870
rect 450972 4868 450996 4870
rect 451052 4868 451076 4870
rect 451132 4868 451156 4870
rect 451212 4868 451236 4870
rect 451292 4868 451316 4870
rect 451372 4868 451386 4870
rect 450822 4848 451386 4868
rect 452476 4140 452528 4146
rect 452476 4082 452528 4088
rect 448980 4072 449032 4078
rect 448980 4014 449032 4020
rect 448612 3188 448664 3194
rect 448612 3130 448664 3136
rect 448992 480 449020 4014
rect 450822 3836 451386 3856
rect 450822 3834 450836 3836
rect 450892 3834 450916 3836
rect 450972 3834 450996 3836
rect 451052 3834 451076 3836
rect 451132 3834 451156 3836
rect 451212 3834 451236 3836
rect 451292 3834 451316 3836
rect 451372 3834 451386 3836
rect 451066 3782 451076 3834
rect 451132 3782 451142 3834
rect 450822 3780 450836 3782
rect 450892 3780 450916 3782
rect 450972 3780 450996 3782
rect 451052 3780 451076 3782
rect 451132 3780 451156 3782
rect 451212 3780 451236 3782
rect 451292 3780 451316 3782
rect 451372 3780 451386 3782
rect 450822 3760 451386 3780
rect 451464 3188 451516 3194
rect 451464 3130 451516 3136
rect 450176 3120 450228 3126
rect 450176 3062 450228 3068
rect 450188 480 450216 3062
rect 450822 2748 451386 2768
rect 450822 2746 450836 2748
rect 450892 2746 450916 2748
rect 450972 2746 450996 2748
rect 451052 2746 451076 2748
rect 451132 2746 451156 2748
rect 451212 2746 451236 2748
rect 451292 2746 451316 2748
rect 451372 2746 451386 2748
rect 451066 2694 451076 2746
rect 451132 2694 451142 2746
rect 450822 2692 450836 2694
rect 450892 2692 450916 2694
rect 450972 2692 450996 2694
rect 451052 2692 451076 2694
rect 451132 2692 451156 2694
rect 451212 2692 451236 2694
rect 451292 2692 451316 2694
rect 451372 2692 451386 2694
rect 450822 2672 451386 2692
rect 451476 2530 451504 3130
rect 451292 2502 451504 2530
rect 451292 480 451320 2502
rect 452488 480 452516 4082
rect 453132 3398 453160 6734
rect 454144 6594 454172 8092
rect 453672 6588 453724 6594
rect 453672 6530 453724 6536
rect 454132 6588 454184 6594
rect 454132 6530 454184 6536
rect 453684 4146 453712 6530
rect 454132 6316 454184 6322
rect 454132 6258 454184 6264
rect 453672 4140 453724 4146
rect 453672 4082 453724 4088
rect 453672 3460 453724 3466
rect 453672 3402 453724 3408
rect 453120 3392 453172 3398
rect 453120 3334 453172 3340
rect 453684 480 453712 3402
rect 454144 3194 454172 6258
rect 455248 6118 455276 8092
rect 455236 6112 455288 6118
rect 455236 6054 455288 6060
rect 454684 5908 454736 5914
rect 454684 5850 454736 5856
rect 454132 3188 454184 3194
rect 454132 3130 454184 3136
rect 454696 3126 454724 5850
rect 456352 5574 456380 8092
rect 456800 6656 456852 6662
rect 456800 6598 456852 6604
rect 456340 5568 456392 5574
rect 456340 5510 456392 5516
rect 456064 4140 456116 4146
rect 456064 4082 456116 4088
rect 454868 3392 454920 3398
rect 454868 3334 454920 3340
rect 454684 3120 454736 3126
rect 454684 3062 454736 3068
rect 454880 480 454908 3334
rect 456076 480 456104 4082
rect 456812 3602 456840 6598
rect 457548 6526 457576 8092
rect 457536 6520 457588 6526
rect 457536 6462 457588 6468
rect 458180 6452 458232 6458
rect 458180 6394 458232 6400
rect 458192 4078 458220 6394
rect 458652 6322 458680 8092
rect 459560 6724 459612 6730
rect 459560 6666 459612 6672
rect 458640 6316 458692 6322
rect 458640 6258 458692 6264
rect 458272 6248 458324 6254
rect 458272 6190 458324 6196
rect 458180 4072 458232 4078
rect 458180 4014 458232 4020
rect 456800 3596 456852 3602
rect 456800 3538 456852 3544
rect 458284 3194 458312 6190
rect 458640 5568 458692 5574
rect 458640 5510 458692 5516
rect 458652 3466 458680 5510
rect 459572 4146 459600 6666
rect 459756 5914 459784 8092
rect 460952 6730 460980 8092
rect 462056 6798 462084 8092
rect 462044 6792 462096 6798
rect 462044 6734 462096 6740
rect 460940 6724 460992 6730
rect 460940 6666 460992 6672
rect 462228 6384 462280 6390
rect 462228 6326 462280 6332
rect 459744 5908 459796 5914
rect 459744 5850 459796 5856
rect 459560 4140 459612 4146
rect 459560 4082 459612 4088
rect 462044 4072 462096 4078
rect 462044 4014 462096 4020
rect 459652 3596 459704 3602
rect 459652 3538 459704 3544
rect 458640 3460 458692 3466
rect 458640 3402 458692 3408
rect 457260 3188 457312 3194
rect 457260 3130 457312 3136
rect 458272 3188 458324 3194
rect 458272 3130 458324 3136
rect 457272 480 457300 3130
rect 458456 3120 458508 3126
rect 458456 3062 458508 3068
rect 458468 480 458496 3062
rect 459664 480 459692 3538
rect 460848 3188 460900 3194
rect 460848 3130 460900 3136
rect 460860 480 460888 3130
rect 462056 480 462084 4014
rect 462240 3466 462268 6326
rect 463160 6254 463188 8092
rect 463332 6860 463384 6866
rect 463332 6802 463384 6808
rect 463148 6248 463200 6254
rect 463148 6190 463200 6196
rect 463240 4140 463292 4146
rect 463240 4082 463292 4088
rect 462228 3460 462280 3466
rect 462228 3402 462280 3408
rect 463252 480 463280 4082
rect 463344 3602 463372 6802
rect 464264 6662 464292 8092
rect 464252 6656 464304 6662
rect 464252 6598 464304 6604
rect 464436 6588 464488 6594
rect 464436 6530 464488 6536
rect 463700 6180 463752 6186
rect 463700 6122 463752 6128
rect 463332 3596 463384 3602
rect 463332 3538 463384 3544
rect 463712 3126 463740 6122
rect 464252 6112 464304 6118
rect 464252 6054 464304 6060
rect 463700 3120 463752 3126
rect 463700 3062 463752 3068
rect 464264 3058 464292 6054
rect 464448 3738 464476 6530
rect 465460 6118 465488 8092
rect 466564 6458 466592 8092
rect 467668 6594 467696 8092
rect 467656 6588 467708 6594
rect 467656 6530 467708 6536
rect 467840 6520 467892 6526
rect 467840 6462 467892 6468
rect 466552 6452 466604 6458
rect 466552 6394 466604 6400
rect 465448 6112 465500 6118
rect 465448 6054 465500 6060
rect 467852 4078 467880 6462
rect 468864 6390 468892 8092
rect 468852 6384 468904 6390
rect 468852 6326 468904 6332
rect 469496 6316 469548 6322
rect 469496 6258 469548 6264
rect 469404 5908 469456 5914
rect 469404 5850 469456 5856
rect 468822 5468 469386 5488
rect 468822 5466 468836 5468
rect 468892 5466 468916 5468
rect 468972 5466 468996 5468
rect 469052 5466 469076 5468
rect 469132 5466 469156 5468
rect 469212 5466 469236 5468
rect 469292 5466 469316 5468
rect 469372 5466 469386 5468
rect 469066 5414 469076 5466
rect 469132 5414 469142 5466
rect 468822 5412 468836 5414
rect 468892 5412 468916 5414
rect 468972 5412 468996 5414
rect 469052 5412 469076 5414
rect 469132 5412 469156 5414
rect 469212 5412 469236 5414
rect 469292 5412 469316 5414
rect 469372 5412 469386 5414
rect 468822 5392 469386 5412
rect 468822 4380 469386 4400
rect 468822 4378 468836 4380
rect 468892 4378 468916 4380
rect 468972 4378 468996 4380
rect 469052 4378 469076 4380
rect 469132 4378 469156 4380
rect 469212 4378 469236 4380
rect 469292 4378 469316 4380
rect 469372 4378 469386 4380
rect 469066 4326 469076 4378
rect 469132 4326 469142 4378
rect 468822 4324 468836 4326
rect 468892 4324 468916 4326
rect 468972 4324 468996 4326
rect 469052 4324 469076 4326
rect 469132 4324 469156 4326
rect 469212 4324 469236 4326
rect 469292 4324 469316 4326
rect 469372 4324 469386 4326
rect 468822 4304 469386 4324
rect 467840 4072 467892 4078
rect 467840 4014 467892 4020
rect 464436 3732 464488 3738
rect 464436 3674 464488 3680
rect 467932 3732 467984 3738
rect 467932 3674 467984 3680
rect 465632 3596 465684 3602
rect 465632 3538 465684 3544
rect 464436 3460 464488 3466
rect 464436 3402 464488 3408
rect 464252 3052 464304 3058
rect 464252 2994 464304 3000
rect 464448 480 464476 3402
rect 465644 480 465672 3538
rect 466828 3120 466880 3126
rect 466828 3062 466880 3068
rect 466840 480 466868 3062
rect 467944 480 467972 3674
rect 469416 3466 469444 5850
rect 469508 3738 469536 6258
rect 469968 5846 469996 8092
rect 469956 5840 470008 5846
rect 469956 5782 470008 5788
rect 471072 5574 471100 8092
rect 472268 6526 472296 8092
rect 473372 6866 473400 8092
rect 473360 6860 473412 6866
rect 473360 6802 473412 6808
rect 472900 6792 472952 6798
rect 472900 6734 472952 6740
rect 472532 6724 472584 6730
rect 472532 6666 472584 6672
rect 472256 6520 472308 6526
rect 472256 6462 472308 6468
rect 471060 5568 471112 5574
rect 471060 5510 471112 5516
rect 472544 4146 472572 6666
rect 472532 4140 472584 4146
rect 472532 4082 472584 4088
rect 471520 4072 471572 4078
rect 471520 4014 471572 4020
rect 469496 3732 469548 3738
rect 469496 3674 469548 3680
rect 469404 3460 469456 3466
rect 469404 3402 469456 3408
rect 470324 3392 470376 3398
rect 470324 3334 470376 3340
rect 468822 3292 469386 3312
rect 468822 3290 468836 3292
rect 468892 3290 468916 3292
rect 468972 3290 468996 3292
rect 469052 3290 469076 3292
rect 469132 3290 469156 3292
rect 469212 3290 469236 3292
rect 469292 3290 469316 3292
rect 469372 3290 469386 3292
rect 469066 3238 469076 3290
rect 469132 3238 469142 3290
rect 468822 3236 468836 3238
rect 468892 3236 468916 3238
rect 468972 3236 468996 3238
rect 469052 3236 469076 3238
rect 469132 3236 469156 3238
rect 469212 3236 469236 3238
rect 469292 3236 469316 3238
rect 469372 3236 469386 3238
rect 468822 3216 469386 3236
rect 468668 3052 468720 3058
rect 468668 2994 468720 3000
rect 468680 1986 468708 2994
rect 468822 2204 469386 2224
rect 468822 2202 468836 2204
rect 468892 2202 468916 2204
rect 468972 2202 468996 2204
rect 469052 2202 469076 2204
rect 469132 2202 469156 2204
rect 469212 2202 469236 2204
rect 469292 2202 469316 2204
rect 469372 2202 469386 2204
rect 469066 2150 469076 2202
rect 469132 2150 469142 2202
rect 468822 2148 468836 2150
rect 468892 2148 468916 2150
rect 468972 2148 468996 2150
rect 469052 2148 469076 2150
rect 469132 2148 469156 2150
rect 469212 2148 469236 2150
rect 469292 2148 469316 2150
rect 469372 2148 469386 2150
rect 468822 2128 469386 2148
rect 468680 1958 469168 1986
rect 469140 480 469168 1958
rect 470336 480 470364 3334
rect 471532 480 471560 4014
rect 472716 3732 472768 3738
rect 472716 3674 472768 3680
rect 472728 480 472756 3674
rect 472912 3670 472940 6734
rect 474096 6248 474148 6254
rect 474096 6190 474148 6196
rect 474108 3738 474136 6190
rect 474476 6186 474504 8092
rect 474740 6656 474792 6662
rect 474740 6598 474792 6604
rect 474464 6180 474516 6186
rect 474464 6122 474516 6128
rect 474648 5568 474700 5574
rect 474648 5510 474700 5516
rect 474096 3732 474148 3738
rect 474096 3674 474148 3680
rect 472900 3664 472952 3670
rect 472900 3606 472952 3612
rect 474660 3534 474688 5510
rect 474648 3528 474700 3534
rect 474648 3470 474700 3476
rect 474752 3466 474780 6598
rect 475672 6254 475700 8092
rect 476776 6730 476804 8092
rect 476764 6724 476816 6730
rect 476764 6666 476816 6672
rect 477880 6662 477908 8092
rect 479076 6798 479104 8092
rect 479064 6792 479116 6798
rect 479064 6734 479116 6740
rect 477868 6656 477920 6662
rect 477868 6598 477920 6604
rect 477592 6588 477644 6594
rect 477592 6530 477644 6536
rect 477500 6452 477552 6458
rect 477500 6394 477552 6400
rect 475660 6248 475712 6254
rect 475660 6190 475712 6196
rect 476120 6112 476172 6118
rect 476120 6054 476172 6060
rect 475108 4140 475160 4146
rect 475108 4082 475160 4088
rect 473912 3460 473964 3466
rect 473912 3402 473964 3408
rect 474740 3460 474792 3466
rect 474740 3402 474792 3408
rect 473924 480 473952 3402
rect 475120 480 475148 4082
rect 476132 4078 476160 6054
rect 477512 4146 477540 6394
rect 477500 4140 477552 4146
rect 477500 4082 477552 4088
rect 476120 4072 476172 4078
rect 476120 4014 476172 4020
rect 477500 3732 477552 3738
rect 477500 3674 477552 3680
rect 476304 3664 476356 3670
rect 476304 3606 476356 3612
rect 476316 480 476344 3606
rect 477512 480 477540 3674
rect 477604 3398 477632 6530
rect 478972 6384 479024 6390
rect 478972 6326 479024 6332
rect 478880 5840 478932 5846
rect 478880 5782 478932 5788
rect 478892 3534 478920 5782
rect 478984 3670 479012 6326
rect 480180 6322 480208 8092
rect 481284 6458 481312 8092
rect 482480 6594 482508 8092
rect 482468 6588 482520 6594
rect 482468 6530 482520 6536
rect 483296 6520 483348 6526
rect 483296 6462 483348 6468
rect 481272 6452 481324 6458
rect 481272 6394 481324 6400
rect 480168 6316 480220 6322
rect 480168 6258 480220 6264
rect 481088 4140 481140 4146
rect 481088 4082 481140 4088
rect 479892 4072 479944 4078
rect 479892 4014 479944 4020
rect 478972 3664 479024 3670
rect 478972 3606 479024 3612
rect 478880 3528 478932 3534
rect 478880 3470 478932 3476
rect 478696 3460 478748 3466
rect 478696 3402 478748 3408
rect 477592 3392 477644 3398
rect 477592 3334 477644 3340
rect 478708 480 478736 3402
rect 479904 480 479932 4014
rect 481100 480 481128 4082
rect 482284 3392 482336 3398
rect 482284 3334 482336 3340
rect 482296 480 482324 3334
rect 483308 3194 483336 6462
rect 483584 6390 483612 8092
rect 484400 6860 484452 6866
rect 484400 6802 484452 6808
rect 483572 6384 483624 6390
rect 483572 6326 483624 6332
rect 484412 4146 484440 6802
rect 484688 6526 484716 8092
rect 485884 6866 485912 8092
rect 485872 6860 485924 6866
rect 485872 6802 485924 6808
rect 484676 6520 484728 6526
rect 484676 6462 484728 6468
rect 486988 6254 487016 8092
rect 487436 6724 487488 6730
rect 487436 6666 487488 6672
rect 484676 6248 484728 6254
rect 484676 6190 484728 6196
rect 486976 6248 487028 6254
rect 486976 6190 487028 6196
rect 484400 4140 484452 4146
rect 484400 4082 484452 4088
rect 483480 3664 483532 3670
rect 483480 3606 483532 3612
rect 483296 3188 483348 3194
rect 483296 3130 483348 3136
rect 483492 480 483520 3606
rect 484584 3528 484636 3534
rect 484584 3470 484636 3476
rect 484596 480 484624 3470
rect 484688 3126 484716 6190
rect 486822 6012 487386 6032
rect 486822 6010 486836 6012
rect 486892 6010 486916 6012
rect 486972 6010 486996 6012
rect 487052 6010 487076 6012
rect 487132 6010 487156 6012
rect 487212 6010 487236 6012
rect 487292 6010 487316 6012
rect 487372 6010 487386 6012
rect 487066 5958 487076 6010
rect 487132 5958 487142 6010
rect 486822 5956 486836 5958
rect 486892 5956 486916 5958
rect 486972 5956 486996 5958
rect 487052 5956 487076 5958
rect 487132 5956 487156 5958
rect 487212 5956 487236 5958
rect 487292 5956 487316 5958
rect 487372 5956 487386 5958
rect 486822 5936 487386 5956
rect 486822 4924 487386 4944
rect 486822 4922 486836 4924
rect 486892 4922 486916 4924
rect 486972 4922 486996 4924
rect 487052 4922 487076 4924
rect 487132 4922 487156 4924
rect 487212 4922 487236 4924
rect 487292 4922 487316 4924
rect 487372 4922 487386 4924
rect 487066 4870 487076 4922
rect 487132 4870 487142 4922
rect 486822 4868 486836 4870
rect 486892 4868 486916 4870
rect 486972 4868 486996 4870
rect 487052 4868 487076 4870
rect 487132 4868 487156 4870
rect 487212 4868 487236 4870
rect 487292 4868 487316 4870
rect 487372 4868 487386 4870
rect 486822 4848 487386 4868
rect 486822 3836 487386 3856
rect 486822 3834 486836 3836
rect 486892 3834 486916 3836
rect 486972 3834 486996 3836
rect 487052 3834 487076 3836
rect 487132 3834 487156 3836
rect 487212 3834 487236 3836
rect 487292 3834 487316 3836
rect 487372 3834 487386 3836
rect 487066 3782 487076 3834
rect 487132 3782 487142 3834
rect 486822 3780 486836 3782
rect 486892 3780 486916 3782
rect 486972 3780 486996 3782
rect 487052 3780 487076 3782
rect 487132 3780 487156 3782
rect 487212 3780 487236 3782
rect 487292 3780 487316 3782
rect 487372 3780 487386 3782
rect 486822 3760 487386 3780
rect 485780 3460 485832 3466
rect 485780 3402 485832 3408
rect 484676 3120 484728 3126
rect 484676 3062 484728 3068
rect 485792 480 485820 3402
rect 487448 3398 487476 6666
rect 488092 5642 488120 8092
rect 488540 6656 488592 6662
rect 488540 6598 488592 6604
rect 488080 5636 488132 5642
rect 488080 5578 488132 5584
rect 488172 4140 488224 4146
rect 488172 4082 488224 4088
rect 487436 3392 487488 3398
rect 487436 3334 487488 3340
rect 486700 3188 486752 3194
rect 486700 3130 486752 3136
rect 486712 2530 486740 3130
rect 486822 2748 487386 2768
rect 486822 2746 486836 2748
rect 486892 2746 486916 2748
rect 486972 2746 486996 2748
rect 487052 2746 487076 2748
rect 487132 2746 487156 2748
rect 487212 2746 487236 2748
rect 487292 2746 487316 2748
rect 487372 2746 487386 2748
rect 487066 2694 487076 2746
rect 487132 2694 487142 2746
rect 486822 2692 486836 2694
rect 486892 2692 486916 2694
rect 486972 2692 486996 2694
rect 487052 2692 487076 2694
rect 487132 2692 487156 2694
rect 487212 2692 487236 2694
rect 487292 2692 487316 2694
rect 487372 2692 487386 2694
rect 486822 2672 487386 2692
rect 486712 2502 487016 2530
rect 486988 480 487016 2502
rect 488184 480 488212 4082
rect 488552 3602 488580 6598
rect 489288 6186 489316 8092
rect 489184 6180 489236 6186
rect 489184 6122 489236 6128
rect 489276 6180 489328 6186
rect 489276 6122 489328 6128
rect 489196 6066 489224 6122
rect 489196 6038 489408 6066
rect 488540 3596 488592 3602
rect 488540 3538 488592 3544
rect 489380 480 489408 6038
rect 490392 5778 490420 8092
rect 491116 6792 491168 6798
rect 491116 6734 491168 6740
rect 490748 6316 490800 6322
rect 490748 6258 490800 6264
rect 490380 5772 490432 5778
rect 490380 5714 490432 5720
rect 490760 4078 490788 6258
rect 490748 4072 490800 4078
rect 490748 4014 490800 4020
rect 490564 3120 490616 3126
rect 490564 3062 490616 3068
rect 490576 480 490604 3062
rect 491128 2922 491156 6734
rect 491496 6390 491524 8092
rect 491484 6384 491536 6390
rect 491484 6326 491536 6332
rect 492692 5914 492720 8092
rect 493796 6730 493824 8092
rect 493784 6724 493836 6730
rect 493784 6666 493836 6672
rect 494900 6322 494928 8092
rect 494888 6316 494940 6322
rect 494888 6258 494940 6264
rect 496096 6118 496124 8092
rect 496820 6860 496872 6866
rect 496820 6802 496872 6808
rect 496544 6452 496596 6458
rect 496544 6394 496596 6400
rect 494152 6112 494204 6118
rect 494152 6054 494204 6060
rect 496084 6112 496136 6118
rect 496084 6054 496136 6060
rect 492680 5908 492732 5914
rect 492680 5850 492732 5856
rect 491208 5636 491260 5642
rect 491208 5578 491260 5584
rect 491220 3466 491248 5578
rect 492956 3596 493008 3602
rect 492956 3538 493008 3544
rect 491208 3460 491260 3466
rect 491208 3402 491260 3408
rect 491760 3392 491812 3398
rect 491760 3334 491812 3340
rect 491116 2916 491168 2922
rect 491116 2858 491168 2864
rect 491772 480 491800 3334
rect 492968 480 492996 3538
rect 494164 3058 494192 6054
rect 495348 4072 495400 4078
rect 495348 4014 495400 4020
rect 494152 3052 494204 3058
rect 494152 2994 494204 3000
rect 494152 2916 494204 2922
rect 494152 2858 494204 2864
rect 494164 480 494192 2858
rect 495360 480 495388 4014
rect 496556 480 496584 6394
rect 496832 3602 496860 6802
rect 497200 6458 497228 8092
rect 498304 6798 498332 8092
rect 499500 6866 499528 8092
rect 500604 6882 500632 8092
rect 499488 6860 499540 6866
rect 499488 6802 499540 6808
rect 500512 6854 500632 6882
rect 498292 6792 498344 6798
rect 498292 6734 498344 6740
rect 497740 6588 497792 6594
rect 497740 6530 497792 6536
rect 497188 6452 497240 6458
rect 497188 6394 497240 6400
rect 496820 3596 496872 3602
rect 496820 3538 496872 3544
rect 497752 480 497780 6530
rect 500132 6520 500184 6526
rect 500132 6462 500184 6468
rect 498936 3052 498988 3058
rect 498936 2994 498988 3000
rect 498948 480 498976 2994
rect 500144 480 500172 6462
rect 500512 5846 500540 6854
rect 501708 6186 501736 8092
rect 502812 6594 502840 8092
rect 503904 6724 503956 6730
rect 503904 6666 503956 6672
rect 502800 6588 502852 6594
rect 502800 6530 502852 6536
rect 502432 6248 502484 6254
rect 502432 6190 502484 6196
rect 500592 6180 500644 6186
rect 500592 6122 500644 6128
rect 501696 6180 501748 6186
rect 501696 6122 501748 6128
rect 500500 5840 500552 5846
rect 500500 5782 500552 5788
rect 500604 3126 500632 6122
rect 501236 3596 501288 3602
rect 501236 3538 501288 3544
rect 500592 3120 500644 3126
rect 500592 3062 500644 3068
rect 501248 480 501276 3538
rect 502444 480 502472 6190
rect 503628 3460 503680 3466
rect 503628 3402 503680 3408
rect 503640 480 503668 3402
rect 503916 3398 503944 6666
rect 504008 6526 504036 8092
rect 505112 6730 505140 8092
rect 505100 6724 505152 6730
rect 505100 6666 505152 6672
rect 506216 6662 506244 8092
rect 506204 6656 506256 6662
rect 506204 6598 506256 6604
rect 503996 6520 504048 6526
rect 503996 6462 504048 6468
rect 507412 6390 507440 8092
rect 507216 6384 507268 6390
rect 507216 6326 507268 6332
rect 507400 6384 507452 6390
rect 507400 6326 507452 6332
rect 506480 6112 506532 6118
rect 506480 6054 506532 6060
rect 503996 5908 504048 5914
rect 503996 5850 504048 5856
rect 503904 3392 503956 3398
rect 503904 3334 503956 3340
rect 504008 3058 504036 5850
rect 506020 5772 506072 5778
rect 506020 5714 506072 5720
rect 504822 5468 505386 5488
rect 504822 5466 504836 5468
rect 504892 5466 504916 5468
rect 504972 5466 504996 5468
rect 505052 5466 505076 5468
rect 505132 5466 505156 5468
rect 505212 5466 505236 5468
rect 505292 5466 505316 5468
rect 505372 5466 505386 5468
rect 505066 5414 505076 5466
rect 505132 5414 505142 5466
rect 504822 5412 504836 5414
rect 504892 5412 504916 5414
rect 504972 5412 504996 5414
rect 505052 5412 505076 5414
rect 505132 5412 505156 5414
rect 505212 5412 505236 5414
rect 505292 5412 505316 5414
rect 505372 5412 505386 5414
rect 504822 5392 505386 5412
rect 504822 4380 505386 4400
rect 504822 4378 504836 4380
rect 504892 4378 504916 4380
rect 504972 4378 504996 4380
rect 505052 4378 505076 4380
rect 505132 4378 505156 4380
rect 505212 4378 505236 4380
rect 505292 4378 505316 4380
rect 505372 4378 505386 4380
rect 505066 4326 505076 4378
rect 505132 4326 505142 4378
rect 504822 4324 504836 4326
rect 504892 4324 504916 4326
rect 504972 4324 504996 4326
rect 505052 4324 505076 4326
rect 505132 4324 505156 4326
rect 505212 4324 505236 4326
rect 505292 4324 505316 4326
rect 505372 4324 505386 4326
rect 504822 4304 505386 4324
rect 504822 3292 505386 3312
rect 504822 3290 504836 3292
rect 504892 3290 504916 3292
rect 504972 3290 504996 3292
rect 505052 3290 505076 3292
rect 505132 3290 505156 3292
rect 505212 3290 505236 3292
rect 505292 3290 505316 3292
rect 505372 3290 505386 3292
rect 505066 3238 505076 3290
rect 505132 3238 505142 3290
rect 504822 3236 504836 3238
rect 504892 3236 504916 3238
rect 504972 3236 504996 3238
rect 505052 3236 505076 3238
rect 505132 3236 505156 3238
rect 505212 3236 505236 3238
rect 505292 3236 505316 3238
rect 505372 3236 505386 3238
rect 504822 3216 505386 3236
rect 504732 3120 504784 3126
rect 504732 3062 504784 3068
rect 503996 3052 504048 3058
rect 503996 2994 504048 3000
rect 504744 1986 504772 3062
rect 504822 2204 505386 2224
rect 504822 2202 504836 2204
rect 504892 2202 504916 2204
rect 504972 2202 504996 2204
rect 505052 2202 505076 2204
rect 505132 2202 505156 2204
rect 505212 2202 505236 2204
rect 505292 2202 505316 2204
rect 505372 2202 505386 2204
rect 505066 2150 505076 2202
rect 505132 2150 505142 2202
rect 504822 2148 504836 2150
rect 504892 2148 504916 2150
rect 504972 2148 504996 2150
rect 505052 2148 505076 2150
rect 505132 2148 505156 2150
rect 505212 2148 505236 2150
rect 505292 2148 505316 2150
rect 505372 2148 505386 2150
rect 504822 2128 505386 2148
rect 504744 1958 504864 1986
rect 504836 480 504864 1958
rect 506032 480 506060 5714
rect 506492 3534 506520 6054
rect 506480 3528 506532 3534
rect 506480 3470 506532 3476
rect 507228 480 507256 6326
rect 508516 6254 508544 8092
rect 508504 6248 508556 6254
rect 508504 6190 508556 6196
rect 509620 6118 509648 8092
rect 510436 6860 510488 6866
rect 510436 6802 510488 6808
rect 509608 6112 509660 6118
rect 509608 6054 509660 6060
rect 510448 3738 510476 6802
rect 510528 6792 510580 6798
rect 510528 6734 510580 6740
rect 510436 3732 510488 3738
rect 510436 3674 510488 3680
rect 510540 3602 510568 6734
rect 510816 6474 510844 8092
rect 510724 6446 510844 6474
rect 510724 5914 510752 6446
rect 510804 6316 510856 6322
rect 510804 6258 510856 6264
rect 510712 5908 510764 5914
rect 510712 5850 510764 5856
rect 510528 3596 510580 3602
rect 510528 3538 510580 3544
rect 509608 3392 509660 3398
rect 509608 3334 509660 3340
rect 508412 3052 508464 3058
rect 508412 2994 508464 3000
rect 508424 480 508452 2994
rect 509620 480 509648 3334
rect 510816 480 510844 6258
rect 511920 5930 511948 8092
rect 511736 5902 511948 5930
rect 511736 3466 511764 5902
rect 513024 5846 513052 8092
rect 514220 6866 514248 8092
rect 514208 6860 514260 6866
rect 514208 6802 514260 6808
rect 515324 6798 515352 8092
rect 515312 6792 515364 6798
rect 515312 6734 515364 6740
rect 514760 6520 514812 6526
rect 514760 6462 514812 6468
rect 513196 6452 513248 6458
rect 513196 6394 513248 6400
rect 511908 5840 511960 5846
rect 511908 5782 511960 5788
rect 513012 5840 513064 5846
rect 513012 5782 513064 5788
rect 511724 3460 511776 3466
rect 511724 3402 511776 3408
rect 511920 2990 511948 5782
rect 512000 3528 512052 3534
rect 512000 3470 512052 3476
rect 511908 2984 511960 2990
rect 511908 2926 511960 2932
rect 512012 480 512040 3470
rect 513208 480 513236 6394
rect 514392 3596 514444 3602
rect 514392 3538 514444 3544
rect 514404 480 514432 3538
rect 514772 3194 514800 6462
rect 516428 6322 516456 8092
rect 517624 6526 517652 8092
rect 517612 6520 517664 6526
rect 517612 6462 517664 6468
rect 516416 6316 516468 6322
rect 516416 6258 516468 6264
rect 517888 6180 517940 6186
rect 517888 6122 517940 6128
rect 515588 3732 515640 3738
rect 515588 3674 515640 3680
rect 514760 3188 514812 3194
rect 514760 3130 514812 3136
rect 515600 480 515628 3674
rect 516784 2984 516836 2990
rect 516784 2926 516836 2932
rect 516796 480 516824 2926
rect 517900 480 517928 6122
rect 518728 3670 518756 8092
rect 519084 6588 519136 6594
rect 519084 6530 519136 6536
rect 518716 3664 518768 3670
rect 518716 3606 518768 3612
rect 519096 480 519124 6530
rect 519832 3602 519860 8092
rect 520832 6656 520884 6662
rect 520832 6598 520884 6604
rect 519820 3596 519872 3602
rect 519820 3538 519872 3544
rect 520844 3398 520872 6598
rect 521028 6594 521056 8092
rect 521476 6724 521528 6730
rect 521476 6666 521528 6672
rect 521016 6588 521068 6594
rect 521016 6530 521068 6536
rect 521200 6112 521252 6118
rect 521200 6054 521252 6060
rect 520832 3392 520884 3398
rect 520832 3334 520884 3340
rect 520280 3188 520332 3194
rect 520280 3130 520332 3136
rect 520292 480 520320 3130
rect 521212 3058 521240 6054
rect 521200 3052 521252 3058
rect 521200 2994 521252 3000
rect 521488 480 521516 6666
rect 522132 6186 522160 8092
rect 523236 6730 523264 8092
rect 523224 6724 523276 6730
rect 523224 6666 523276 6672
rect 524432 6662 524460 8092
rect 524512 6860 524564 6866
rect 524512 6802 524564 6808
rect 524420 6656 524472 6662
rect 524420 6598 524472 6604
rect 523868 6384 523920 6390
rect 523868 6326 523920 6332
rect 522120 6180 522172 6186
rect 522120 6122 522172 6128
rect 522822 6012 523386 6032
rect 522822 6010 522836 6012
rect 522892 6010 522916 6012
rect 522972 6010 522996 6012
rect 523052 6010 523076 6012
rect 523132 6010 523156 6012
rect 523212 6010 523236 6012
rect 523292 6010 523316 6012
rect 523372 6010 523386 6012
rect 523066 5958 523076 6010
rect 523132 5958 523142 6010
rect 522822 5956 522836 5958
rect 522892 5956 522916 5958
rect 522972 5956 522996 5958
rect 523052 5956 523076 5958
rect 523132 5956 523156 5958
rect 523212 5956 523236 5958
rect 523292 5956 523316 5958
rect 523372 5956 523386 5958
rect 522822 5936 523386 5956
rect 522396 5908 522448 5914
rect 522396 5850 522448 5856
rect 522408 2990 522436 5850
rect 522822 4924 523386 4944
rect 522822 4922 522836 4924
rect 522892 4922 522916 4924
rect 522972 4922 522996 4924
rect 523052 4922 523076 4924
rect 523132 4922 523156 4924
rect 523212 4922 523236 4924
rect 523292 4922 523316 4924
rect 523372 4922 523386 4924
rect 523066 4870 523076 4922
rect 523132 4870 523142 4922
rect 522822 4868 522836 4870
rect 522892 4868 522916 4870
rect 522972 4868 522996 4870
rect 523052 4868 523076 4870
rect 523132 4868 523156 4870
rect 523212 4868 523236 4870
rect 523292 4868 523316 4870
rect 523372 4868 523386 4870
rect 522822 4848 523386 4868
rect 522822 3836 523386 3856
rect 522822 3834 522836 3836
rect 522892 3834 522916 3836
rect 522972 3834 522996 3836
rect 523052 3834 523076 3836
rect 523132 3834 523156 3836
rect 523212 3834 523236 3836
rect 523292 3834 523316 3836
rect 523372 3834 523386 3836
rect 523066 3782 523076 3834
rect 523132 3782 523142 3834
rect 522822 3780 522836 3782
rect 522892 3780 522916 3782
rect 522972 3780 522996 3782
rect 523052 3780 523076 3782
rect 523132 3780 523156 3782
rect 523212 3780 523236 3782
rect 523292 3780 523316 3782
rect 523372 3780 523386 3782
rect 522822 3760 523386 3780
rect 522672 3392 522724 3398
rect 522672 3334 522724 3340
rect 522396 2984 522448 2990
rect 522396 2926 522448 2932
rect 522684 480 522712 3334
rect 522822 2748 523386 2768
rect 522822 2746 522836 2748
rect 522892 2746 522916 2748
rect 522972 2746 522996 2748
rect 523052 2746 523076 2748
rect 523132 2746 523156 2748
rect 523212 2746 523236 2748
rect 523292 2746 523316 2748
rect 523372 2746 523386 2748
rect 523066 2694 523076 2746
rect 523132 2694 523142 2746
rect 522822 2692 522836 2694
rect 522892 2692 522916 2694
rect 522972 2692 522996 2694
rect 523052 2692 523076 2694
rect 523132 2692 523156 2694
rect 523212 2692 523236 2694
rect 523292 2692 523316 2694
rect 523372 2692 523386 2694
rect 522822 2672 523386 2692
rect 523880 480 523908 6326
rect 524524 3738 524552 6802
rect 525064 6248 525116 6254
rect 525064 6190 525116 6196
rect 524512 3732 524564 3738
rect 524512 3674 524564 3680
rect 525076 480 525104 6190
rect 525536 3942 525564 8092
rect 525800 6792 525852 6798
rect 525800 6734 525852 6740
rect 525812 4010 525840 6734
rect 525800 4004 525852 4010
rect 525800 3946 525852 3952
rect 525524 3936 525576 3942
rect 525524 3878 525576 3884
rect 526640 3126 526668 8092
rect 527836 3534 527864 8092
rect 527824 3528 527876 3534
rect 527824 3470 527876 3476
rect 528652 3460 528704 3466
rect 528652 3402 528704 3408
rect 526628 3120 526680 3126
rect 526628 3062 526680 3068
rect 526260 3052 526312 3058
rect 526260 2994 526312 3000
rect 526272 480 526300 2994
rect 527456 2984 527508 2990
rect 527456 2926 527508 2932
rect 527468 480 527496 2926
rect 528664 480 528692 3402
rect 528940 2922 528968 8092
rect 530044 6254 530072 8092
rect 530032 6248 530084 6254
rect 530032 6190 530084 6196
rect 529848 5840 529900 5846
rect 529848 5782 529900 5788
rect 528928 2916 528980 2922
rect 528928 2858 528980 2864
rect 529860 480 529888 5782
rect 531240 3738 531268 8092
rect 532240 4004 532292 4010
rect 532240 3946 532292 3952
rect 531044 3732 531096 3738
rect 531044 3674 531096 3680
rect 531228 3732 531280 3738
rect 531228 3674 531280 3680
rect 531056 480 531084 3674
rect 532252 480 532280 3946
rect 532344 2854 532372 8092
rect 533344 6316 533396 6322
rect 533344 6258 533396 6264
rect 533356 3890 533384 6258
rect 533448 4010 533476 8092
rect 534540 6520 534592 6526
rect 534540 6462 534592 6468
rect 533436 4004 533488 4010
rect 533436 3946 533488 3952
rect 533356 3862 533476 3890
rect 532332 2848 532384 2854
rect 532332 2790 532384 2796
rect 533448 480 533476 3862
rect 534552 480 534580 6462
rect 534644 3466 534672 8092
rect 535748 4146 535776 8092
rect 536748 6656 536800 6662
rect 536748 6598 536800 6604
rect 535920 6588 535972 6594
rect 535920 6530 535972 6536
rect 535736 4140 535788 4146
rect 535736 4082 535788 4088
rect 535932 3942 535960 6530
rect 535920 3936 535972 3942
rect 535920 3878 535972 3884
rect 535736 3664 535788 3670
rect 535736 3606 535788 3612
rect 534632 3460 534684 3466
rect 534632 3402 534684 3408
rect 535748 480 535776 3606
rect 536760 2990 536788 6598
rect 536852 3058 536880 8092
rect 538048 3670 538076 8092
rect 538128 3936 538180 3942
rect 538128 3878 538180 3884
rect 538036 3664 538088 3670
rect 538036 3606 538088 3612
rect 536932 3596 536984 3602
rect 536932 3538 536984 3544
rect 536840 3052 536892 3058
rect 536840 2994 536892 3000
rect 536748 2984 536800 2990
rect 536748 2926 536800 2932
rect 536944 480 536972 3538
rect 538140 480 538168 3878
rect 539152 3466 539180 8092
rect 539324 6180 539376 6186
rect 539324 6122 539376 6128
rect 539140 3460 539192 3466
rect 539140 3402 539192 3408
rect 539336 480 539364 6122
rect 540256 3194 540284 8092
rect 541374 8078 541664 8106
rect 540520 6724 540572 6730
rect 540520 6666 540572 6672
rect 540244 3188 540296 3194
rect 540244 3130 540296 3136
rect 540532 480 540560 6666
rect 541440 6248 541492 6254
rect 541440 6190 541492 6196
rect 540822 5468 541386 5488
rect 540822 5466 540836 5468
rect 540892 5466 540916 5468
rect 540972 5466 540996 5468
rect 541052 5466 541076 5468
rect 541132 5466 541156 5468
rect 541212 5466 541236 5468
rect 541292 5466 541316 5468
rect 541372 5466 541386 5468
rect 541066 5414 541076 5466
rect 541132 5414 541142 5466
rect 540822 5412 540836 5414
rect 540892 5412 540916 5414
rect 540972 5412 540996 5414
rect 541052 5412 541076 5414
rect 541132 5412 541156 5414
rect 541212 5412 541236 5414
rect 541292 5412 541316 5414
rect 541372 5412 541386 5414
rect 540822 5392 541386 5412
rect 540822 4380 541386 4400
rect 540822 4378 540836 4380
rect 540892 4378 540916 4380
rect 540972 4378 540996 4380
rect 541052 4378 541076 4380
rect 541132 4378 541156 4380
rect 541212 4378 541236 4380
rect 541292 4378 541316 4380
rect 541372 4378 541386 4380
rect 541066 4326 541076 4378
rect 541132 4326 541142 4378
rect 540822 4324 540836 4326
rect 540892 4324 540916 4326
rect 540972 4324 540996 4326
rect 541052 4324 541076 4326
rect 541132 4324 541156 4326
rect 541212 4324 541236 4326
rect 541292 4324 541316 4326
rect 541372 4324 541386 4326
rect 540822 4304 541386 4324
rect 541452 4078 541480 6190
rect 541440 4072 541492 4078
rect 541440 4014 541492 4020
rect 541636 3942 541664 8078
rect 541624 3936 541676 3942
rect 541624 3878 541676 3884
rect 542556 3602 542584 8092
rect 542544 3596 542596 3602
rect 542544 3538 542596 3544
rect 543660 3398 543688 8092
rect 544764 3466 544792 8092
rect 545960 4078 545988 8092
rect 545948 4072 546000 4078
rect 545948 4014 546000 4020
rect 547064 3534 547092 8092
rect 547616 3602 547828 3618
rect 547616 3596 547840 3602
rect 547616 3590 547788 3596
rect 545304 3528 545356 3534
rect 545304 3470 545356 3476
rect 546592 3528 546644 3534
rect 546592 3470 546644 3476
rect 547052 3528 547104 3534
rect 547052 3470 547104 3476
rect 544752 3460 544804 3466
rect 544752 3402 544804 3408
rect 542912 3392 542964 3398
rect 542912 3334 542964 3340
rect 543648 3392 543700 3398
rect 543648 3334 543700 3340
rect 540822 3292 541386 3312
rect 540822 3290 540836 3292
rect 540892 3290 540916 3292
rect 540972 3290 540996 3292
rect 541052 3290 541076 3292
rect 541132 3290 541156 3292
rect 541212 3290 541236 3292
rect 541292 3290 541316 3292
rect 541372 3290 541386 3292
rect 541066 3238 541076 3290
rect 541132 3238 541142 3290
rect 540822 3236 540836 3238
rect 540892 3236 540916 3238
rect 540972 3236 540996 3238
rect 541052 3236 541076 3238
rect 541132 3236 541156 3238
rect 541212 3236 541236 3238
rect 541292 3236 541316 3238
rect 541372 3236 541386 3238
rect 540822 3216 541386 3236
rect 541716 2984 541768 2990
rect 541716 2926 541768 2932
rect 540822 2204 541386 2224
rect 540822 2202 540836 2204
rect 540892 2202 540916 2204
rect 540972 2202 540996 2204
rect 541052 2202 541076 2204
rect 541132 2202 541156 2204
rect 541212 2202 541236 2204
rect 541292 2202 541316 2204
rect 541372 2202 541386 2204
rect 541066 2150 541076 2202
rect 541132 2150 541142 2202
rect 540822 2148 540836 2150
rect 540892 2148 540916 2150
rect 540972 2148 540996 2150
rect 541052 2148 541076 2150
rect 541132 2148 541156 2150
rect 541212 2148 541236 2150
rect 541292 2148 541316 2150
rect 541372 2148 541386 2150
rect 540822 2128 541386 2148
rect 541728 480 541756 2926
rect 542924 480 542952 3334
rect 544108 3120 544160 3126
rect 544108 3062 544160 3068
rect 544120 480 544148 3062
rect 545316 480 545344 3470
rect 546604 2922 546632 3470
rect 547616 3466 547644 3590
rect 547788 3538 547840 3544
rect 547604 3460 547656 3466
rect 547604 3402 547656 3408
rect 547788 3392 547840 3398
rect 547788 3334 547840 3340
rect 547800 3210 547828 3334
rect 547708 3194 547828 3210
rect 547696 3188 547828 3194
rect 547748 3182 547828 3188
rect 547696 3130 547748 3136
rect 548168 2922 548196 8092
rect 549364 6118 549392 8092
rect 549352 6112 549404 6118
rect 549352 6054 549404 6060
rect 550468 3738 550496 8092
rect 550548 6112 550600 6118
rect 550548 6054 550600 6060
rect 548892 3732 548944 3738
rect 548892 3674 548944 3680
rect 550456 3732 550508 3738
rect 550456 3674 550508 3680
rect 546500 2916 546552 2922
rect 546500 2858 546552 2864
rect 546592 2916 546644 2922
rect 546592 2858 546644 2864
rect 547696 2916 547748 2922
rect 547696 2858 547748 2864
rect 548156 2916 548208 2922
rect 548156 2858 548208 2864
rect 546512 480 546540 2858
rect 547708 480 547736 2858
rect 548904 480 548932 3674
rect 550560 2854 550588 6054
rect 551572 4010 551600 8092
rect 551192 4004 551244 4010
rect 551192 3946 551244 3952
rect 551560 4004 551612 4010
rect 551560 3946 551612 3952
rect 550088 2848 550140 2854
rect 550088 2790 550140 2796
rect 550548 2848 550600 2854
rect 550548 2790 550600 2796
rect 550100 480 550128 2790
rect 551204 480 551232 3946
rect 552768 3738 552796 8092
rect 553872 4146 553900 8092
rect 553584 4140 553636 4146
rect 553584 4082 553636 4088
rect 553860 4140 553912 4146
rect 553860 4082 553912 4088
rect 552756 3732 552808 3738
rect 552756 3674 552808 3680
rect 552388 2984 552440 2990
rect 552388 2926 552440 2932
rect 552400 480 552428 2926
rect 553596 480 553624 4082
rect 554976 2990 555004 8092
rect 556172 3126 556200 8092
rect 557276 4146 557304 8092
rect 557264 4140 557316 4146
rect 557264 4082 557316 4088
rect 558380 3942 558408 8092
rect 558822 6012 559386 6032
rect 558822 6010 558836 6012
rect 558892 6010 558916 6012
rect 558972 6010 558996 6012
rect 559052 6010 559076 6012
rect 559132 6010 559156 6012
rect 559212 6010 559236 6012
rect 559292 6010 559316 6012
rect 559372 6010 559386 6012
rect 559066 5958 559076 6010
rect 559132 5958 559142 6010
rect 558822 5956 558836 5958
rect 558892 5956 558916 5958
rect 558972 5956 558996 5958
rect 559052 5956 559076 5958
rect 559132 5956 559156 5958
rect 559212 5956 559236 5958
rect 559292 5956 559316 5958
rect 559372 5956 559386 5958
rect 558822 5936 559386 5956
rect 558822 4924 559386 4944
rect 558822 4922 558836 4924
rect 558892 4922 558916 4924
rect 558972 4922 558996 4924
rect 559052 4922 559076 4924
rect 559132 4922 559156 4924
rect 559212 4922 559236 4924
rect 559292 4922 559316 4924
rect 559372 4922 559386 4924
rect 559066 4870 559076 4922
rect 559132 4870 559142 4922
rect 558822 4868 558836 4870
rect 558892 4868 558916 4870
rect 558972 4868 558996 4870
rect 559052 4868 559076 4870
rect 559132 4868 559156 4870
rect 559212 4868 559236 4870
rect 559292 4868 559316 4870
rect 559372 4868 559386 4870
rect 558822 4848 559386 4868
rect 558368 3936 558420 3942
rect 558368 3878 558420 3884
rect 558822 3836 559386 3856
rect 558822 3834 558836 3836
rect 558892 3834 558916 3836
rect 558972 3834 558996 3836
rect 559052 3834 559076 3836
rect 559132 3834 559156 3836
rect 559212 3834 559236 3836
rect 559292 3834 559316 3836
rect 559372 3834 559386 3836
rect 559066 3782 559076 3834
rect 559132 3782 559142 3834
rect 558822 3780 558836 3782
rect 558892 3780 558916 3782
rect 558972 3780 558996 3782
rect 559052 3780 559076 3782
rect 559132 3780 559156 3782
rect 559212 3780 559236 3782
rect 559292 3780 559316 3782
rect 559372 3780 559386 3782
rect 558822 3760 559386 3780
rect 559576 3670 559604 8092
rect 560680 4078 560708 8092
rect 560576 4072 560628 4078
rect 560576 4014 560628 4020
rect 560668 4072 560720 4078
rect 560668 4014 560720 4020
rect 560588 3890 560616 4014
rect 560588 3862 560800 3890
rect 559472 3664 559524 3670
rect 559472 3606 559524 3612
rect 559564 3664 559616 3670
rect 559564 3606 559616 3612
rect 559484 3482 559512 3606
rect 559484 3454 559604 3482
rect 558368 3392 558420 3398
rect 558368 3334 558420 3340
rect 557172 3188 557224 3194
rect 557172 3130 557224 3136
rect 555976 3120 556028 3126
rect 555976 3062 556028 3068
rect 556160 3120 556212 3126
rect 556160 3062 556212 3068
rect 554964 2984 555016 2990
rect 554964 2926 555016 2932
rect 554780 2644 554832 2650
rect 554780 2586 554832 2592
rect 554792 480 554820 2586
rect 555988 480 556016 3062
rect 557184 480 557212 3130
rect 558380 480 558408 3334
rect 558822 2748 559386 2768
rect 558822 2746 558836 2748
rect 558892 2746 558916 2748
rect 558972 2746 558996 2748
rect 559052 2746 559076 2748
rect 559132 2746 559156 2748
rect 559212 2746 559236 2748
rect 559292 2746 559316 2748
rect 559372 2746 559386 2748
rect 559066 2694 559076 2746
rect 559132 2694 559142 2746
rect 558822 2692 558836 2694
rect 558892 2692 558916 2694
rect 558972 2692 558996 2694
rect 559052 2692 559076 2694
rect 559132 2692 559156 2694
rect 559212 2692 559236 2694
rect 559292 2692 559316 2694
rect 559372 2692 559386 2694
rect 558822 2672 559386 2692
rect 559576 480 559604 3454
rect 560772 480 560800 3862
rect 561678 3496 561734 3505
rect 561784 3466 561812 8092
rect 562980 3942 563008 8092
rect 576822 5468 577386 5488
rect 576822 5466 576836 5468
rect 576892 5466 576916 5468
rect 576972 5466 576996 5468
rect 577052 5466 577076 5468
rect 577132 5466 577156 5468
rect 577212 5466 577236 5468
rect 577292 5466 577316 5468
rect 577372 5466 577386 5468
rect 577066 5414 577076 5466
rect 577132 5414 577142 5466
rect 576822 5412 576836 5414
rect 576892 5412 576916 5414
rect 576972 5412 576996 5414
rect 577052 5412 577076 5414
rect 577132 5412 577156 5414
rect 577212 5412 577236 5414
rect 577292 5412 577316 5414
rect 577372 5412 577386 5414
rect 576822 5392 577386 5412
rect 576822 4380 577386 4400
rect 576822 4378 576836 4380
rect 576892 4378 576916 4380
rect 576972 4378 576996 4380
rect 577052 4378 577076 4380
rect 577132 4378 577156 4380
rect 577212 4378 577236 4380
rect 577292 4378 577316 4380
rect 577372 4378 577386 4380
rect 577066 4326 577076 4378
rect 577132 4326 577142 4378
rect 576822 4324 576836 4326
rect 576892 4324 576916 4326
rect 576972 4324 576996 4326
rect 577052 4324 577076 4326
rect 577132 4324 577156 4326
rect 577212 4324 577236 4326
rect 577292 4324 577316 4326
rect 577372 4324 577386 4326
rect 576822 4304 577386 4324
rect 576216 4140 576268 4146
rect 576216 4082 576268 4088
rect 570236 4004 570288 4010
rect 570236 3946 570288 3952
rect 562968 3936 563020 3942
rect 562968 3878 563020 3884
rect 563152 3596 563204 3602
rect 563152 3538 563204 3544
rect 564532 3596 564584 3602
rect 564532 3538 564584 3544
rect 561678 3431 561680 3440
rect 561732 3431 561734 3440
rect 561772 3460 561824 3466
rect 561680 3402 561732 3408
rect 561772 3402 561824 3408
rect 561956 3392 562008 3398
rect 561956 3334 562008 3340
rect 561968 480 561996 3334
rect 563164 480 563192 3538
rect 564544 3505 564572 3538
rect 569040 3528 569092 3534
rect 564530 3496 564586 3505
rect 569040 3470 569092 3476
rect 564530 3431 564586 3440
rect 566740 3120 566792 3126
rect 566740 3062 566792 3068
rect 564348 2984 564400 2990
rect 564348 2926 564400 2932
rect 564360 480 564388 2926
rect 565544 2916 565596 2922
rect 565544 2858 565596 2864
rect 565556 480 565584 2858
rect 566752 480 566780 3062
rect 567844 2848 567896 2854
rect 567844 2790 567896 2796
rect 567856 480 567884 2790
rect 569052 480 569080 3470
rect 570248 480 570276 3946
rect 571432 3732 571484 3738
rect 571432 3674 571484 3680
rect 571444 480 571472 3674
rect 575020 3188 575072 3194
rect 575020 3130 575072 3136
rect 573824 3120 573876 3126
rect 573824 3062 573876 3068
rect 572628 2984 572680 2990
rect 572628 2926 572680 2932
rect 572640 480 572668 2926
rect 573836 480 573864 3062
rect 575032 480 575060 3130
rect 576228 480 576256 4082
rect 579804 4072 579856 4078
rect 579804 4014 579856 4020
rect 578608 3664 578660 3670
rect 578608 3606 578660 3612
rect 577412 3392 577464 3398
rect 577412 3334 577464 3340
rect 576822 3292 577386 3312
rect 576822 3290 576836 3292
rect 576892 3290 576916 3292
rect 576972 3290 576996 3292
rect 577052 3290 577076 3292
rect 577132 3290 577156 3292
rect 577212 3290 577236 3292
rect 577292 3290 577316 3292
rect 577372 3290 577386 3292
rect 577066 3238 577076 3290
rect 577132 3238 577142 3290
rect 576822 3236 576836 3238
rect 576892 3236 576916 3238
rect 576972 3236 576996 3238
rect 577052 3236 577076 3238
rect 577132 3236 577156 3238
rect 577212 3236 577236 3238
rect 577292 3236 577316 3238
rect 577372 3236 577386 3238
rect 576822 3216 577386 3236
rect 576822 2204 577386 2224
rect 576822 2202 576836 2204
rect 576892 2202 576916 2204
rect 576972 2202 576996 2204
rect 577052 2202 577076 2204
rect 577132 2202 577156 2204
rect 577212 2202 577236 2204
rect 577292 2202 577316 2204
rect 577372 2202 577386 2204
rect 577066 2150 577076 2202
rect 577132 2150 577142 2202
rect 576822 2148 576836 2150
rect 576892 2148 576916 2150
rect 576972 2148 576996 2150
rect 577052 2148 577076 2150
rect 577132 2148 577156 2150
rect 577212 2148 577236 2150
rect 577292 2148 577316 2150
rect 577372 2148 577386 2150
rect 576822 2128 577386 2148
rect 577424 480 577452 3334
rect 578620 480 578648 3606
rect 579816 480 579844 4014
rect 582196 3936 582248 3942
rect 582196 3878 582248 3884
rect 581000 3460 581052 3466
rect 581000 3402 581052 3408
rect 581012 480 581040 3402
rect 582208 480 582236 3878
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 18836 701242 18892 701244
rect 18916 701242 18972 701244
rect 18996 701242 19052 701244
rect 19076 701242 19132 701244
rect 19156 701242 19212 701244
rect 19236 701242 19292 701244
rect 19316 701242 19372 701244
rect 18836 701190 18874 701242
rect 18874 701190 18886 701242
rect 18886 701190 18892 701242
rect 18916 701190 18938 701242
rect 18938 701190 18950 701242
rect 18950 701190 18972 701242
rect 18996 701190 19002 701242
rect 19002 701190 19014 701242
rect 19014 701190 19052 701242
rect 19076 701190 19078 701242
rect 19078 701190 19130 701242
rect 19130 701190 19132 701242
rect 19156 701190 19194 701242
rect 19194 701190 19206 701242
rect 19206 701190 19212 701242
rect 19236 701190 19258 701242
rect 19258 701190 19270 701242
rect 19270 701190 19292 701242
rect 19316 701190 19322 701242
rect 19322 701190 19334 701242
rect 19334 701190 19372 701242
rect 18836 701188 18892 701190
rect 18916 701188 18972 701190
rect 18996 701188 19052 701190
rect 19076 701188 19132 701190
rect 19156 701188 19212 701190
rect 19236 701188 19292 701190
rect 19316 701188 19372 701190
rect 36836 701786 36892 701788
rect 36916 701786 36972 701788
rect 36996 701786 37052 701788
rect 37076 701786 37132 701788
rect 37156 701786 37212 701788
rect 37236 701786 37292 701788
rect 37316 701786 37372 701788
rect 36836 701734 36874 701786
rect 36874 701734 36886 701786
rect 36886 701734 36892 701786
rect 36916 701734 36938 701786
rect 36938 701734 36950 701786
rect 36950 701734 36972 701786
rect 36996 701734 37002 701786
rect 37002 701734 37014 701786
rect 37014 701734 37052 701786
rect 37076 701734 37078 701786
rect 37078 701734 37130 701786
rect 37130 701734 37132 701786
rect 37156 701734 37194 701786
rect 37194 701734 37206 701786
rect 37206 701734 37212 701786
rect 37236 701734 37258 701786
rect 37258 701734 37270 701786
rect 37270 701734 37292 701786
rect 37316 701734 37322 701786
rect 37322 701734 37334 701786
rect 37334 701734 37372 701786
rect 36836 701732 36892 701734
rect 36916 701732 36972 701734
rect 36996 701732 37052 701734
rect 37076 701732 37132 701734
rect 37156 701732 37212 701734
rect 37236 701732 37292 701734
rect 37316 701732 37372 701734
rect 54836 701242 54892 701244
rect 54916 701242 54972 701244
rect 54996 701242 55052 701244
rect 55076 701242 55132 701244
rect 55156 701242 55212 701244
rect 55236 701242 55292 701244
rect 55316 701242 55372 701244
rect 54836 701190 54874 701242
rect 54874 701190 54886 701242
rect 54886 701190 54892 701242
rect 54916 701190 54938 701242
rect 54938 701190 54950 701242
rect 54950 701190 54972 701242
rect 54996 701190 55002 701242
rect 55002 701190 55014 701242
rect 55014 701190 55052 701242
rect 55076 701190 55078 701242
rect 55078 701190 55130 701242
rect 55130 701190 55132 701242
rect 55156 701190 55194 701242
rect 55194 701190 55206 701242
rect 55206 701190 55212 701242
rect 55236 701190 55258 701242
rect 55258 701190 55270 701242
rect 55270 701190 55292 701242
rect 55316 701190 55322 701242
rect 55322 701190 55334 701242
rect 55334 701190 55372 701242
rect 54836 701188 54892 701190
rect 54916 701188 54972 701190
rect 54996 701188 55052 701190
rect 55076 701188 55132 701190
rect 55156 701188 55212 701190
rect 55236 701188 55292 701190
rect 55316 701188 55372 701190
rect 40498 700984 40554 701040
rect 36836 700698 36892 700700
rect 36916 700698 36972 700700
rect 36996 700698 37052 700700
rect 37076 700698 37132 700700
rect 37156 700698 37212 700700
rect 37236 700698 37292 700700
rect 37316 700698 37372 700700
rect 36836 700646 36874 700698
rect 36874 700646 36886 700698
rect 36886 700646 36892 700698
rect 36916 700646 36938 700698
rect 36938 700646 36950 700698
rect 36950 700646 36972 700698
rect 36996 700646 37002 700698
rect 37002 700646 37014 700698
rect 37014 700646 37052 700698
rect 37076 700646 37078 700698
rect 37078 700646 37130 700698
rect 37130 700646 37132 700698
rect 37156 700646 37194 700698
rect 37194 700646 37206 700698
rect 37206 700646 37212 700698
rect 37236 700646 37258 700698
rect 37258 700646 37270 700698
rect 37270 700646 37292 700698
rect 37316 700646 37322 700698
rect 37322 700646 37334 700698
rect 37334 700646 37372 700698
rect 36836 700644 36892 700646
rect 36916 700644 36972 700646
rect 36996 700644 37052 700646
rect 37076 700644 37132 700646
rect 37156 700644 37212 700646
rect 37236 700644 37292 700646
rect 37316 700644 37372 700646
rect 24306 700440 24362 700496
rect 8114 700304 8170 700360
rect 72836 701786 72892 701788
rect 72916 701786 72972 701788
rect 72996 701786 73052 701788
rect 73076 701786 73132 701788
rect 73156 701786 73212 701788
rect 73236 701786 73292 701788
rect 73316 701786 73372 701788
rect 72836 701734 72874 701786
rect 72874 701734 72886 701786
rect 72886 701734 72892 701786
rect 72916 701734 72938 701786
rect 72938 701734 72950 701786
rect 72950 701734 72972 701786
rect 72996 701734 73002 701786
rect 73002 701734 73014 701786
rect 73014 701734 73052 701786
rect 73076 701734 73078 701786
rect 73078 701734 73130 701786
rect 73130 701734 73132 701786
rect 73156 701734 73194 701786
rect 73194 701734 73206 701786
rect 73206 701734 73212 701786
rect 73236 701734 73258 701786
rect 73258 701734 73270 701786
rect 73270 701734 73292 701786
rect 73316 701734 73322 701786
rect 73322 701734 73334 701786
rect 73334 701734 73372 701786
rect 72836 701732 72892 701734
rect 72916 701732 72972 701734
rect 72996 701732 73052 701734
rect 73076 701732 73132 701734
rect 73156 701732 73212 701734
rect 73236 701732 73292 701734
rect 73316 701732 73372 701734
rect 72836 700698 72892 700700
rect 72916 700698 72972 700700
rect 72996 700698 73052 700700
rect 73076 700698 73132 700700
rect 73156 700698 73212 700700
rect 73236 700698 73292 700700
rect 73316 700698 73372 700700
rect 72836 700646 72874 700698
rect 72874 700646 72886 700698
rect 72886 700646 72892 700698
rect 72916 700646 72938 700698
rect 72938 700646 72950 700698
rect 72950 700646 72972 700698
rect 72996 700646 73002 700698
rect 73002 700646 73014 700698
rect 73014 700646 73052 700698
rect 73076 700646 73078 700698
rect 73078 700646 73130 700698
rect 73130 700646 73132 700698
rect 73156 700646 73194 700698
rect 73194 700646 73206 700698
rect 73206 700646 73212 700698
rect 73236 700646 73258 700698
rect 73258 700646 73270 700698
rect 73270 700646 73292 700698
rect 73316 700646 73322 700698
rect 73322 700646 73334 700698
rect 73334 700646 73372 700698
rect 72836 700644 72892 700646
rect 72916 700644 72972 700646
rect 72996 700644 73052 700646
rect 73076 700644 73132 700646
rect 73156 700644 73212 700646
rect 73236 700644 73292 700646
rect 73316 700644 73372 700646
rect 90836 701242 90892 701244
rect 90916 701242 90972 701244
rect 90996 701242 91052 701244
rect 91076 701242 91132 701244
rect 91156 701242 91212 701244
rect 91236 701242 91292 701244
rect 91316 701242 91372 701244
rect 90836 701190 90874 701242
rect 90874 701190 90886 701242
rect 90886 701190 90892 701242
rect 90916 701190 90938 701242
rect 90938 701190 90950 701242
rect 90950 701190 90972 701242
rect 90996 701190 91002 701242
rect 91002 701190 91014 701242
rect 91014 701190 91052 701242
rect 91076 701190 91078 701242
rect 91078 701190 91130 701242
rect 91130 701190 91132 701242
rect 91156 701190 91194 701242
rect 91194 701190 91206 701242
rect 91206 701190 91212 701242
rect 91236 701190 91258 701242
rect 91258 701190 91270 701242
rect 91270 701190 91292 701242
rect 91316 701190 91322 701242
rect 91322 701190 91334 701242
rect 91334 701190 91372 701242
rect 90836 701188 90892 701190
rect 90916 701188 90972 701190
rect 90996 701188 91052 701190
rect 91076 701188 91132 701190
rect 91156 701188 91212 701190
rect 91236 701188 91292 701190
rect 91316 701188 91372 701190
rect 108836 701786 108892 701788
rect 108916 701786 108972 701788
rect 108996 701786 109052 701788
rect 109076 701786 109132 701788
rect 109156 701786 109212 701788
rect 109236 701786 109292 701788
rect 109316 701786 109372 701788
rect 108836 701734 108874 701786
rect 108874 701734 108886 701786
rect 108886 701734 108892 701786
rect 108916 701734 108938 701786
rect 108938 701734 108950 701786
rect 108950 701734 108972 701786
rect 108996 701734 109002 701786
rect 109002 701734 109014 701786
rect 109014 701734 109052 701786
rect 109076 701734 109078 701786
rect 109078 701734 109130 701786
rect 109130 701734 109132 701786
rect 109156 701734 109194 701786
rect 109194 701734 109206 701786
rect 109206 701734 109212 701786
rect 109236 701734 109258 701786
rect 109258 701734 109270 701786
rect 109270 701734 109292 701786
rect 109316 701734 109322 701786
rect 109322 701734 109334 701786
rect 109334 701734 109372 701786
rect 108836 701732 108892 701734
rect 108916 701732 108972 701734
rect 108996 701732 109052 701734
rect 109076 701732 109132 701734
rect 109156 701732 109212 701734
rect 109236 701732 109292 701734
rect 109316 701732 109372 701734
rect 126836 701242 126892 701244
rect 126916 701242 126972 701244
rect 126996 701242 127052 701244
rect 127076 701242 127132 701244
rect 127156 701242 127212 701244
rect 127236 701242 127292 701244
rect 127316 701242 127372 701244
rect 126836 701190 126874 701242
rect 126874 701190 126886 701242
rect 126886 701190 126892 701242
rect 126916 701190 126938 701242
rect 126938 701190 126950 701242
rect 126950 701190 126972 701242
rect 126996 701190 127002 701242
rect 127002 701190 127014 701242
rect 127014 701190 127052 701242
rect 127076 701190 127078 701242
rect 127078 701190 127130 701242
rect 127130 701190 127132 701242
rect 127156 701190 127194 701242
rect 127194 701190 127206 701242
rect 127206 701190 127212 701242
rect 127236 701190 127258 701242
rect 127258 701190 127270 701242
rect 127270 701190 127292 701242
rect 127316 701190 127322 701242
rect 127322 701190 127334 701242
rect 127334 701190 127372 701242
rect 126836 701188 126892 701190
rect 126916 701188 126972 701190
rect 126996 701188 127052 701190
rect 127076 701188 127132 701190
rect 127156 701188 127212 701190
rect 127236 701188 127292 701190
rect 127316 701188 127372 701190
rect 144836 701786 144892 701788
rect 144916 701786 144972 701788
rect 144996 701786 145052 701788
rect 145076 701786 145132 701788
rect 145156 701786 145212 701788
rect 145236 701786 145292 701788
rect 145316 701786 145372 701788
rect 144836 701734 144874 701786
rect 144874 701734 144886 701786
rect 144886 701734 144892 701786
rect 144916 701734 144938 701786
rect 144938 701734 144950 701786
rect 144950 701734 144972 701786
rect 144996 701734 145002 701786
rect 145002 701734 145014 701786
rect 145014 701734 145052 701786
rect 145076 701734 145078 701786
rect 145078 701734 145130 701786
rect 145130 701734 145132 701786
rect 145156 701734 145194 701786
rect 145194 701734 145206 701786
rect 145206 701734 145212 701786
rect 145236 701734 145258 701786
rect 145258 701734 145270 701786
rect 145270 701734 145292 701786
rect 145316 701734 145322 701786
rect 145322 701734 145334 701786
rect 145334 701734 145372 701786
rect 144836 701732 144892 701734
rect 144916 701732 144972 701734
rect 144996 701732 145052 701734
rect 145076 701732 145132 701734
rect 145156 701732 145212 701734
rect 145236 701732 145292 701734
rect 145316 701732 145372 701734
rect 162836 701242 162892 701244
rect 162916 701242 162972 701244
rect 162996 701242 163052 701244
rect 163076 701242 163132 701244
rect 163156 701242 163212 701244
rect 163236 701242 163292 701244
rect 163316 701242 163372 701244
rect 162836 701190 162874 701242
rect 162874 701190 162886 701242
rect 162886 701190 162892 701242
rect 162916 701190 162938 701242
rect 162938 701190 162950 701242
rect 162950 701190 162972 701242
rect 162996 701190 163002 701242
rect 163002 701190 163014 701242
rect 163014 701190 163052 701242
rect 163076 701190 163078 701242
rect 163078 701190 163130 701242
rect 163130 701190 163132 701242
rect 163156 701190 163194 701242
rect 163194 701190 163206 701242
rect 163206 701190 163212 701242
rect 163236 701190 163258 701242
rect 163258 701190 163270 701242
rect 163270 701190 163292 701242
rect 163316 701190 163322 701242
rect 163322 701190 163334 701242
rect 163334 701190 163372 701242
rect 162836 701188 162892 701190
rect 162916 701188 162972 701190
rect 162996 701188 163052 701190
rect 163076 701188 163132 701190
rect 163156 701188 163212 701190
rect 163236 701188 163292 701190
rect 163316 701188 163372 701190
rect 108836 700698 108892 700700
rect 108916 700698 108972 700700
rect 108996 700698 109052 700700
rect 109076 700698 109132 700700
rect 109156 700698 109212 700700
rect 109236 700698 109292 700700
rect 109316 700698 109372 700700
rect 108836 700646 108874 700698
rect 108874 700646 108886 700698
rect 108886 700646 108892 700698
rect 108916 700646 108938 700698
rect 108938 700646 108950 700698
rect 108950 700646 108972 700698
rect 108996 700646 109002 700698
rect 109002 700646 109014 700698
rect 109014 700646 109052 700698
rect 109076 700646 109078 700698
rect 109078 700646 109130 700698
rect 109130 700646 109132 700698
rect 109156 700646 109194 700698
rect 109194 700646 109206 700698
rect 109206 700646 109212 700698
rect 109236 700646 109258 700698
rect 109258 700646 109270 700698
rect 109270 700646 109292 700698
rect 109316 700646 109322 700698
rect 109322 700646 109334 700698
rect 109334 700646 109372 700698
rect 108836 700644 108892 700646
rect 108916 700644 108972 700646
rect 108996 700644 109052 700646
rect 109076 700644 109132 700646
rect 109156 700644 109212 700646
rect 109236 700644 109292 700646
rect 109316 700644 109372 700646
rect 144836 700698 144892 700700
rect 144916 700698 144972 700700
rect 144996 700698 145052 700700
rect 145076 700698 145132 700700
rect 145156 700698 145212 700700
rect 145236 700698 145292 700700
rect 145316 700698 145372 700700
rect 144836 700646 144874 700698
rect 144874 700646 144886 700698
rect 144886 700646 144892 700698
rect 144916 700646 144938 700698
rect 144938 700646 144950 700698
rect 144950 700646 144972 700698
rect 144996 700646 145002 700698
rect 145002 700646 145014 700698
rect 145014 700646 145052 700698
rect 145076 700646 145078 700698
rect 145078 700646 145130 700698
rect 145130 700646 145132 700698
rect 145156 700646 145194 700698
rect 145194 700646 145206 700698
rect 145206 700646 145212 700698
rect 145236 700646 145258 700698
rect 145258 700646 145270 700698
rect 145270 700646 145292 700698
rect 145316 700646 145322 700698
rect 145322 700646 145334 700698
rect 145334 700646 145372 700698
rect 144836 700644 144892 700646
rect 144916 700644 144972 700646
rect 144996 700644 145052 700646
rect 145076 700644 145132 700646
rect 145156 700644 145212 700646
rect 145236 700644 145292 700646
rect 145316 700644 145372 700646
rect 18836 700154 18892 700156
rect 18916 700154 18972 700156
rect 18996 700154 19052 700156
rect 19076 700154 19132 700156
rect 19156 700154 19212 700156
rect 19236 700154 19292 700156
rect 19316 700154 19372 700156
rect 18836 700102 18874 700154
rect 18874 700102 18886 700154
rect 18886 700102 18892 700154
rect 18916 700102 18938 700154
rect 18938 700102 18950 700154
rect 18950 700102 18972 700154
rect 18996 700102 19002 700154
rect 19002 700102 19014 700154
rect 19014 700102 19052 700154
rect 19076 700102 19078 700154
rect 19078 700102 19130 700154
rect 19130 700102 19132 700154
rect 19156 700102 19194 700154
rect 19194 700102 19206 700154
rect 19206 700102 19212 700154
rect 19236 700102 19258 700154
rect 19258 700102 19270 700154
rect 19270 700102 19292 700154
rect 19316 700102 19322 700154
rect 19322 700102 19334 700154
rect 19334 700102 19372 700154
rect 18836 700100 18892 700102
rect 18916 700100 18972 700102
rect 18996 700100 19052 700102
rect 19076 700100 19132 700102
rect 19156 700100 19212 700102
rect 19236 700100 19292 700102
rect 19316 700100 19372 700102
rect 54836 700154 54892 700156
rect 54916 700154 54972 700156
rect 54996 700154 55052 700156
rect 55076 700154 55132 700156
rect 55156 700154 55212 700156
rect 55236 700154 55292 700156
rect 55316 700154 55372 700156
rect 54836 700102 54874 700154
rect 54874 700102 54886 700154
rect 54886 700102 54892 700154
rect 54916 700102 54938 700154
rect 54938 700102 54950 700154
rect 54950 700102 54972 700154
rect 54996 700102 55002 700154
rect 55002 700102 55014 700154
rect 55014 700102 55052 700154
rect 55076 700102 55078 700154
rect 55078 700102 55130 700154
rect 55130 700102 55132 700154
rect 55156 700102 55194 700154
rect 55194 700102 55206 700154
rect 55206 700102 55212 700154
rect 55236 700102 55258 700154
rect 55258 700102 55270 700154
rect 55270 700102 55292 700154
rect 55316 700102 55322 700154
rect 55322 700102 55334 700154
rect 55334 700102 55372 700154
rect 54836 700100 54892 700102
rect 54916 700100 54972 700102
rect 54996 700100 55052 700102
rect 55076 700100 55132 700102
rect 55156 700100 55212 700102
rect 55236 700100 55292 700102
rect 55316 700100 55372 700102
rect 90836 700154 90892 700156
rect 90916 700154 90972 700156
rect 90996 700154 91052 700156
rect 91076 700154 91132 700156
rect 91156 700154 91212 700156
rect 91236 700154 91292 700156
rect 91316 700154 91372 700156
rect 90836 700102 90874 700154
rect 90874 700102 90886 700154
rect 90886 700102 90892 700154
rect 90916 700102 90938 700154
rect 90938 700102 90950 700154
rect 90950 700102 90972 700154
rect 90996 700102 91002 700154
rect 91002 700102 91014 700154
rect 91014 700102 91052 700154
rect 91076 700102 91078 700154
rect 91078 700102 91130 700154
rect 91130 700102 91132 700154
rect 91156 700102 91194 700154
rect 91194 700102 91206 700154
rect 91206 700102 91212 700154
rect 91236 700102 91258 700154
rect 91258 700102 91270 700154
rect 91270 700102 91292 700154
rect 91316 700102 91322 700154
rect 91322 700102 91334 700154
rect 91334 700102 91372 700154
rect 90836 700100 90892 700102
rect 90916 700100 90972 700102
rect 90996 700100 91052 700102
rect 91076 700100 91132 700102
rect 91156 700100 91212 700102
rect 91236 700100 91292 700102
rect 91316 700100 91372 700102
rect 126836 700154 126892 700156
rect 126916 700154 126972 700156
rect 126996 700154 127052 700156
rect 127076 700154 127132 700156
rect 127156 700154 127212 700156
rect 127236 700154 127292 700156
rect 127316 700154 127372 700156
rect 126836 700102 126874 700154
rect 126874 700102 126886 700154
rect 126886 700102 126892 700154
rect 126916 700102 126938 700154
rect 126938 700102 126950 700154
rect 126950 700102 126972 700154
rect 126996 700102 127002 700154
rect 127002 700102 127014 700154
rect 127014 700102 127052 700154
rect 127076 700102 127078 700154
rect 127078 700102 127130 700154
rect 127130 700102 127132 700154
rect 127156 700102 127194 700154
rect 127194 700102 127206 700154
rect 127206 700102 127212 700154
rect 127236 700102 127258 700154
rect 127258 700102 127270 700154
rect 127270 700102 127292 700154
rect 127316 700102 127322 700154
rect 127322 700102 127334 700154
rect 127334 700102 127372 700154
rect 126836 700100 126892 700102
rect 126916 700100 126972 700102
rect 126996 700100 127052 700102
rect 127076 700100 127132 700102
rect 127156 700100 127212 700102
rect 127236 700100 127292 700102
rect 127316 700100 127372 700102
rect 162836 700154 162892 700156
rect 162916 700154 162972 700156
rect 162996 700154 163052 700156
rect 163076 700154 163132 700156
rect 163156 700154 163212 700156
rect 163236 700154 163292 700156
rect 163316 700154 163372 700156
rect 162836 700102 162874 700154
rect 162874 700102 162886 700154
rect 162886 700102 162892 700154
rect 162916 700102 162938 700154
rect 162938 700102 162950 700154
rect 162950 700102 162972 700154
rect 162996 700102 163002 700154
rect 163002 700102 163014 700154
rect 163014 700102 163052 700154
rect 163076 700102 163078 700154
rect 163078 700102 163130 700154
rect 163130 700102 163132 700154
rect 163156 700102 163194 700154
rect 163194 700102 163206 700154
rect 163206 700102 163212 700154
rect 163236 700102 163258 700154
rect 163258 700102 163270 700154
rect 163270 700102 163292 700154
rect 163316 700102 163322 700154
rect 163322 700102 163334 700154
rect 163334 700102 163372 700154
rect 162836 700100 162892 700102
rect 162916 700100 162972 700102
rect 162996 700100 163052 700102
rect 163076 700100 163132 700102
rect 163156 700100 163212 700102
rect 163236 700100 163292 700102
rect 163316 700100 163372 700102
rect 180836 701786 180892 701788
rect 180916 701786 180972 701788
rect 180996 701786 181052 701788
rect 181076 701786 181132 701788
rect 181156 701786 181212 701788
rect 181236 701786 181292 701788
rect 181316 701786 181372 701788
rect 180836 701734 180874 701786
rect 180874 701734 180886 701786
rect 180886 701734 180892 701786
rect 180916 701734 180938 701786
rect 180938 701734 180950 701786
rect 180950 701734 180972 701786
rect 180996 701734 181002 701786
rect 181002 701734 181014 701786
rect 181014 701734 181052 701786
rect 181076 701734 181078 701786
rect 181078 701734 181130 701786
rect 181130 701734 181132 701786
rect 181156 701734 181194 701786
rect 181194 701734 181206 701786
rect 181206 701734 181212 701786
rect 181236 701734 181258 701786
rect 181258 701734 181270 701786
rect 181270 701734 181292 701786
rect 181316 701734 181322 701786
rect 181322 701734 181334 701786
rect 181334 701734 181372 701786
rect 180836 701732 180892 701734
rect 180916 701732 180972 701734
rect 180996 701732 181052 701734
rect 181076 701732 181132 701734
rect 181156 701732 181212 701734
rect 181236 701732 181292 701734
rect 181316 701732 181372 701734
rect 198836 701242 198892 701244
rect 198916 701242 198972 701244
rect 198996 701242 199052 701244
rect 199076 701242 199132 701244
rect 199156 701242 199212 701244
rect 199236 701242 199292 701244
rect 199316 701242 199372 701244
rect 198836 701190 198874 701242
rect 198874 701190 198886 701242
rect 198886 701190 198892 701242
rect 198916 701190 198938 701242
rect 198938 701190 198950 701242
rect 198950 701190 198972 701242
rect 198996 701190 199002 701242
rect 199002 701190 199014 701242
rect 199014 701190 199052 701242
rect 199076 701190 199078 701242
rect 199078 701190 199130 701242
rect 199130 701190 199132 701242
rect 199156 701190 199194 701242
rect 199194 701190 199206 701242
rect 199206 701190 199212 701242
rect 199236 701190 199258 701242
rect 199258 701190 199270 701242
rect 199270 701190 199292 701242
rect 199316 701190 199322 701242
rect 199322 701190 199334 701242
rect 199334 701190 199372 701242
rect 198836 701188 198892 701190
rect 198916 701188 198972 701190
rect 198996 701188 199052 701190
rect 199076 701188 199132 701190
rect 199156 701188 199212 701190
rect 199236 701188 199292 701190
rect 199316 701188 199372 701190
rect 180836 700698 180892 700700
rect 180916 700698 180972 700700
rect 180996 700698 181052 700700
rect 181076 700698 181132 700700
rect 181156 700698 181212 700700
rect 181236 700698 181292 700700
rect 181316 700698 181372 700700
rect 180836 700646 180874 700698
rect 180874 700646 180886 700698
rect 180886 700646 180892 700698
rect 180916 700646 180938 700698
rect 180938 700646 180950 700698
rect 180950 700646 180972 700698
rect 180996 700646 181002 700698
rect 181002 700646 181014 700698
rect 181014 700646 181052 700698
rect 181076 700646 181078 700698
rect 181078 700646 181130 700698
rect 181130 700646 181132 700698
rect 181156 700646 181194 700698
rect 181194 700646 181206 700698
rect 181206 700646 181212 700698
rect 181236 700646 181258 700698
rect 181258 700646 181270 700698
rect 181270 700646 181292 700698
rect 181316 700646 181322 700698
rect 181322 700646 181334 700698
rect 181334 700646 181372 700698
rect 180836 700644 180892 700646
rect 180916 700644 180972 700646
rect 180996 700644 181052 700646
rect 181076 700644 181132 700646
rect 181156 700644 181212 700646
rect 181236 700644 181292 700646
rect 181316 700644 181372 700646
rect 216836 701786 216892 701788
rect 216916 701786 216972 701788
rect 216996 701786 217052 701788
rect 217076 701786 217132 701788
rect 217156 701786 217212 701788
rect 217236 701786 217292 701788
rect 217316 701786 217372 701788
rect 216836 701734 216874 701786
rect 216874 701734 216886 701786
rect 216886 701734 216892 701786
rect 216916 701734 216938 701786
rect 216938 701734 216950 701786
rect 216950 701734 216972 701786
rect 216996 701734 217002 701786
rect 217002 701734 217014 701786
rect 217014 701734 217052 701786
rect 217076 701734 217078 701786
rect 217078 701734 217130 701786
rect 217130 701734 217132 701786
rect 217156 701734 217194 701786
rect 217194 701734 217206 701786
rect 217206 701734 217212 701786
rect 217236 701734 217258 701786
rect 217258 701734 217270 701786
rect 217270 701734 217292 701786
rect 217316 701734 217322 701786
rect 217322 701734 217334 701786
rect 217334 701734 217372 701786
rect 216836 701732 216892 701734
rect 216916 701732 216972 701734
rect 216996 701732 217052 701734
rect 217076 701732 217132 701734
rect 217156 701732 217212 701734
rect 217236 701732 217292 701734
rect 217316 701732 217372 701734
rect 216836 700698 216892 700700
rect 216916 700698 216972 700700
rect 216996 700698 217052 700700
rect 217076 700698 217132 700700
rect 217156 700698 217212 700700
rect 217236 700698 217292 700700
rect 217316 700698 217372 700700
rect 216836 700646 216874 700698
rect 216874 700646 216886 700698
rect 216886 700646 216892 700698
rect 216916 700646 216938 700698
rect 216938 700646 216950 700698
rect 216950 700646 216972 700698
rect 216996 700646 217002 700698
rect 217002 700646 217014 700698
rect 217014 700646 217052 700698
rect 217076 700646 217078 700698
rect 217078 700646 217130 700698
rect 217130 700646 217132 700698
rect 217156 700646 217194 700698
rect 217194 700646 217206 700698
rect 217206 700646 217212 700698
rect 217236 700646 217258 700698
rect 217258 700646 217270 700698
rect 217270 700646 217292 700698
rect 217316 700646 217322 700698
rect 217322 700646 217334 700698
rect 217334 700646 217372 700698
rect 216836 700644 216892 700646
rect 216916 700644 216972 700646
rect 216996 700644 217052 700646
rect 217076 700644 217132 700646
rect 217156 700644 217212 700646
rect 217236 700644 217292 700646
rect 217316 700644 217372 700646
rect 198836 700154 198892 700156
rect 198916 700154 198972 700156
rect 198996 700154 199052 700156
rect 199076 700154 199132 700156
rect 199156 700154 199212 700156
rect 199236 700154 199292 700156
rect 199316 700154 199372 700156
rect 198836 700102 198874 700154
rect 198874 700102 198886 700154
rect 198886 700102 198892 700154
rect 198916 700102 198938 700154
rect 198938 700102 198950 700154
rect 198950 700102 198972 700154
rect 198996 700102 199002 700154
rect 199002 700102 199014 700154
rect 199014 700102 199052 700154
rect 199076 700102 199078 700154
rect 199078 700102 199130 700154
rect 199130 700102 199132 700154
rect 199156 700102 199194 700154
rect 199194 700102 199206 700154
rect 199206 700102 199212 700154
rect 199236 700102 199258 700154
rect 199258 700102 199270 700154
rect 199270 700102 199292 700154
rect 199316 700102 199322 700154
rect 199322 700102 199334 700154
rect 199334 700102 199372 700154
rect 198836 700100 198892 700102
rect 198916 700100 198972 700102
rect 198996 700100 199052 700102
rect 199076 700100 199132 700102
rect 199156 700100 199212 700102
rect 199236 700100 199292 700102
rect 199316 700100 199372 700102
rect 36836 699610 36892 699612
rect 36916 699610 36972 699612
rect 36996 699610 37052 699612
rect 37076 699610 37132 699612
rect 37156 699610 37212 699612
rect 37236 699610 37292 699612
rect 37316 699610 37372 699612
rect 36836 699558 36874 699610
rect 36874 699558 36886 699610
rect 36886 699558 36892 699610
rect 36916 699558 36938 699610
rect 36938 699558 36950 699610
rect 36950 699558 36972 699610
rect 36996 699558 37002 699610
rect 37002 699558 37014 699610
rect 37014 699558 37052 699610
rect 37076 699558 37078 699610
rect 37078 699558 37130 699610
rect 37130 699558 37132 699610
rect 37156 699558 37194 699610
rect 37194 699558 37206 699610
rect 37206 699558 37212 699610
rect 37236 699558 37258 699610
rect 37258 699558 37270 699610
rect 37270 699558 37292 699610
rect 37316 699558 37322 699610
rect 37322 699558 37334 699610
rect 37334 699558 37372 699610
rect 36836 699556 36892 699558
rect 36916 699556 36972 699558
rect 36996 699556 37052 699558
rect 37076 699556 37132 699558
rect 37156 699556 37212 699558
rect 37236 699556 37292 699558
rect 37316 699556 37372 699558
rect 72836 699610 72892 699612
rect 72916 699610 72972 699612
rect 72996 699610 73052 699612
rect 73076 699610 73132 699612
rect 73156 699610 73212 699612
rect 73236 699610 73292 699612
rect 73316 699610 73372 699612
rect 72836 699558 72874 699610
rect 72874 699558 72886 699610
rect 72886 699558 72892 699610
rect 72916 699558 72938 699610
rect 72938 699558 72950 699610
rect 72950 699558 72972 699610
rect 72996 699558 73002 699610
rect 73002 699558 73014 699610
rect 73014 699558 73052 699610
rect 73076 699558 73078 699610
rect 73078 699558 73130 699610
rect 73130 699558 73132 699610
rect 73156 699558 73194 699610
rect 73194 699558 73206 699610
rect 73206 699558 73212 699610
rect 73236 699558 73258 699610
rect 73258 699558 73270 699610
rect 73270 699558 73292 699610
rect 73316 699558 73322 699610
rect 73322 699558 73334 699610
rect 73334 699558 73372 699610
rect 72836 699556 72892 699558
rect 72916 699556 72972 699558
rect 72996 699556 73052 699558
rect 73076 699556 73132 699558
rect 73156 699556 73212 699558
rect 73236 699556 73292 699558
rect 73316 699556 73372 699558
rect 108836 699610 108892 699612
rect 108916 699610 108972 699612
rect 108996 699610 109052 699612
rect 109076 699610 109132 699612
rect 109156 699610 109212 699612
rect 109236 699610 109292 699612
rect 109316 699610 109372 699612
rect 108836 699558 108874 699610
rect 108874 699558 108886 699610
rect 108886 699558 108892 699610
rect 108916 699558 108938 699610
rect 108938 699558 108950 699610
rect 108950 699558 108972 699610
rect 108996 699558 109002 699610
rect 109002 699558 109014 699610
rect 109014 699558 109052 699610
rect 109076 699558 109078 699610
rect 109078 699558 109130 699610
rect 109130 699558 109132 699610
rect 109156 699558 109194 699610
rect 109194 699558 109206 699610
rect 109206 699558 109212 699610
rect 109236 699558 109258 699610
rect 109258 699558 109270 699610
rect 109270 699558 109292 699610
rect 109316 699558 109322 699610
rect 109322 699558 109334 699610
rect 109334 699558 109372 699610
rect 108836 699556 108892 699558
rect 108916 699556 108972 699558
rect 108996 699556 109052 699558
rect 109076 699556 109132 699558
rect 109156 699556 109212 699558
rect 109236 699556 109292 699558
rect 109316 699556 109372 699558
rect 144836 699610 144892 699612
rect 144916 699610 144972 699612
rect 144996 699610 145052 699612
rect 145076 699610 145132 699612
rect 145156 699610 145212 699612
rect 145236 699610 145292 699612
rect 145316 699610 145372 699612
rect 144836 699558 144874 699610
rect 144874 699558 144886 699610
rect 144886 699558 144892 699610
rect 144916 699558 144938 699610
rect 144938 699558 144950 699610
rect 144950 699558 144972 699610
rect 144996 699558 145002 699610
rect 145002 699558 145014 699610
rect 145014 699558 145052 699610
rect 145076 699558 145078 699610
rect 145078 699558 145130 699610
rect 145130 699558 145132 699610
rect 145156 699558 145194 699610
rect 145194 699558 145206 699610
rect 145206 699558 145212 699610
rect 145236 699558 145258 699610
rect 145258 699558 145270 699610
rect 145270 699558 145292 699610
rect 145316 699558 145322 699610
rect 145322 699558 145334 699610
rect 145334 699558 145372 699610
rect 144836 699556 144892 699558
rect 144916 699556 144972 699558
rect 144996 699556 145052 699558
rect 145076 699556 145132 699558
rect 145156 699556 145212 699558
rect 145236 699556 145292 699558
rect 145316 699556 145372 699558
rect 180836 699610 180892 699612
rect 180916 699610 180972 699612
rect 180996 699610 181052 699612
rect 181076 699610 181132 699612
rect 181156 699610 181212 699612
rect 181236 699610 181292 699612
rect 181316 699610 181372 699612
rect 180836 699558 180874 699610
rect 180874 699558 180886 699610
rect 180886 699558 180892 699610
rect 180916 699558 180938 699610
rect 180938 699558 180950 699610
rect 180950 699558 180972 699610
rect 180996 699558 181002 699610
rect 181002 699558 181014 699610
rect 181014 699558 181052 699610
rect 181076 699558 181078 699610
rect 181078 699558 181130 699610
rect 181130 699558 181132 699610
rect 181156 699558 181194 699610
rect 181194 699558 181206 699610
rect 181206 699558 181212 699610
rect 181236 699558 181258 699610
rect 181258 699558 181270 699610
rect 181270 699558 181292 699610
rect 181316 699558 181322 699610
rect 181322 699558 181334 699610
rect 181334 699558 181372 699610
rect 180836 699556 180892 699558
rect 180916 699556 180972 699558
rect 180996 699556 181052 699558
rect 181076 699556 181132 699558
rect 181156 699556 181212 699558
rect 181236 699556 181292 699558
rect 181316 699556 181372 699558
rect 216836 699610 216892 699612
rect 216916 699610 216972 699612
rect 216996 699610 217052 699612
rect 217076 699610 217132 699612
rect 217156 699610 217212 699612
rect 217236 699610 217292 699612
rect 217316 699610 217372 699612
rect 216836 699558 216874 699610
rect 216874 699558 216886 699610
rect 216886 699558 216892 699610
rect 216916 699558 216938 699610
rect 216938 699558 216950 699610
rect 216950 699558 216972 699610
rect 216996 699558 217002 699610
rect 217002 699558 217014 699610
rect 217014 699558 217052 699610
rect 217076 699558 217078 699610
rect 217078 699558 217130 699610
rect 217130 699558 217132 699610
rect 217156 699558 217194 699610
rect 217194 699558 217206 699610
rect 217206 699558 217212 699610
rect 217236 699558 217258 699610
rect 217258 699558 217270 699610
rect 217270 699558 217292 699610
rect 217316 699558 217322 699610
rect 217322 699558 217334 699610
rect 217334 699558 217372 699610
rect 216836 699556 216892 699558
rect 216916 699556 216972 699558
rect 216996 699556 217052 699558
rect 217076 699556 217132 699558
rect 217156 699556 217212 699558
rect 217236 699556 217292 699558
rect 217316 699556 217372 699558
rect 4802 698808 4858 698864
rect 2962 682216 3018 682272
rect 2778 667936 2834 667992
rect 3054 653520 3110 653576
rect 2962 624860 2964 624880
rect 2964 624860 3016 624880
rect 3016 624860 3018 624880
rect 2962 624824 3018 624860
rect 3146 610408 3202 610464
rect 3146 596028 3148 596048
rect 3148 596028 3200 596048
rect 3200 596028 3202 596048
rect 3146 595992 3202 596028
rect 3054 567296 3110 567352
rect 3238 538600 3294 538656
rect 3054 509904 3110 509960
rect 3422 693776 3478 693832
rect 3330 495488 3386 495544
rect 3330 481108 3332 481128
rect 3332 481108 3384 481128
rect 3384 481108 3386 481128
rect 3330 481072 3386 481108
rect 3330 452412 3332 452432
rect 3332 452412 3384 452432
rect 3384 452412 3386 452432
rect 3330 452376 3386 452412
rect 2870 423680 2926 423736
rect 3238 394984 3294 395040
rect 2778 380604 2780 380624
rect 2780 380604 2832 380624
rect 2832 380604 2834 380624
rect 2778 380568 2834 380604
rect 3238 366152 3294 366208
rect 3238 337456 3294 337512
rect 3238 308760 3294 308816
rect 3238 294344 3294 294400
rect 2778 280084 2834 280120
rect 2778 280064 2780 280084
rect 2780 280064 2832 280084
rect 2832 280064 2834 280084
rect 2962 265648 3018 265704
rect 3238 251232 3294 251288
rect 3330 236952 3386 237008
rect 3330 208156 3332 208176
rect 3332 208156 3384 208176
rect 3384 208156 3386 208176
rect 3330 208120 3386 208156
rect 2778 193840 2834 193896
rect 3330 165044 3332 165064
rect 3332 165044 3384 165064
rect 3384 165044 3386 165064
rect 3330 165008 3386 165044
rect 3330 136348 3332 136368
rect 3332 136348 3384 136368
rect 3384 136348 3386 136368
rect 3330 136312 3386 136348
rect 3330 122032 3386 122088
rect 2778 107616 2834 107672
rect 3054 78920 3110 78976
rect 3882 553016 3938 553072
rect 3790 222536 3846 222592
rect 3698 179424 3754 179480
rect 4066 437960 4122 438016
rect 3974 323040 4030 323096
rect 3882 150728 3938 150784
rect 3606 93200 3662 93256
rect 3514 64504 3570 64560
rect 3422 50088 3478 50144
rect 3422 35828 3478 35864
rect 3422 35808 3424 35828
rect 3424 35808 3476 35828
rect 3476 35808 3478 35828
rect 4986 698672 5042 698728
rect 18836 699066 18892 699068
rect 18916 699066 18972 699068
rect 18996 699066 19052 699068
rect 19076 699066 19132 699068
rect 19156 699066 19212 699068
rect 19236 699066 19292 699068
rect 19316 699066 19372 699068
rect 18836 699014 18874 699066
rect 18874 699014 18886 699066
rect 18886 699014 18892 699066
rect 18916 699014 18938 699066
rect 18938 699014 18950 699066
rect 18950 699014 18972 699066
rect 18996 699014 19002 699066
rect 19002 699014 19014 699066
rect 19014 699014 19052 699066
rect 19076 699014 19078 699066
rect 19078 699014 19130 699066
rect 19130 699014 19132 699066
rect 19156 699014 19194 699066
rect 19194 699014 19206 699066
rect 19206 699014 19212 699066
rect 19236 699014 19258 699066
rect 19258 699014 19270 699066
rect 19270 699014 19292 699066
rect 19316 699014 19322 699066
rect 19322 699014 19334 699066
rect 19334 699014 19372 699066
rect 18836 699012 18892 699014
rect 18916 699012 18972 699014
rect 18996 699012 19052 699014
rect 19076 699012 19132 699014
rect 19156 699012 19212 699014
rect 19236 699012 19292 699014
rect 19316 699012 19372 699014
rect 6182 697040 6238 697096
rect 2778 21392 2834 21448
rect 6642 694048 6698 694104
rect 7654 693640 7710 693696
rect 10322 696904 10378 696960
rect 19982 695952 20038 696008
rect 36836 698522 36892 698524
rect 36916 698522 36972 698524
rect 36996 698522 37052 698524
rect 37076 698522 37132 698524
rect 37156 698522 37212 698524
rect 37236 698522 37292 698524
rect 37316 698522 37372 698524
rect 36836 698470 36874 698522
rect 36874 698470 36886 698522
rect 36886 698470 36892 698522
rect 36916 698470 36938 698522
rect 36938 698470 36950 698522
rect 36950 698470 36972 698522
rect 36996 698470 37002 698522
rect 37002 698470 37014 698522
rect 37014 698470 37052 698522
rect 37076 698470 37078 698522
rect 37078 698470 37130 698522
rect 37130 698470 37132 698522
rect 37156 698470 37194 698522
rect 37194 698470 37206 698522
rect 37206 698470 37212 698522
rect 37236 698470 37258 698522
rect 37258 698470 37270 698522
rect 37270 698470 37292 698522
rect 37316 698470 37322 698522
rect 37322 698470 37334 698522
rect 37334 698470 37372 698522
rect 36836 698468 36892 698470
rect 36916 698468 36972 698470
rect 36996 698468 37052 698470
rect 37076 698468 37132 698470
rect 37156 698468 37212 698470
rect 37236 698468 37292 698470
rect 37316 698468 37372 698470
rect 54836 699066 54892 699068
rect 54916 699066 54972 699068
rect 54996 699066 55052 699068
rect 55076 699066 55132 699068
rect 55156 699066 55212 699068
rect 55236 699066 55292 699068
rect 55316 699066 55372 699068
rect 54836 699014 54874 699066
rect 54874 699014 54886 699066
rect 54886 699014 54892 699066
rect 54916 699014 54938 699066
rect 54938 699014 54950 699066
rect 54950 699014 54972 699066
rect 54996 699014 55002 699066
rect 55002 699014 55014 699066
rect 55014 699014 55052 699066
rect 55076 699014 55078 699066
rect 55078 699014 55130 699066
rect 55130 699014 55132 699066
rect 55156 699014 55194 699066
rect 55194 699014 55206 699066
rect 55206 699014 55212 699066
rect 55236 699014 55258 699066
rect 55258 699014 55270 699066
rect 55270 699014 55292 699066
rect 55316 699014 55322 699066
rect 55322 699014 55334 699066
rect 55334 699014 55372 699066
rect 54836 699012 54892 699014
rect 54916 699012 54972 699014
rect 54996 699012 55052 699014
rect 55076 699012 55132 699014
rect 55156 699012 55212 699014
rect 55236 699012 55292 699014
rect 55316 699012 55372 699014
rect 90836 699066 90892 699068
rect 90916 699066 90972 699068
rect 90996 699066 91052 699068
rect 91076 699066 91132 699068
rect 91156 699066 91212 699068
rect 91236 699066 91292 699068
rect 91316 699066 91372 699068
rect 90836 699014 90874 699066
rect 90874 699014 90886 699066
rect 90886 699014 90892 699066
rect 90916 699014 90938 699066
rect 90938 699014 90950 699066
rect 90950 699014 90972 699066
rect 90996 699014 91002 699066
rect 91002 699014 91014 699066
rect 91014 699014 91052 699066
rect 91076 699014 91078 699066
rect 91078 699014 91130 699066
rect 91130 699014 91132 699066
rect 91156 699014 91194 699066
rect 91194 699014 91206 699066
rect 91206 699014 91212 699066
rect 91236 699014 91258 699066
rect 91258 699014 91270 699066
rect 91270 699014 91292 699066
rect 91316 699014 91322 699066
rect 91322 699014 91334 699066
rect 91334 699014 91372 699066
rect 90836 699012 90892 699014
rect 90916 699012 90972 699014
rect 90996 699012 91052 699014
rect 91076 699012 91132 699014
rect 91156 699012 91212 699014
rect 91236 699012 91292 699014
rect 91316 699012 91372 699014
rect 72836 698522 72892 698524
rect 72916 698522 72972 698524
rect 72996 698522 73052 698524
rect 73076 698522 73132 698524
rect 73156 698522 73212 698524
rect 73236 698522 73292 698524
rect 73316 698522 73372 698524
rect 72836 698470 72874 698522
rect 72874 698470 72886 698522
rect 72886 698470 72892 698522
rect 72916 698470 72938 698522
rect 72938 698470 72950 698522
rect 72950 698470 72972 698522
rect 72996 698470 73002 698522
rect 73002 698470 73014 698522
rect 73014 698470 73052 698522
rect 73076 698470 73078 698522
rect 73078 698470 73130 698522
rect 73130 698470 73132 698522
rect 73156 698470 73194 698522
rect 73194 698470 73206 698522
rect 73206 698470 73212 698522
rect 73236 698470 73258 698522
rect 73258 698470 73270 698522
rect 73270 698470 73292 698522
rect 73316 698470 73322 698522
rect 73322 698470 73334 698522
rect 73334 698470 73372 698522
rect 72836 698468 72892 698470
rect 72916 698468 72972 698470
rect 72996 698468 73052 698470
rect 73076 698468 73132 698470
rect 73156 698468 73212 698470
rect 73236 698468 73292 698470
rect 73316 698468 73372 698470
rect 89718 696088 89774 696144
rect 126836 699066 126892 699068
rect 126916 699066 126972 699068
rect 126996 699066 127052 699068
rect 127076 699066 127132 699068
rect 127156 699066 127212 699068
rect 127236 699066 127292 699068
rect 127316 699066 127372 699068
rect 126836 699014 126874 699066
rect 126874 699014 126886 699066
rect 126886 699014 126892 699066
rect 126916 699014 126938 699066
rect 126938 699014 126950 699066
rect 126950 699014 126972 699066
rect 126996 699014 127002 699066
rect 127002 699014 127014 699066
rect 127014 699014 127052 699066
rect 127076 699014 127078 699066
rect 127078 699014 127130 699066
rect 127130 699014 127132 699066
rect 127156 699014 127194 699066
rect 127194 699014 127206 699066
rect 127206 699014 127212 699066
rect 127236 699014 127258 699066
rect 127258 699014 127270 699066
rect 127270 699014 127292 699066
rect 127316 699014 127322 699066
rect 127322 699014 127334 699066
rect 127334 699014 127372 699066
rect 126836 699012 126892 699014
rect 126916 699012 126972 699014
rect 126996 699012 127052 699014
rect 127076 699012 127132 699014
rect 127156 699012 127212 699014
rect 127236 699012 127292 699014
rect 127316 699012 127372 699014
rect 108836 698522 108892 698524
rect 108916 698522 108972 698524
rect 108996 698522 109052 698524
rect 109076 698522 109132 698524
rect 109156 698522 109212 698524
rect 109236 698522 109292 698524
rect 109316 698522 109372 698524
rect 108836 698470 108874 698522
rect 108874 698470 108886 698522
rect 108886 698470 108892 698522
rect 108916 698470 108938 698522
rect 108938 698470 108950 698522
rect 108950 698470 108972 698522
rect 108996 698470 109002 698522
rect 109002 698470 109014 698522
rect 109014 698470 109052 698522
rect 109076 698470 109078 698522
rect 109078 698470 109130 698522
rect 109130 698470 109132 698522
rect 109156 698470 109194 698522
rect 109194 698470 109206 698522
rect 109206 698470 109212 698522
rect 109236 698470 109258 698522
rect 109258 698470 109270 698522
rect 109270 698470 109292 698522
rect 109316 698470 109322 698522
rect 109322 698470 109334 698522
rect 109334 698470 109372 698522
rect 108836 698468 108892 698470
rect 108916 698468 108972 698470
rect 108996 698468 109052 698470
rect 109076 698468 109132 698470
rect 109156 698468 109212 698470
rect 109236 698468 109292 698470
rect 109316 698468 109372 698470
rect 144836 698522 144892 698524
rect 144916 698522 144972 698524
rect 144996 698522 145052 698524
rect 145076 698522 145132 698524
rect 145156 698522 145212 698524
rect 145236 698522 145292 698524
rect 145316 698522 145372 698524
rect 144836 698470 144874 698522
rect 144874 698470 144886 698522
rect 144886 698470 144892 698522
rect 144916 698470 144938 698522
rect 144938 698470 144950 698522
rect 144950 698470 144972 698522
rect 144996 698470 145002 698522
rect 145002 698470 145014 698522
rect 145014 698470 145052 698522
rect 145076 698470 145078 698522
rect 145078 698470 145130 698522
rect 145130 698470 145132 698522
rect 145156 698470 145194 698522
rect 145194 698470 145206 698522
rect 145206 698470 145212 698522
rect 145236 698470 145258 698522
rect 145258 698470 145270 698522
rect 145270 698470 145292 698522
rect 145316 698470 145322 698522
rect 145322 698470 145334 698522
rect 145334 698470 145372 698522
rect 144836 698468 144892 698470
rect 144916 698468 144972 698470
rect 144996 698468 145052 698470
rect 145076 698468 145132 698470
rect 145156 698468 145212 698470
rect 145236 698468 145292 698470
rect 145316 698468 145372 698470
rect 186134 699236 186190 699272
rect 186134 699216 186136 699236
rect 186136 699216 186188 699236
rect 186188 699216 186190 699236
rect 162836 699066 162892 699068
rect 162916 699066 162972 699068
rect 162996 699066 163052 699068
rect 163076 699066 163132 699068
rect 163156 699066 163212 699068
rect 163236 699066 163292 699068
rect 163316 699066 163372 699068
rect 162836 699014 162874 699066
rect 162874 699014 162886 699066
rect 162886 699014 162892 699066
rect 162916 699014 162938 699066
rect 162938 699014 162950 699066
rect 162950 699014 162972 699066
rect 162996 699014 163002 699066
rect 163002 699014 163014 699066
rect 163014 699014 163052 699066
rect 163076 699014 163078 699066
rect 163078 699014 163130 699066
rect 163130 699014 163132 699066
rect 163156 699014 163194 699066
rect 163194 699014 163206 699066
rect 163206 699014 163212 699066
rect 163236 699014 163258 699066
rect 163258 699014 163270 699066
rect 163270 699014 163292 699066
rect 163316 699014 163322 699066
rect 163322 699014 163334 699066
rect 163334 699014 163372 699066
rect 162836 699012 162892 699014
rect 162916 699012 162972 699014
rect 162996 699012 163052 699014
rect 163076 699012 163132 699014
rect 163156 699012 163212 699014
rect 163236 699012 163292 699014
rect 163316 699012 163372 699014
rect 198836 699066 198892 699068
rect 198916 699066 198972 699068
rect 198996 699066 199052 699068
rect 199076 699066 199132 699068
rect 199156 699066 199212 699068
rect 199236 699066 199292 699068
rect 199316 699066 199372 699068
rect 198836 699014 198874 699066
rect 198874 699014 198886 699066
rect 198886 699014 198892 699066
rect 198916 699014 198938 699066
rect 198938 699014 198950 699066
rect 198950 699014 198972 699066
rect 198996 699014 199002 699066
rect 199002 699014 199014 699066
rect 199014 699014 199052 699066
rect 199076 699014 199078 699066
rect 199078 699014 199130 699066
rect 199130 699014 199132 699066
rect 199156 699014 199194 699066
rect 199194 699014 199206 699066
rect 199206 699014 199212 699066
rect 199236 699014 199258 699066
rect 199258 699014 199270 699066
rect 199270 699014 199292 699066
rect 199316 699014 199322 699066
rect 199322 699014 199334 699066
rect 199334 699014 199372 699066
rect 198836 699012 198892 699014
rect 198916 699012 198972 699014
rect 198996 699012 199052 699014
rect 199076 699012 199132 699014
rect 199156 699012 199212 699014
rect 199236 699012 199292 699014
rect 199316 699012 199372 699014
rect 180836 698522 180892 698524
rect 180916 698522 180972 698524
rect 180996 698522 181052 698524
rect 181076 698522 181132 698524
rect 181156 698522 181212 698524
rect 181236 698522 181292 698524
rect 181316 698522 181372 698524
rect 180836 698470 180874 698522
rect 180874 698470 180886 698522
rect 180886 698470 180892 698522
rect 180916 698470 180938 698522
rect 180938 698470 180950 698522
rect 180950 698470 180972 698522
rect 180996 698470 181002 698522
rect 181002 698470 181014 698522
rect 181014 698470 181052 698522
rect 181076 698470 181078 698522
rect 181078 698470 181130 698522
rect 181130 698470 181132 698522
rect 181156 698470 181194 698522
rect 181194 698470 181206 698522
rect 181206 698470 181212 698522
rect 181236 698470 181258 698522
rect 181258 698470 181270 698522
rect 181270 698470 181292 698522
rect 181316 698470 181322 698522
rect 181322 698470 181334 698522
rect 181334 698470 181372 698522
rect 180836 698468 180892 698470
rect 180916 698468 180972 698470
rect 180996 698468 181052 698470
rect 181076 698468 181132 698470
rect 181156 698468 181212 698470
rect 181236 698468 181292 698470
rect 181316 698468 181372 698470
rect 216836 698522 216892 698524
rect 216916 698522 216972 698524
rect 216996 698522 217052 698524
rect 217076 698522 217132 698524
rect 217156 698522 217212 698524
rect 217236 698522 217292 698524
rect 217316 698522 217372 698524
rect 216836 698470 216874 698522
rect 216874 698470 216886 698522
rect 216886 698470 216892 698522
rect 216916 698470 216938 698522
rect 216938 698470 216950 698522
rect 216950 698470 216972 698522
rect 216996 698470 217002 698522
rect 217002 698470 217014 698522
rect 217014 698470 217052 698522
rect 217076 698470 217078 698522
rect 217078 698470 217130 698522
rect 217130 698470 217132 698522
rect 217156 698470 217194 698522
rect 217194 698470 217206 698522
rect 217206 698470 217212 698522
rect 217236 698470 217258 698522
rect 217258 698470 217270 698522
rect 217270 698470 217292 698522
rect 217316 698470 217322 698522
rect 217322 698470 217334 698522
rect 217334 698470 217372 698522
rect 216836 698468 216892 698470
rect 216916 698468 216972 698470
rect 216996 698468 217052 698470
rect 217076 698468 217132 698470
rect 217156 698468 217212 698470
rect 217236 698468 217292 698470
rect 217316 698468 217372 698470
rect 218058 698420 218114 698456
rect 218058 698400 218060 698420
rect 218060 698400 218112 698420
rect 218112 698400 218114 698420
rect 218426 698420 218482 698456
rect 218426 698400 218428 698420
rect 218428 698400 218480 698420
rect 218480 698400 218482 698420
rect 218058 698284 218114 698320
rect 218058 698264 218060 698284
rect 218060 698264 218112 698284
rect 218112 698264 218114 698284
rect 218426 698284 218482 698320
rect 218426 698264 218428 698284
rect 218428 698264 218480 698284
rect 218480 698264 218482 698284
rect 208950 698148 209006 698184
rect 215114 698164 215116 698184
rect 215116 698164 215168 698184
rect 215168 698164 215170 698184
rect 208950 698128 208952 698148
rect 208952 698128 209004 698148
rect 209004 698128 209006 698148
rect 215114 698128 215170 698164
rect 193310 697992 193366 698048
rect 202786 697992 202842 698048
rect 205546 695952 205602 696008
rect 213734 695952 213790 696008
rect 234836 701242 234892 701244
rect 234916 701242 234972 701244
rect 234996 701242 235052 701244
rect 235076 701242 235132 701244
rect 235156 701242 235212 701244
rect 235236 701242 235292 701244
rect 235316 701242 235372 701244
rect 234836 701190 234874 701242
rect 234874 701190 234886 701242
rect 234886 701190 234892 701242
rect 234916 701190 234938 701242
rect 234938 701190 234950 701242
rect 234950 701190 234972 701242
rect 234996 701190 235002 701242
rect 235002 701190 235014 701242
rect 235014 701190 235052 701242
rect 235076 701190 235078 701242
rect 235078 701190 235130 701242
rect 235130 701190 235132 701242
rect 235156 701190 235194 701242
rect 235194 701190 235206 701242
rect 235206 701190 235212 701242
rect 235236 701190 235258 701242
rect 235258 701190 235270 701242
rect 235270 701190 235292 701242
rect 235316 701190 235322 701242
rect 235322 701190 235334 701242
rect 235334 701190 235372 701242
rect 234836 701188 234892 701190
rect 234916 701188 234972 701190
rect 234996 701188 235052 701190
rect 235076 701188 235132 701190
rect 235156 701188 235212 701190
rect 235236 701188 235292 701190
rect 235316 701188 235372 701190
rect 227994 700848 228050 700904
rect 226338 698264 226394 698320
rect 224958 696380 225014 696416
rect 224958 696360 224960 696380
rect 224960 696360 225012 696380
rect 225012 696360 225014 696380
rect 234836 700154 234892 700156
rect 234916 700154 234972 700156
rect 234996 700154 235052 700156
rect 235076 700154 235132 700156
rect 235156 700154 235212 700156
rect 235236 700154 235292 700156
rect 235316 700154 235372 700156
rect 234836 700102 234874 700154
rect 234874 700102 234886 700154
rect 234886 700102 234892 700154
rect 234916 700102 234938 700154
rect 234938 700102 234950 700154
rect 234950 700102 234972 700154
rect 234996 700102 235002 700154
rect 235002 700102 235014 700154
rect 235014 700102 235052 700154
rect 235076 700102 235078 700154
rect 235078 700102 235130 700154
rect 235130 700102 235132 700154
rect 235156 700102 235194 700154
rect 235194 700102 235206 700154
rect 235206 700102 235212 700154
rect 235236 700102 235258 700154
rect 235258 700102 235270 700154
rect 235270 700102 235292 700154
rect 235316 700102 235322 700154
rect 235322 700102 235334 700154
rect 235334 700102 235372 700154
rect 234836 700100 234892 700102
rect 234916 700100 234972 700102
rect 234996 700100 235052 700102
rect 235076 700100 235132 700102
rect 235156 700100 235212 700102
rect 235236 700100 235292 700102
rect 235316 700100 235372 700102
rect 234836 699066 234892 699068
rect 234916 699066 234972 699068
rect 234996 699066 235052 699068
rect 235076 699066 235132 699068
rect 235156 699066 235212 699068
rect 235236 699066 235292 699068
rect 235316 699066 235372 699068
rect 234836 699014 234874 699066
rect 234874 699014 234886 699066
rect 234886 699014 234892 699066
rect 234916 699014 234938 699066
rect 234938 699014 234950 699066
rect 234950 699014 234972 699066
rect 234996 699014 235002 699066
rect 235002 699014 235014 699066
rect 235014 699014 235052 699066
rect 235076 699014 235078 699066
rect 235078 699014 235130 699066
rect 235130 699014 235132 699066
rect 235156 699014 235194 699066
rect 235194 699014 235206 699066
rect 235206 699014 235212 699066
rect 235236 699014 235258 699066
rect 235258 699014 235270 699066
rect 235270 699014 235292 699066
rect 235316 699014 235322 699066
rect 235322 699014 235334 699066
rect 235334 699014 235372 699066
rect 234836 699012 234892 699014
rect 234916 699012 234972 699014
rect 234996 699012 235052 699014
rect 235076 699012 235132 699014
rect 235156 699012 235212 699014
rect 235236 699012 235292 699014
rect 235316 699012 235372 699014
rect 235906 698264 235962 698320
rect 237378 698164 237380 698184
rect 237380 698164 237432 698184
rect 237432 698164 237434 698184
rect 237378 698128 237434 698164
rect 232962 696768 233018 696824
rect 229006 695952 229062 696008
rect 230386 695952 230442 696008
rect 234526 696788 234582 696824
rect 234526 696768 234528 696788
rect 234528 696768 234580 696788
rect 234580 696768 234582 696788
rect 234526 696380 234582 696416
rect 234526 696360 234528 696380
rect 234528 696360 234580 696380
rect 234580 696360 234582 696380
rect 237562 698164 237564 698184
rect 237564 698164 237616 698184
rect 237616 698164 237618 698184
rect 237562 698128 237618 698164
rect 244094 699216 244150 699272
rect 244094 698964 244150 699000
rect 244278 699216 244334 699272
rect 244094 698944 244096 698964
rect 244096 698944 244148 698964
rect 244148 698944 244150 698964
rect 244370 698964 244426 699000
rect 244370 698944 244372 698964
rect 244372 698944 244424 698964
rect 244424 698944 244426 698964
rect 244278 696788 244334 696824
rect 244278 696768 244280 696788
rect 244280 696768 244332 696788
rect 244332 696768 244334 696788
rect 244278 696380 244334 696416
rect 244278 696360 244280 696380
rect 244280 696360 244332 696380
rect 244332 696360 244334 696380
rect 248326 698264 248382 698320
rect 248418 696768 248474 696824
rect 251086 695952 251142 696008
rect 252836 701786 252892 701788
rect 252916 701786 252972 701788
rect 252996 701786 253052 701788
rect 253076 701786 253132 701788
rect 253156 701786 253212 701788
rect 253236 701786 253292 701788
rect 253316 701786 253372 701788
rect 252836 701734 252874 701786
rect 252874 701734 252886 701786
rect 252886 701734 252892 701786
rect 252916 701734 252938 701786
rect 252938 701734 252950 701786
rect 252950 701734 252972 701786
rect 252996 701734 253002 701786
rect 253002 701734 253014 701786
rect 253014 701734 253052 701786
rect 253076 701734 253078 701786
rect 253078 701734 253130 701786
rect 253130 701734 253132 701786
rect 253156 701734 253194 701786
rect 253194 701734 253206 701786
rect 253206 701734 253212 701786
rect 253236 701734 253258 701786
rect 253258 701734 253270 701786
rect 253270 701734 253292 701786
rect 253316 701734 253322 701786
rect 253322 701734 253334 701786
rect 253334 701734 253372 701786
rect 252836 701732 252892 701734
rect 252916 701732 252972 701734
rect 252996 701732 253052 701734
rect 253076 701732 253132 701734
rect 253156 701732 253212 701734
rect 253236 701732 253292 701734
rect 253316 701732 253372 701734
rect 252836 700698 252892 700700
rect 252916 700698 252972 700700
rect 252996 700698 253052 700700
rect 253076 700698 253132 700700
rect 253156 700698 253212 700700
rect 253236 700698 253292 700700
rect 253316 700698 253372 700700
rect 252836 700646 252874 700698
rect 252874 700646 252886 700698
rect 252886 700646 252892 700698
rect 252916 700646 252938 700698
rect 252938 700646 252950 700698
rect 252950 700646 252972 700698
rect 252996 700646 253002 700698
rect 253002 700646 253014 700698
rect 253014 700646 253052 700698
rect 253076 700646 253078 700698
rect 253078 700646 253130 700698
rect 253130 700646 253132 700698
rect 253156 700646 253194 700698
rect 253194 700646 253206 700698
rect 253206 700646 253212 700698
rect 253236 700646 253258 700698
rect 253258 700646 253270 700698
rect 253270 700646 253292 700698
rect 253316 700646 253322 700698
rect 253322 700646 253334 700698
rect 253334 700646 253372 700698
rect 252836 700644 252892 700646
rect 252916 700644 252972 700646
rect 252996 700644 253052 700646
rect 253076 700644 253132 700646
rect 253156 700644 253212 700646
rect 253236 700644 253292 700646
rect 253316 700644 253372 700646
rect 252836 699610 252892 699612
rect 252916 699610 252972 699612
rect 252996 699610 253052 699612
rect 253076 699610 253132 699612
rect 253156 699610 253212 699612
rect 253236 699610 253292 699612
rect 253316 699610 253372 699612
rect 252836 699558 252874 699610
rect 252874 699558 252886 699610
rect 252886 699558 252892 699610
rect 252916 699558 252938 699610
rect 252938 699558 252950 699610
rect 252950 699558 252972 699610
rect 252996 699558 253002 699610
rect 253002 699558 253014 699610
rect 253014 699558 253052 699610
rect 253076 699558 253078 699610
rect 253078 699558 253130 699610
rect 253130 699558 253132 699610
rect 253156 699558 253194 699610
rect 253194 699558 253206 699610
rect 253206 699558 253212 699610
rect 253236 699558 253258 699610
rect 253258 699558 253270 699610
rect 253270 699558 253292 699610
rect 253316 699558 253322 699610
rect 253322 699558 253334 699610
rect 253334 699558 253372 699610
rect 252836 699556 252892 699558
rect 252916 699556 252972 699558
rect 252996 699556 253052 699558
rect 253076 699556 253132 699558
rect 253156 699556 253212 699558
rect 253236 699556 253292 699558
rect 253316 699556 253372 699558
rect 253754 698964 253810 699000
rect 253754 698944 253756 698964
rect 253756 698944 253808 698964
rect 253808 698944 253810 698964
rect 252836 698522 252892 698524
rect 252916 698522 252972 698524
rect 252996 698522 253052 698524
rect 253076 698522 253132 698524
rect 253156 698522 253212 698524
rect 253236 698522 253292 698524
rect 253316 698522 253372 698524
rect 252836 698470 252874 698522
rect 252874 698470 252886 698522
rect 252886 698470 252892 698522
rect 252916 698470 252938 698522
rect 252938 698470 252950 698522
rect 252950 698470 252972 698522
rect 252996 698470 253002 698522
rect 253002 698470 253014 698522
rect 253014 698470 253052 698522
rect 253076 698470 253078 698522
rect 253078 698470 253130 698522
rect 253130 698470 253132 698522
rect 253156 698470 253194 698522
rect 253194 698470 253206 698522
rect 253206 698470 253212 698522
rect 253236 698470 253258 698522
rect 253258 698470 253270 698522
rect 253270 698470 253292 698522
rect 253316 698470 253322 698522
rect 253322 698470 253334 698522
rect 253334 698470 253372 698522
rect 252836 698468 252892 698470
rect 252916 698468 252972 698470
rect 252996 698468 253052 698470
rect 253076 698468 253132 698470
rect 253156 698468 253212 698470
rect 253236 698468 253292 698470
rect 253316 698468 253372 698470
rect 253846 698264 253902 698320
rect 253846 698164 253848 698184
rect 253848 698164 253900 698184
rect 253900 698164 253902 698184
rect 253846 698128 253902 698164
rect 254030 698164 254032 698184
rect 254032 698164 254084 698184
rect 254084 698164 254086 698184
rect 254030 698128 254086 698164
rect 253846 696380 253902 696416
rect 253846 696360 253848 696380
rect 253848 696360 253900 696380
rect 253900 696360 253902 696380
rect 259458 699488 259514 699544
rect 263598 696380 263654 696416
rect 263598 696360 263600 696380
rect 263600 696360 263652 696380
rect 263652 696360 263654 696380
rect 265622 695952 265678 696008
rect 270836 701242 270892 701244
rect 270916 701242 270972 701244
rect 270996 701242 271052 701244
rect 271076 701242 271132 701244
rect 271156 701242 271212 701244
rect 271236 701242 271292 701244
rect 271316 701242 271372 701244
rect 270836 701190 270874 701242
rect 270874 701190 270886 701242
rect 270886 701190 270892 701242
rect 270916 701190 270938 701242
rect 270938 701190 270950 701242
rect 270950 701190 270972 701242
rect 270996 701190 271002 701242
rect 271002 701190 271014 701242
rect 271014 701190 271052 701242
rect 271076 701190 271078 701242
rect 271078 701190 271130 701242
rect 271130 701190 271132 701242
rect 271156 701190 271194 701242
rect 271194 701190 271206 701242
rect 271206 701190 271212 701242
rect 271236 701190 271258 701242
rect 271258 701190 271270 701242
rect 271270 701190 271292 701242
rect 271316 701190 271322 701242
rect 271322 701190 271334 701242
rect 271334 701190 271372 701242
rect 270836 701188 270892 701190
rect 270916 701188 270972 701190
rect 270996 701188 271052 701190
rect 271076 701188 271132 701190
rect 271156 701188 271212 701190
rect 271236 701188 271292 701190
rect 271316 701188 271372 701190
rect 270836 700154 270892 700156
rect 270916 700154 270972 700156
rect 270996 700154 271052 700156
rect 271076 700154 271132 700156
rect 271156 700154 271212 700156
rect 271236 700154 271292 700156
rect 271316 700154 271372 700156
rect 270836 700102 270874 700154
rect 270874 700102 270886 700154
rect 270886 700102 270892 700154
rect 270916 700102 270938 700154
rect 270938 700102 270950 700154
rect 270950 700102 270972 700154
rect 270996 700102 271002 700154
rect 271002 700102 271014 700154
rect 271014 700102 271052 700154
rect 271076 700102 271078 700154
rect 271078 700102 271130 700154
rect 271130 700102 271132 700154
rect 271156 700102 271194 700154
rect 271194 700102 271206 700154
rect 271206 700102 271212 700154
rect 271236 700102 271258 700154
rect 271258 700102 271270 700154
rect 271270 700102 271292 700154
rect 271316 700102 271322 700154
rect 271322 700102 271334 700154
rect 271334 700102 271372 700154
rect 270836 700100 270892 700102
rect 270916 700100 270972 700102
rect 270996 700100 271052 700102
rect 271076 700100 271132 700102
rect 271156 700100 271212 700102
rect 271236 700100 271292 700102
rect 271316 700100 271372 700102
rect 283102 700032 283158 700088
rect 267646 699236 267702 699272
rect 267646 699216 267648 699236
rect 267648 699216 267700 699236
rect 267700 699216 267702 699236
rect 273902 699780 273958 699816
rect 273902 699760 273904 699780
rect 273904 699760 273956 699780
rect 273956 699760 273958 699780
rect 280066 699624 280122 699680
rect 283010 699660 283012 699680
rect 283012 699660 283064 699680
rect 283064 699660 283066 699680
rect 273258 699352 273314 699408
rect 273350 699216 273406 699272
rect 277398 699216 277454 699272
rect 270836 699066 270892 699068
rect 270916 699066 270972 699068
rect 270996 699066 271052 699068
rect 271076 699066 271132 699068
rect 271156 699066 271212 699068
rect 271236 699066 271292 699068
rect 271316 699066 271372 699068
rect 270836 699014 270874 699066
rect 270874 699014 270886 699066
rect 270886 699014 270892 699066
rect 270916 699014 270938 699066
rect 270938 699014 270950 699066
rect 270950 699014 270972 699066
rect 270996 699014 271002 699066
rect 271002 699014 271014 699066
rect 271014 699014 271052 699066
rect 271076 699014 271078 699066
rect 271078 699014 271130 699066
rect 271130 699014 271132 699066
rect 271156 699014 271194 699066
rect 271194 699014 271206 699066
rect 271206 699014 271212 699066
rect 271236 699014 271258 699066
rect 271258 699014 271270 699066
rect 271270 699014 271292 699066
rect 271316 699014 271322 699066
rect 271322 699014 271334 699066
rect 271334 699014 271372 699066
rect 270836 699012 270892 699014
rect 270916 699012 270972 699014
rect 270996 699012 271052 699014
rect 271076 699012 271132 699014
rect 271156 699012 271212 699014
rect 271236 699012 271292 699014
rect 271316 699012 271372 699014
rect 275742 698128 275798 698184
rect 277398 698128 277454 698184
rect 273166 696380 273222 696416
rect 273166 696360 273168 696380
rect 273168 696360 273220 696380
rect 273220 696360 273222 696380
rect 283010 699624 283066 699660
rect 283010 699372 283066 699408
rect 283010 699352 283012 699372
rect 283012 699352 283064 699372
rect 283064 699352 283066 699372
rect 282918 699080 282974 699136
rect 283746 699780 283802 699816
rect 288836 701786 288892 701788
rect 288916 701786 288972 701788
rect 288996 701786 289052 701788
rect 289076 701786 289132 701788
rect 289156 701786 289212 701788
rect 289236 701786 289292 701788
rect 289316 701786 289372 701788
rect 288836 701734 288874 701786
rect 288874 701734 288886 701786
rect 288886 701734 288892 701786
rect 288916 701734 288938 701786
rect 288938 701734 288950 701786
rect 288950 701734 288972 701786
rect 288996 701734 289002 701786
rect 289002 701734 289014 701786
rect 289014 701734 289052 701786
rect 289076 701734 289078 701786
rect 289078 701734 289130 701786
rect 289130 701734 289132 701786
rect 289156 701734 289194 701786
rect 289194 701734 289206 701786
rect 289206 701734 289212 701786
rect 289236 701734 289258 701786
rect 289258 701734 289270 701786
rect 289270 701734 289292 701786
rect 289316 701734 289322 701786
rect 289322 701734 289334 701786
rect 289334 701734 289372 701786
rect 288836 701732 288892 701734
rect 288916 701732 288972 701734
rect 288996 701732 289052 701734
rect 289076 701732 289132 701734
rect 289156 701732 289212 701734
rect 289236 701732 289292 701734
rect 289316 701732 289372 701734
rect 288836 700698 288892 700700
rect 288916 700698 288972 700700
rect 288996 700698 289052 700700
rect 289076 700698 289132 700700
rect 289156 700698 289212 700700
rect 289236 700698 289292 700700
rect 289316 700698 289372 700700
rect 288836 700646 288874 700698
rect 288874 700646 288886 700698
rect 288886 700646 288892 700698
rect 288916 700646 288938 700698
rect 288938 700646 288950 700698
rect 288950 700646 288972 700698
rect 288996 700646 289002 700698
rect 289002 700646 289014 700698
rect 289014 700646 289052 700698
rect 289076 700646 289078 700698
rect 289078 700646 289130 700698
rect 289130 700646 289132 700698
rect 289156 700646 289194 700698
rect 289194 700646 289206 700698
rect 289206 700646 289212 700698
rect 289236 700646 289258 700698
rect 289258 700646 289270 700698
rect 289270 700646 289292 700698
rect 289316 700646 289322 700698
rect 289322 700646 289334 700698
rect 289334 700646 289372 700698
rect 288836 700644 288892 700646
rect 288916 700644 288972 700646
rect 288996 700644 289052 700646
rect 289076 700644 289132 700646
rect 289156 700644 289212 700646
rect 289236 700644 289292 700646
rect 289316 700644 289372 700646
rect 296534 700168 296590 700224
rect 298650 700168 298706 700224
rect 296626 700032 296682 700088
rect 298006 699916 298062 699952
rect 298006 699896 298008 699916
rect 298008 699896 298060 699916
rect 298060 699896 298062 699916
rect 283746 699760 283748 699780
rect 283748 699760 283800 699780
rect 283800 699760 283802 699780
rect 288714 699760 288770 699816
rect 296718 699760 296774 699816
rect 282918 696380 282974 696416
rect 282918 696360 282920 696380
rect 282920 696360 282972 696380
rect 282972 696360 282974 696380
rect 288836 699610 288892 699612
rect 288916 699610 288972 699612
rect 288996 699610 289052 699612
rect 289076 699610 289132 699612
rect 289156 699610 289212 699612
rect 289236 699610 289292 699612
rect 289316 699610 289372 699612
rect 288836 699558 288874 699610
rect 288874 699558 288886 699610
rect 288886 699558 288892 699610
rect 288916 699558 288938 699610
rect 288938 699558 288950 699610
rect 288950 699558 288972 699610
rect 288996 699558 289002 699610
rect 289002 699558 289014 699610
rect 289014 699558 289052 699610
rect 289076 699558 289078 699610
rect 289078 699558 289130 699610
rect 289130 699558 289132 699610
rect 289156 699558 289194 699610
rect 289194 699558 289206 699610
rect 289206 699558 289212 699610
rect 289236 699558 289258 699610
rect 289258 699558 289270 699610
rect 289270 699558 289292 699610
rect 289316 699558 289322 699610
rect 289322 699558 289334 699610
rect 289334 699558 289372 699610
rect 288836 699556 288892 699558
rect 288916 699556 288972 699558
rect 288996 699556 289052 699558
rect 289076 699556 289132 699558
rect 289156 699556 289212 699558
rect 289236 699556 289292 699558
rect 289316 699556 289372 699558
rect 289726 699488 289782 699544
rect 288836 698522 288892 698524
rect 288916 698522 288972 698524
rect 288996 698522 289052 698524
rect 289076 698522 289132 698524
rect 289156 698522 289212 698524
rect 289236 698522 289292 698524
rect 289316 698522 289372 698524
rect 288836 698470 288874 698522
rect 288874 698470 288886 698522
rect 288886 698470 288892 698522
rect 288916 698470 288938 698522
rect 288938 698470 288950 698522
rect 288950 698470 288972 698522
rect 288996 698470 289002 698522
rect 289002 698470 289014 698522
rect 289014 698470 289052 698522
rect 289076 698470 289078 698522
rect 289078 698470 289130 698522
rect 289130 698470 289132 698522
rect 289156 698470 289194 698522
rect 289194 698470 289206 698522
rect 289206 698470 289212 698522
rect 289236 698470 289258 698522
rect 289258 698470 289270 698522
rect 289270 698470 289292 698522
rect 289316 698470 289322 698522
rect 289322 698470 289334 698522
rect 289334 698470 289372 698522
rect 288836 698468 288892 698470
rect 288916 698468 288972 698470
rect 288996 698468 289052 698470
rect 289076 698468 289132 698470
rect 289156 698468 289212 698470
rect 289236 698468 289292 698470
rect 289316 698468 289372 698470
rect 292394 699352 292450 699408
rect 296902 699488 296958 699544
rect 294050 699352 294106 699408
rect 292486 699216 292542 699272
rect 119986 695680 120042 695736
rect 120170 695544 120226 695600
rect 176198 695544 176254 695600
rect 205546 695544 205602 695600
rect 213734 695544 213790 695600
rect 215206 695544 215262 695600
rect 234618 695680 234674 695736
rect 230386 695544 230442 695600
rect 234526 695544 234582 695600
rect 292486 696380 292542 696416
rect 292486 696360 292488 696380
rect 292488 696360 292540 696380
rect 292540 696360 292542 696380
rect 296534 699216 296590 699272
rect 296626 699080 296682 699136
rect 324836 701786 324892 701788
rect 324916 701786 324972 701788
rect 324996 701786 325052 701788
rect 325076 701786 325132 701788
rect 325156 701786 325212 701788
rect 325236 701786 325292 701788
rect 325316 701786 325372 701788
rect 324836 701734 324874 701786
rect 324874 701734 324886 701786
rect 324886 701734 324892 701786
rect 324916 701734 324938 701786
rect 324938 701734 324950 701786
rect 324950 701734 324972 701786
rect 324996 701734 325002 701786
rect 325002 701734 325014 701786
rect 325014 701734 325052 701786
rect 325076 701734 325078 701786
rect 325078 701734 325130 701786
rect 325130 701734 325132 701786
rect 325156 701734 325194 701786
rect 325194 701734 325206 701786
rect 325206 701734 325212 701786
rect 325236 701734 325258 701786
rect 325258 701734 325270 701786
rect 325270 701734 325292 701786
rect 325316 701734 325322 701786
rect 325322 701734 325334 701786
rect 325334 701734 325372 701786
rect 324836 701732 324892 701734
rect 324916 701732 324972 701734
rect 324996 701732 325052 701734
rect 325076 701732 325132 701734
rect 325156 701732 325212 701734
rect 325236 701732 325292 701734
rect 325316 701732 325372 701734
rect 306836 701242 306892 701244
rect 306916 701242 306972 701244
rect 306996 701242 307052 701244
rect 307076 701242 307132 701244
rect 307156 701242 307212 701244
rect 307236 701242 307292 701244
rect 307316 701242 307372 701244
rect 306836 701190 306874 701242
rect 306874 701190 306886 701242
rect 306886 701190 306892 701242
rect 306916 701190 306938 701242
rect 306938 701190 306950 701242
rect 306950 701190 306972 701242
rect 306996 701190 307002 701242
rect 307002 701190 307014 701242
rect 307014 701190 307052 701242
rect 307076 701190 307078 701242
rect 307078 701190 307130 701242
rect 307130 701190 307132 701242
rect 307156 701190 307194 701242
rect 307194 701190 307206 701242
rect 307206 701190 307212 701242
rect 307236 701190 307258 701242
rect 307258 701190 307270 701242
rect 307270 701190 307292 701242
rect 307316 701190 307322 701242
rect 307322 701190 307334 701242
rect 307334 701190 307372 701242
rect 306836 701188 306892 701190
rect 306916 701188 306972 701190
rect 306996 701188 307052 701190
rect 307076 701188 307132 701190
rect 307156 701188 307212 701190
rect 307236 701188 307292 701190
rect 307316 701188 307372 701190
rect 306836 700154 306892 700156
rect 306916 700154 306972 700156
rect 306996 700154 307052 700156
rect 307076 700154 307132 700156
rect 307156 700154 307212 700156
rect 307236 700154 307292 700156
rect 307316 700154 307372 700156
rect 306836 700102 306874 700154
rect 306874 700102 306886 700154
rect 306886 700102 306892 700154
rect 306916 700102 306938 700154
rect 306938 700102 306950 700154
rect 306950 700102 306972 700154
rect 306996 700102 307002 700154
rect 307002 700102 307014 700154
rect 307014 700102 307052 700154
rect 307076 700102 307078 700154
rect 307078 700102 307130 700154
rect 307130 700102 307132 700154
rect 307156 700102 307194 700154
rect 307194 700102 307206 700154
rect 307206 700102 307212 700154
rect 307236 700102 307258 700154
rect 307258 700102 307270 700154
rect 307270 700102 307292 700154
rect 307316 700102 307322 700154
rect 307322 700102 307334 700154
rect 307334 700102 307372 700154
rect 306836 700100 306892 700102
rect 306916 700100 306972 700102
rect 306996 700100 307052 700102
rect 307076 700100 307132 700102
rect 307156 700100 307212 700102
rect 307236 700100 307292 700102
rect 307316 700100 307372 700102
rect 300122 699896 300178 699952
rect 302330 699896 302386 699952
rect 303618 699760 303674 699816
rect 302330 699236 302386 699272
rect 302330 699216 302332 699236
rect 302332 699216 302384 699236
rect 302384 699216 302386 699236
rect 299478 696632 299534 696688
rect 306836 699066 306892 699068
rect 306916 699066 306972 699068
rect 306996 699066 307052 699068
rect 307076 699066 307132 699068
rect 307156 699066 307212 699068
rect 307236 699066 307292 699068
rect 307316 699066 307372 699068
rect 306836 699014 306874 699066
rect 306874 699014 306886 699066
rect 306886 699014 306892 699066
rect 306916 699014 306938 699066
rect 306938 699014 306950 699066
rect 306950 699014 306972 699066
rect 306996 699014 307002 699066
rect 307002 699014 307014 699066
rect 307014 699014 307052 699066
rect 307076 699014 307078 699066
rect 307078 699014 307130 699066
rect 307130 699014 307132 699066
rect 307156 699014 307194 699066
rect 307194 699014 307206 699066
rect 307206 699014 307212 699066
rect 307236 699014 307258 699066
rect 307258 699014 307270 699066
rect 307270 699014 307292 699066
rect 307316 699014 307322 699066
rect 307322 699014 307334 699066
rect 307334 699014 307372 699066
rect 306836 699012 306892 699014
rect 306916 699012 306972 699014
rect 306996 699012 307052 699014
rect 307076 699012 307132 699014
rect 307156 699012 307212 699014
rect 307236 699012 307292 699014
rect 307316 699012 307372 699014
rect 308586 699896 308642 699952
rect 311990 699216 312046 699272
rect 311990 698944 312046 699000
rect 309138 696804 309140 696824
rect 309140 696804 309192 696824
rect 309192 696804 309194 696824
rect 309138 696768 309194 696804
rect 309046 696632 309102 696688
rect 321650 699216 321706 699272
rect 321558 699080 321614 699136
rect 321650 698964 321706 699000
rect 321650 698944 321652 698964
rect 321652 698944 321704 698964
rect 321704 698944 321706 698964
rect 318614 696768 318670 696824
rect 318798 696632 318854 696688
rect 321558 696632 321614 696688
rect 324836 700698 324892 700700
rect 324916 700698 324972 700700
rect 324996 700698 325052 700700
rect 325076 700698 325132 700700
rect 325156 700698 325212 700700
rect 325236 700698 325292 700700
rect 325316 700698 325372 700700
rect 324836 700646 324874 700698
rect 324874 700646 324886 700698
rect 324886 700646 324892 700698
rect 324916 700646 324938 700698
rect 324938 700646 324950 700698
rect 324950 700646 324972 700698
rect 324996 700646 325002 700698
rect 325002 700646 325014 700698
rect 325014 700646 325052 700698
rect 325076 700646 325078 700698
rect 325078 700646 325130 700698
rect 325130 700646 325132 700698
rect 325156 700646 325194 700698
rect 325194 700646 325206 700698
rect 325206 700646 325212 700698
rect 325236 700646 325258 700698
rect 325258 700646 325270 700698
rect 325270 700646 325292 700698
rect 325316 700646 325322 700698
rect 325322 700646 325334 700698
rect 325334 700646 325372 700698
rect 324836 700644 324892 700646
rect 324916 700644 324972 700646
rect 324996 700644 325052 700646
rect 325076 700644 325132 700646
rect 325156 700644 325212 700646
rect 325236 700644 325292 700646
rect 325316 700644 325372 700646
rect 324836 699610 324892 699612
rect 324916 699610 324972 699612
rect 324996 699610 325052 699612
rect 325076 699610 325132 699612
rect 325156 699610 325212 699612
rect 325236 699610 325292 699612
rect 325316 699610 325372 699612
rect 324836 699558 324874 699610
rect 324874 699558 324886 699610
rect 324886 699558 324892 699610
rect 324916 699558 324938 699610
rect 324938 699558 324950 699610
rect 324950 699558 324972 699610
rect 324996 699558 325002 699610
rect 325002 699558 325014 699610
rect 325014 699558 325052 699610
rect 325076 699558 325078 699610
rect 325078 699558 325130 699610
rect 325130 699558 325132 699610
rect 325156 699558 325194 699610
rect 325194 699558 325206 699610
rect 325206 699558 325212 699610
rect 325236 699558 325258 699610
rect 325258 699558 325270 699610
rect 325270 699558 325292 699610
rect 325316 699558 325322 699610
rect 325322 699558 325334 699610
rect 325334 699558 325372 699610
rect 324836 699556 324892 699558
rect 324916 699556 324972 699558
rect 324996 699556 325052 699558
rect 325076 699556 325132 699558
rect 325156 699556 325212 699558
rect 325236 699556 325292 699558
rect 325316 699556 325372 699558
rect 324836 698522 324892 698524
rect 324916 698522 324972 698524
rect 324996 698522 325052 698524
rect 325076 698522 325132 698524
rect 325156 698522 325212 698524
rect 325236 698522 325292 698524
rect 325316 698522 325372 698524
rect 324836 698470 324874 698522
rect 324874 698470 324886 698522
rect 324886 698470 324892 698522
rect 324916 698470 324938 698522
rect 324938 698470 324950 698522
rect 324950 698470 324972 698522
rect 324996 698470 325002 698522
rect 325002 698470 325014 698522
rect 325014 698470 325052 698522
rect 325076 698470 325078 698522
rect 325078 698470 325130 698522
rect 325130 698470 325132 698522
rect 325156 698470 325194 698522
rect 325194 698470 325206 698522
rect 325206 698470 325212 698522
rect 325236 698470 325258 698522
rect 325258 698470 325270 698522
rect 325270 698470 325292 698522
rect 325316 698470 325322 698522
rect 325322 698470 325334 698522
rect 325334 698470 325372 698522
rect 324836 698468 324892 698470
rect 324916 698468 324972 698470
rect 324996 698468 325052 698470
rect 325076 698468 325132 698470
rect 325156 698468 325212 698470
rect 325236 698468 325292 698470
rect 325316 698468 325372 698470
rect 331034 699216 331090 699272
rect 331310 699216 331366 699272
rect 331126 699116 331128 699136
rect 331128 699116 331180 699136
rect 331180 699116 331182 699136
rect 331126 699080 331182 699116
rect 328458 696632 328514 696688
rect 328366 695952 328422 696008
rect 342836 701242 342892 701244
rect 342916 701242 342972 701244
rect 342996 701242 343052 701244
rect 343076 701242 343132 701244
rect 343156 701242 343212 701244
rect 343236 701242 343292 701244
rect 343316 701242 343372 701244
rect 342836 701190 342874 701242
rect 342874 701190 342886 701242
rect 342886 701190 342892 701242
rect 342916 701190 342938 701242
rect 342938 701190 342950 701242
rect 342950 701190 342972 701242
rect 342996 701190 343002 701242
rect 343002 701190 343014 701242
rect 343014 701190 343052 701242
rect 343076 701190 343078 701242
rect 343078 701190 343130 701242
rect 343130 701190 343132 701242
rect 343156 701190 343194 701242
rect 343194 701190 343206 701242
rect 343206 701190 343212 701242
rect 343236 701190 343258 701242
rect 343258 701190 343270 701242
rect 343270 701190 343292 701242
rect 343316 701190 343322 701242
rect 343322 701190 343334 701242
rect 343334 701190 343372 701242
rect 342836 701188 342892 701190
rect 342916 701188 342972 701190
rect 342996 701188 343052 701190
rect 343076 701188 343132 701190
rect 343156 701188 343212 701190
rect 343236 701188 343292 701190
rect 343316 701188 343372 701190
rect 336922 700984 336978 701040
rect 346306 700440 346362 700496
rect 341614 700304 341670 700360
rect 340694 699216 340750 699272
rect 338118 696768 338174 696824
rect 338026 696632 338082 696688
rect 342836 700154 342892 700156
rect 342916 700154 342972 700156
rect 342996 700154 343052 700156
rect 343076 700154 343132 700156
rect 343156 700154 343212 700156
rect 343236 700154 343292 700156
rect 343316 700154 343372 700156
rect 342836 700102 342874 700154
rect 342874 700102 342886 700154
rect 342886 700102 342892 700154
rect 342916 700102 342938 700154
rect 342938 700102 342950 700154
rect 342950 700102 342972 700154
rect 342996 700102 343002 700154
rect 343002 700102 343014 700154
rect 343014 700102 343052 700154
rect 343076 700102 343078 700154
rect 343078 700102 343130 700154
rect 343130 700102 343132 700154
rect 343156 700102 343194 700154
rect 343194 700102 343206 700154
rect 343206 700102 343212 700154
rect 343236 700102 343258 700154
rect 343258 700102 343270 700154
rect 343270 700102 343292 700154
rect 343316 700102 343322 700154
rect 343322 700102 343334 700154
rect 343334 700102 343372 700154
rect 342836 700100 342892 700102
rect 342916 700100 342972 700102
rect 342996 700100 343052 700102
rect 343076 700100 343132 700102
rect 343156 700100 343212 700102
rect 343236 700100 343292 700102
rect 343316 700100 343372 700102
rect 344926 699216 344982 699272
rect 342836 699066 342892 699068
rect 342916 699066 342972 699068
rect 342996 699066 343052 699068
rect 343076 699066 343132 699068
rect 343156 699066 343212 699068
rect 343236 699066 343292 699068
rect 343316 699066 343372 699068
rect 342836 699014 342874 699066
rect 342874 699014 342886 699066
rect 342886 699014 342892 699066
rect 342916 699014 342938 699066
rect 342938 699014 342950 699066
rect 342950 699014 342972 699066
rect 342996 699014 343002 699066
rect 343002 699014 343014 699066
rect 343014 699014 343052 699066
rect 343076 699014 343078 699066
rect 343078 699014 343130 699066
rect 343130 699014 343132 699066
rect 343156 699014 343194 699066
rect 343194 699014 343206 699066
rect 343206 699014 343212 699066
rect 343236 699014 343258 699066
rect 343258 699014 343270 699066
rect 343270 699014 343292 699066
rect 343316 699014 343322 699066
rect 343322 699014 343334 699066
rect 343334 699014 343372 699066
rect 342836 699012 342892 699014
rect 342916 699012 342972 699014
rect 342996 699012 343052 699014
rect 343076 699012 343132 699014
rect 343156 699012 343212 699014
rect 343236 699012 343292 699014
rect 343316 699012 343372 699014
rect 342626 696788 342682 696824
rect 342626 696768 342628 696788
rect 342628 696768 342680 696788
rect 342680 696768 342682 696788
rect 360836 701786 360892 701788
rect 360916 701786 360972 701788
rect 360996 701786 361052 701788
rect 361076 701786 361132 701788
rect 361156 701786 361212 701788
rect 361236 701786 361292 701788
rect 361316 701786 361372 701788
rect 360836 701734 360874 701786
rect 360874 701734 360886 701786
rect 360886 701734 360892 701786
rect 360916 701734 360938 701786
rect 360938 701734 360950 701786
rect 360950 701734 360972 701786
rect 360996 701734 361002 701786
rect 361002 701734 361014 701786
rect 361014 701734 361052 701786
rect 361076 701734 361078 701786
rect 361078 701734 361130 701786
rect 361130 701734 361132 701786
rect 361156 701734 361194 701786
rect 361194 701734 361206 701786
rect 361206 701734 361212 701786
rect 361236 701734 361258 701786
rect 361258 701734 361270 701786
rect 361270 701734 361292 701786
rect 361316 701734 361322 701786
rect 361322 701734 361334 701786
rect 361334 701734 361372 701786
rect 360836 701732 360892 701734
rect 360916 701732 360972 701734
rect 360996 701732 361052 701734
rect 361076 701732 361132 701734
rect 361156 701732 361212 701734
rect 361236 701732 361292 701734
rect 361316 701732 361372 701734
rect 360836 700698 360892 700700
rect 360916 700698 360972 700700
rect 360996 700698 361052 700700
rect 361076 700698 361132 700700
rect 361156 700698 361212 700700
rect 361236 700698 361292 700700
rect 361316 700698 361372 700700
rect 360836 700646 360874 700698
rect 360874 700646 360886 700698
rect 360886 700646 360892 700698
rect 360916 700646 360938 700698
rect 360938 700646 360950 700698
rect 360950 700646 360972 700698
rect 360996 700646 361002 700698
rect 361002 700646 361014 700698
rect 361014 700646 361052 700698
rect 361076 700646 361078 700698
rect 361078 700646 361130 700698
rect 361130 700646 361132 700698
rect 361156 700646 361194 700698
rect 361194 700646 361206 700698
rect 361206 700646 361212 700698
rect 361236 700646 361258 700698
rect 361258 700646 361270 700698
rect 361270 700646 361292 700698
rect 361316 700646 361322 700698
rect 361322 700646 361334 700698
rect 361334 700646 361372 700698
rect 360836 700644 360892 700646
rect 360916 700644 360972 700646
rect 360996 700644 361052 700646
rect 361076 700644 361132 700646
rect 361156 700644 361212 700646
rect 361236 700644 361292 700646
rect 361316 700644 361372 700646
rect 396836 701786 396892 701788
rect 396916 701786 396972 701788
rect 396996 701786 397052 701788
rect 397076 701786 397132 701788
rect 397156 701786 397212 701788
rect 397236 701786 397292 701788
rect 397316 701786 397372 701788
rect 396836 701734 396874 701786
rect 396874 701734 396886 701786
rect 396886 701734 396892 701786
rect 396916 701734 396938 701786
rect 396938 701734 396950 701786
rect 396950 701734 396972 701786
rect 396996 701734 397002 701786
rect 397002 701734 397014 701786
rect 397014 701734 397052 701786
rect 397076 701734 397078 701786
rect 397078 701734 397130 701786
rect 397130 701734 397132 701786
rect 397156 701734 397194 701786
rect 397194 701734 397206 701786
rect 397206 701734 397212 701786
rect 397236 701734 397258 701786
rect 397258 701734 397270 701786
rect 397270 701734 397292 701786
rect 397316 701734 397322 701786
rect 397322 701734 397334 701786
rect 397334 701734 397372 701786
rect 396836 701732 396892 701734
rect 396916 701732 396972 701734
rect 396996 701732 397052 701734
rect 397076 701732 397132 701734
rect 397156 701732 397212 701734
rect 397236 701732 397292 701734
rect 397316 701732 397372 701734
rect 378836 701242 378892 701244
rect 378916 701242 378972 701244
rect 378996 701242 379052 701244
rect 379076 701242 379132 701244
rect 379156 701242 379212 701244
rect 379236 701242 379292 701244
rect 379316 701242 379372 701244
rect 378836 701190 378874 701242
rect 378874 701190 378886 701242
rect 378886 701190 378892 701242
rect 378916 701190 378938 701242
rect 378938 701190 378950 701242
rect 378950 701190 378972 701242
rect 378996 701190 379002 701242
rect 379002 701190 379014 701242
rect 379014 701190 379052 701242
rect 379076 701190 379078 701242
rect 379078 701190 379130 701242
rect 379130 701190 379132 701242
rect 379156 701190 379194 701242
rect 379194 701190 379206 701242
rect 379206 701190 379212 701242
rect 379236 701190 379258 701242
rect 379258 701190 379270 701242
rect 379270 701190 379292 701242
rect 379316 701190 379322 701242
rect 379322 701190 379334 701242
rect 379334 701190 379372 701242
rect 378836 701188 378892 701190
rect 378916 701188 378972 701190
rect 378996 701188 379052 701190
rect 379076 701188 379132 701190
rect 379156 701188 379212 701190
rect 379236 701188 379292 701190
rect 379316 701188 379372 701190
rect 396836 700698 396892 700700
rect 396916 700698 396972 700700
rect 396996 700698 397052 700700
rect 397076 700698 397132 700700
rect 397156 700698 397212 700700
rect 397236 700698 397292 700700
rect 397316 700698 397372 700700
rect 396836 700646 396874 700698
rect 396874 700646 396886 700698
rect 396886 700646 396892 700698
rect 396916 700646 396938 700698
rect 396938 700646 396950 700698
rect 396950 700646 396972 700698
rect 396996 700646 397002 700698
rect 397002 700646 397014 700698
rect 397014 700646 397052 700698
rect 397076 700646 397078 700698
rect 397078 700646 397130 700698
rect 397130 700646 397132 700698
rect 397156 700646 397194 700698
rect 397194 700646 397206 700698
rect 397206 700646 397212 700698
rect 397236 700646 397258 700698
rect 397258 700646 397270 700698
rect 397270 700646 397292 700698
rect 397316 700646 397322 700698
rect 397322 700646 397334 700698
rect 397334 700646 397372 700698
rect 396836 700644 396892 700646
rect 396916 700644 396972 700646
rect 396996 700644 397052 700646
rect 397076 700644 397132 700646
rect 397156 700644 397212 700646
rect 397236 700644 397292 700646
rect 397316 700644 397372 700646
rect 432836 701786 432892 701788
rect 432916 701786 432972 701788
rect 432996 701786 433052 701788
rect 433076 701786 433132 701788
rect 433156 701786 433212 701788
rect 433236 701786 433292 701788
rect 433316 701786 433372 701788
rect 432836 701734 432874 701786
rect 432874 701734 432886 701786
rect 432886 701734 432892 701786
rect 432916 701734 432938 701786
rect 432938 701734 432950 701786
rect 432950 701734 432972 701786
rect 432996 701734 433002 701786
rect 433002 701734 433014 701786
rect 433014 701734 433052 701786
rect 433076 701734 433078 701786
rect 433078 701734 433130 701786
rect 433130 701734 433132 701786
rect 433156 701734 433194 701786
rect 433194 701734 433206 701786
rect 433206 701734 433212 701786
rect 433236 701734 433258 701786
rect 433258 701734 433270 701786
rect 433270 701734 433292 701786
rect 433316 701734 433322 701786
rect 433322 701734 433334 701786
rect 433334 701734 433372 701786
rect 432836 701732 432892 701734
rect 432916 701732 432972 701734
rect 432996 701732 433052 701734
rect 433076 701732 433132 701734
rect 433156 701732 433212 701734
rect 433236 701732 433292 701734
rect 433316 701732 433372 701734
rect 414836 701242 414892 701244
rect 414916 701242 414972 701244
rect 414996 701242 415052 701244
rect 415076 701242 415132 701244
rect 415156 701242 415212 701244
rect 415236 701242 415292 701244
rect 415316 701242 415372 701244
rect 414836 701190 414874 701242
rect 414874 701190 414886 701242
rect 414886 701190 414892 701242
rect 414916 701190 414938 701242
rect 414938 701190 414950 701242
rect 414950 701190 414972 701242
rect 414996 701190 415002 701242
rect 415002 701190 415014 701242
rect 415014 701190 415052 701242
rect 415076 701190 415078 701242
rect 415078 701190 415130 701242
rect 415130 701190 415132 701242
rect 415156 701190 415194 701242
rect 415194 701190 415206 701242
rect 415206 701190 415212 701242
rect 415236 701190 415258 701242
rect 415258 701190 415270 701242
rect 415270 701190 415292 701242
rect 415316 701190 415322 701242
rect 415322 701190 415334 701242
rect 415334 701190 415372 701242
rect 414836 701188 414892 701190
rect 414916 701188 414972 701190
rect 414996 701188 415052 701190
rect 415076 701188 415132 701190
rect 415156 701188 415212 701190
rect 415236 701188 415292 701190
rect 415316 701188 415372 701190
rect 450836 701242 450892 701244
rect 450916 701242 450972 701244
rect 450996 701242 451052 701244
rect 451076 701242 451132 701244
rect 451156 701242 451212 701244
rect 451236 701242 451292 701244
rect 451316 701242 451372 701244
rect 450836 701190 450874 701242
rect 450874 701190 450886 701242
rect 450886 701190 450892 701242
rect 450916 701190 450938 701242
rect 450938 701190 450950 701242
rect 450950 701190 450972 701242
rect 450996 701190 451002 701242
rect 451002 701190 451014 701242
rect 451014 701190 451052 701242
rect 451076 701190 451078 701242
rect 451078 701190 451130 701242
rect 451130 701190 451132 701242
rect 451156 701190 451194 701242
rect 451194 701190 451206 701242
rect 451206 701190 451212 701242
rect 451236 701190 451258 701242
rect 451258 701190 451270 701242
rect 451270 701190 451292 701242
rect 451316 701190 451322 701242
rect 451322 701190 451334 701242
rect 451334 701190 451372 701242
rect 450836 701188 450892 701190
rect 450916 701188 450972 701190
rect 450996 701188 451052 701190
rect 451076 701188 451132 701190
rect 451156 701188 451212 701190
rect 451236 701188 451292 701190
rect 451316 701188 451372 701190
rect 432836 700698 432892 700700
rect 432916 700698 432972 700700
rect 432996 700698 433052 700700
rect 433076 700698 433132 700700
rect 433156 700698 433212 700700
rect 433236 700698 433292 700700
rect 433316 700698 433372 700700
rect 432836 700646 432874 700698
rect 432874 700646 432886 700698
rect 432886 700646 432892 700698
rect 432916 700646 432938 700698
rect 432938 700646 432950 700698
rect 432950 700646 432972 700698
rect 432996 700646 433002 700698
rect 433002 700646 433014 700698
rect 433014 700646 433052 700698
rect 433076 700646 433078 700698
rect 433078 700646 433130 700698
rect 433130 700646 433132 700698
rect 433156 700646 433194 700698
rect 433194 700646 433206 700698
rect 433206 700646 433212 700698
rect 433236 700646 433258 700698
rect 433258 700646 433270 700698
rect 433270 700646 433292 700698
rect 433316 700646 433322 700698
rect 433322 700646 433334 700698
rect 433334 700646 433372 700698
rect 432836 700644 432892 700646
rect 432916 700644 432972 700646
rect 432996 700644 433052 700646
rect 433076 700644 433132 700646
rect 433156 700644 433212 700646
rect 433236 700644 433292 700646
rect 433316 700644 433372 700646
rect 468836 701786 468892 701788
rect 468916 701786 468972 701788
rect 468996 701786 469052 701788
rect 469076 701786 469132 701788
rect 469156 701786 469212 701788
rect 469236 701786 469292 701788
rect 469316 701786 469372 701788
rect 468836 701734 468874 701786
rect 468874 701734 468886 701786
rect 468886 701734 468892 701786
rect 468916 701734 468938 701786
rect 468938 701734 468950 701786
rect 468950 701734 468972 701786
rect 468996 701734 469002 701786
rect 469002 701734 469014 701786
rect 469014 701734 469052 701786
rect 469076 701734 469078 701786
rect 469078 701734 469130 701786
rect 469130 701734 469132 701786
rect 469156 701734 469194 701786
rect 469194 701734 469206 701786
rect 469206 701734 469212 701786
rect 469236 701734 469258 701786
rect 469258 701734 469270 701786
rect 469270 701734 469292 701786
rect 469316 701734 469322 701786
rect 469322 701734 469334 701786
rect 469334 701734 469372 701786
rect 468836 701732 468892 701734
rect 468916 701732 468972 701734
rect 468996 701732 469052 701734
rect 469076 701732 469132 701734
rect 469156 701732 469212 701734
rect 469236 701732 469292 701734
rect 469316 701732 469372 701734
rect 468836 700698 468892 700700
rect 468916 700698 468972 700700
rect 468996 700698 469052 700700
rect 469076 700698 469132 700700
rect 469156 700698 469212 700700
rect 469236 700698 469292 700700
rect 469316 700698 469372 700700
rect 468836 700646 468874 700698
rect 468874 700646 468886 700698
rect 468886 700646 468892 700698
rect 468916 700646 468938 700698
rect 468938 700646 468950 700698
rect 468950 700646 468972 700698
rect 468996 700646 469002 700698
rect 469002 700646 469014 700698
rect 469014 700646 469052 700698
rect 469076 700646 469078 700698
rect 469078 700646 469130 700698
rect 469130 700646 469132 700698
rect 469156 700646 469194 700698
rect 469194 700646 469206 700698
rect 469206 700646 469212 700698
rect 469236 700646 469258 700698
rect 469258 700646 469270 700698
rect 469270 700646 469292 700698
rect 469316 700646 469322 700698
rect 469322 700646 469334 700698
rect 469334 700646 469372 700698
rect 468836 700644 468892 700646
rect 468916 700644 468972 700646
rect 468996 700644 469052 700646
rect 469076 700644 469132 700646
rect 469156 700644 469212 700646
rect 469236 700644 469292 700646
rect 469316 700644 469372 700646
rect 504836 701786 504892 701788
rect 504916 701786 504972 701788
rect 504996 701786 505052 701788
rect 505076 701786 505132 701788
rect 505156 701786 505212 701788
rect 505236 701786 505292 701788
rect 505316 701786 505372 701788
rect 504836 701734 504874 701786
rect 504874 701734 504886 701786
rect 504886 701734 504892 701786
rect 504916 701734 504938 701786
rect 504938 701734 504950 701786
rect 504950 701734 504972 701786
rect 504996 701734 505002 701786
rect 505002 701734 505014 701786
rect 505014 701734 505052 701786
rect 505076 701734 505078 701786
rect 505078 701734 505130 701786
rect 505130 701734 505132 701786
rect 505156 701734 505194 701786
rect 505194 701734 505206 701786
rect 505206 701734 505212 701786
rect 505236 701734 505258 701786
rect 505258 701734 505270 701786
rect 505270 701734 505292 701786
rect 505316 701734 505322 701786
rect 505322 701734 505334 701786
rect 505334 701734 505372 701786
rect 504836 701732 504892 701734
rect 504916 701732 504972 701734
rect 504996 701732 505052 701734
rect 505076 701732 505132 701734
rect 505156 701732 505212 701734
rect 505236 701732 505292 701734
rect 505316 701732 505372 701734
rect 486836 701242 486892 701244
rect 486916 701242 486972 701244
rect 486996 701242 487052 701244
rect 487076 701242 487132 701244
rect 487156 701242 487212 701244
rect 487236 701242 487292 701244
rect 487316 701242 487372 701244
rect 486836 701190 486874 701242
rect 486874 701190 486886 701242
rect 486886 701190 486892 701242
rect 486916 701190 486938 701242
rect 486938 701190 486950 701242
rect 486950 701190 486972 701242
rect 486996 701190 487002 701242
rect 487002 701190 487014 701242
rect 487014 701190 487052 701242
rect 487076 701190 487078 701242
rect 487078 701190 487130 701242
rect 487130 701190 487132 701242
rect 487156 701190 487194 701242
rect 487194 701190 487206 701242
rect 487206 701190 487212 701242
rect 487236 701190 487258 701242
rect 487258 701190 487270 701242
rect 487270 701190 487292 701242
rect 487316 701190 487322 701242
rect 487322 701190 487334 701242
rect 487334 701190 487372 701242
rect 486836 701188 486892 701190
rect 486916 701188 486972 701190
rect 486996 701188 487052 701190
rect 487076 701188 487132 701190
rect 487156 701188 487212 701190
rect 487236 701188 487292 701190
rect 487316 701188 487372 701190
rect 522836 701242 522892 701244
rect 522916 701242 522972 701244
rect 522996 701242 523052 701244
rect 523076 701242 523132 701244
rect 523156 701242 523212 701244
rect 523236 701242 523292 701244
rect 523316 701242 523372 701244
rect 522836 701190 522874 701242
rect 522874 701190 522886 701242
rect 522886 701190 522892 701242
rect 522916 701190 522938 701242
rect 522938 701190 522950 701242
rect 522950 701190 522972 701242
rect 522996 701190 523002 701242
rect 523002 701190 523014 701242
rect 523014 701190 523052 701242
rect 523076 701190 523078 701242
rect 523078 701190 523130 701242
rect 523130 701190 523132 701242
rect 523156 701190 523194 701242
rect 523194 701190 523206 701242
rect 523206 701190 523212 701242
rect 523236 701190 523258 701242
rect 523258 701190 523270 701242
rect 523270 701190 523292 701242
rect 523316 701190 523322 701242
rect 523322 701190 523334 701242
rect 523334 701190 523372 701242
rect 522836 701188 522892 701190
rect 522916 701188 522972 701190
rect 522996 701188 523052 701190
rect 523076 701188 523132 701190
rect 523156 701188 523212 701190
rect 523236 701188 523292 701190
rect 523316 701188 523372 701190
rect 540836 701786 540892 701788
rect 540916 701786 540972 701788
rect 540996 701786 541052 701788
rect 541076 701786 541132 701788
rect 541156 701786 541212 701788
rect 541236 701786 541292 701788
rect 541316 701786 541372 701788
rect 540836 701734 540874 701786
rect 540874 701734 540886 701786
rect 540886 701734 540892 701786
rect 540916 701734 540938 701786
rect 540938 701734 540950 701786
rect 540950 701734 540972 701786
rect 540996 701734 541002 701786
rect 541002 701734 541014 701786
rect 541014 701734 541052 701786
rect 541076 701734 541078 701786
rect 541078 701734 541130 701786
rect 541130 701734 541132 701786
rect 541156 701734 541194 701786
rect 541194 701734 541206 701786
rect 541206 701734 541212 701786
rect 541236 701734 541258 701786
rect 541258 701734 541270 701786
rect 541270 701734 541292 701786
rect 541316 701734 541322 701786
rect 541322 701734 541334 701786
rect 541334 701734 541372 701786
rect 540836 701732 540892 701734
rect 540916 701732 540972 701734
rect 540996 701732 541052 701734
rect 541076 701732 541132 701734
rect 541156 701732 541212 701734
rect 541236 701732 541292 701734
rect 541316 701732 541372 701734
rect 527178 700848 527234 700904
rect 504836 700698 504892 700700
rect 504916 700698 504972 700700
rect 504996 700698 505052 700700
rect 505076 700698 505132 700700
rect 505156 700698 505212 700700
rect 505236 700698 505292 700700
rect 505316 700698 505372 700700
rect 504836 700646 504874 700698
rect 504874 700646 504886 700698
rect 504886 700646 504892 700698
rect 504916 700646 504938 700698
rect 504938 700646 504950 700698
rect 504950 700646 504972 700698
rect 504996 700646 505002 700698
rect 505002 700646 505014 700698
rect 505014 700646 505052 700698
rect 505076 700646 505078 700698
rect 505078 700646 505130 700698
rect 505130 700646 505132 700698
rect 505156 700646 505194 700698
rect 505194 700646 505206 700698
rect 505206 700646 505212 700698
rect 505236 700646 505258 700698
rect 505258 700646 505270 700698
rect 505270 700646 505292 700698
rect 505316 700646 505322 700698
rect 505322 700646 505334 700698
rect 505334 700646 505372 700698
rect 504836 700644 504892 700646
rect 504916 700644 504972 700646
rect 504996 700644 505052 700646
rect 505076 700644 505132 700646
rect 505156 700644 505212 700646
rect 505236 700644 505292 700646
rect 505316 700644 505372 700646
rect 540836 700698 540892 700700
rect 540916 700698 540972 700700
rect 540996 700698 541052 700700
rect 541076 700698 541132 700700
rect 541156 700698 541212 700700
rect 541236 700698 541292 700700
rect 541316 700698 541372 700700
rect 540836 700646 540874 700698
rect 540874 700646 540886 700698
rect 540886 700646 540892 700698
rect 540916 700646 540938 700698
rect 540938 700646 540950 700698
rect 540950 700646 540972 700698
rect 540996 700646 541002 700698
rect 541002 700646 541014 700698
rect 541014 700646 541052 700698
rect 541076 700646 541078 700698
rect 541078 700646 541130 700698
rect 541130 700646 541132 700698
rect 541156 700646 541194 700698
rect 541194 700646 541206 700698
rect 541206 700646 541212 700698
rect 541236 700646 541258 700698
rect 541258 700646 541270 700698
rect 541270 700646 541292 700698
rect 541316 700646 541322 700698
rect 541322 700646 541334 700698
rect 541334 700646 541372 700698
rect 540836 700644 540892 700646
rect 540916 700644 540972 700646
rect 540996 700644 541052 700646
rect 541076 700644 541132 700646
rect 541156 700644 541212 700646
rect 541236 700644 541292 700646
rect 541316 700644 541372 700646
rect 576836 701786 576892 701788
rect 576916 701786 576972 701788
rect 576996 701786 577052 701788
rect 577076 701786 577132 701788
rect 577156 701786 577212 701788
rect 577236 701786 577292 701788
rect 577316 701786 577372 701788
rect 576836 701734 576874 701786
rect 576874 701734 576886 701786
rect 576886 701734 576892 701786
rect 576916 701734 576938 701786
rect 576938 701734 576950 701786
rect 576950 701734 576972 701786
rect 576996 701734 577002 701786
rect 577002 701734 577014 701786
rect 577014 701734 577052 701786
rect 577076 701734 577078 701786
rect 577078 701734 577130 701786
rect 577130 701734 577132 701786
rect 577156 701734 577194 701786
rect 577194 701734 577206 701786
rect 577206 701734 577212 701786
rect 577236 701734 577258 701786
rect 577258 701734 577270 701786
rect 577270 701734 577292 701786
rect 577316 701734 577322 701786
rect 577322 701734 577334 701786
rect 577334 701734 577372 701786
rect 576836 701732 576892 701734
rect 576916 701732 576972 701734
rect 576996 701732 577052 701734
rect 577076 701732 577132 701734
rect 577156 701732 577212 701734
rect 577236 701732 577292 701734
rect 577316 701732 577372 701734
rect 558836 701242 558892 701244
rect 558916 701242 558972 701244
rect 558996 701242 559052 701244
rect 559076 701242 559132 701244
rect 559156 701242 559212 701244
rect 559236 701242 559292 701244
rect 559316 701242 559372 701244
rect 558836 701190 558874 701242
rect 558874 701190 558886 701242
rect 558886 701190 558892 701242
rect 558916 701190 558938 701242
rect 558938 701190 558950 701242
rect 558950 701190 558972 701242
rect 558996 701190 559002 701242
rect 559002 701190 559014 701242
rect 559014 701190 559052 701242
rect 559076 701190 559078 701242
rect 559078 701190 559130 701242
rect 559130 701190 559132 701242
rect 559156 701190 559194 701242
rect 559194 701190 559206 701242
rect 559206 701190 559212 701242
rect 559236 701190 559258 701242
rect 559258 701190 559270 701242
rect 559270 701190 559292 701242
rect 559316 701190 559322 701242
rect 559322 701190 559334 701242
rect 559334 701190 559372 701242
rect 558836 701188 558892 701190
rect 558916 701188 558972 701190
rect 558996 701188 559052 701190
rect 559076 701188 559132 701190
rect 559156 701188 559212 701190
rect 559236 701188 559292 701190
rect 559316 701188 559372 701190
rect 576836 700698 576892 700700
rect 576916 700698 576972 700700
rect 576996 700698 577052 700700
rect 577076 700698 577132 700700
rect 577156 700698 577212 700700
rect 577236 700698 577292 700700
rect 577316 700698 577372 700700
rect 576836 700646 576874 700698
rect 576874 700646 576886 700698
rect 576886 700646 576892 700698
rect 576916 700646 576938 700698
rect 576938 700646 576950 700698
rect 576950 700646 576972 700698
rect 576996 700646 577002 700698
rect 577002 700646 577014 700698
rect 577014 700646 577052 700698
rect 577076 700646 577078 700698
rect 577078 700646 577130 700698
rect 577130 700646 577132 700698
rect 577156 700646 577194 700698
rect 577194 700646 577206 700698
rect 577206 700646 577212 700698
rect 577236 700646 577258 700698
rect 577258 700646 577270 700698
rect 577270 700646 577292 700698
rect 577316 700646 577322 700698
rect 577322 700646 577334 700698
rect 577334 700646 577372 700698
rect 576836 700644 576892 700646
rect 576916 700644 576972 700646
rect 576996 700644 577052 700646
rect 577076 700644 577132 700646
rect 577156 700644 577212 700646
rect 577236 700644 577292 700646
rect 577316 700644 577372 700646
rect 378836 700154 378892 700156
rect 378916 700154 378972 700156
rect 378996 700154 379052 700156
rect 379076 700154 379132 700156
rect 379156 700154 379212 700156
rect 379236 700154 379292 700156
rect 379316 700154 379372 700156
rect 378836 700102 378874 700154
rect 378874 700102 378886 700154
rect 378886 700102 378892 700154
rect 378916 700102 378938 700154
rect 378938 700102 378950 700154
rect 378950 700102 378972 700154
rect 378996 700102 379002 700154
rect 379002 700102 379014 700154
rect 379014 700102 379052 700154
rect 379076 700102 379078 700154
rect 379078 700102 379130 700154
rect 379130 700102 379132 700154
rect 379156 700102 379194 700154
rect 379194 700102 379206 700154
rect 379206 700102 379212 700154
rect 379236 700102 379258 700154
rect 379258 700102 379270 700154
rect 379270 700102 379292 700154
rect 379316 700102 379322 700154
rect 379322 700102 379334 700154
rect 379334 700102 379372 700154
rect 378836 700100 378892 700102
rect 378916 700100 378972 700102
rect 378996 700100 379052 700102
rect 379076 700100 379132 700102
rect 379156 700100 379212 700102
rect 379236 700100 379292 700102
rect 379316 700100 379372 700102
rect 414836 700154 414892 700156
rect 414916 700154 414972 700156
rect 414996 700154 415052 700156
rect 415076 700154 415132 700156
rect 415156 700154 415212 700156
rect 415236 700154 415292 700156
rect 415316 700154 415372 700156
rect 414836 700102 414874 700154
rect 414874 700102 414886 700154
rect 414886 700102 414892 700154
rect 414916 700102 414938 700154
rect 414938 700102 414950 700154
rect 414950 700102 414972 700154
rect 414996 700102 415002 700154
rect 415002 700102 415014 700154
rect 415014 700102 415052 700154
rect 415076 700102 415078 700154
rect 415078 700102 415130 700154
rect 415130 700102 415132 700154
rect 415156 700102 415194 700154
rect 415194 700102 415206 700154
rect 415206 700102 415212 700154
rect 415236 700102 415258 700154
rect 415258 700102 415270 700154
rect 415270 700102 415292 700154
rect 415316 700102 415322 700154
rect 415322 700102 415334 700154
rect 415334 700102 415372 700154
rect 414836 700100 414892 700102
rect 414916 700100 414972 700102
rect 414996 700100 415052 700102
rect 415076 700100 415132 700102
rect 415156 700100 415212 700102
rect 415236 700100 415292 700102
rect 415316 700100 415372 700102
rect 450836 700154 450892 700156
rect 450916 700154 450972 700156
rect 450996 700154 451052 700156
rect 451076 700154 451132 700156
rect 451156 700154 451212 700156
rect 451236 700154 451292 700156
rect 451316 700154 451372 700156
rect 450836 700102 450874 700154
rect 450874 700102 450886 700154
rect 450886 700102 450892 700154
rect 450916 700102 450938 700154
rect 450938 700102 450950 700154
rect 450950 700102 450972 700154
rect 450996 700102 451002 700154
rect 451002 700102 451014 700154
rect 451014 700102 451052 700154
rect 451076 700102 451078 700154
rect 451078 700102 451130 700154
rect 451130 700102 451132 700154
rect 451156 700102 451194 700154
rect 451194 700102 451206 700154
rect 451206 700102 451212 700154
rect 451236 700102 451258 700154
rect 451258 700102 451270 700154
rect 451270 700102 451292 700154
rect 451316 700102 451322 700154
rect 451322 700102 451334 700154
rect 451334 700102 451372 700154
rect 450836 700100 450892 700102
rect 450916 700100 450972 700102
rect 450996 700100 451052 700102
rect 451076 700100 451132 700102
rect 451156 700100 451212 700102
rect 451236 700100 451292 700102
rect 451316 700100 451372 700102
rect 486836 700154 486892 700156
rect 486916 700154 486972 700156
rect 486996 700154 487052 700156
rect 487076 700154 487132 700156
rect 487156 700154 487212 700156
rect 487236 700154 487292 700156
rect 487316 700154 487372 700156
rect 486836 700102 486874 700154
rect 486874 700102 486886 700154
rect 486886 700102 486892 700154
rect 486916 700102 486938 700154
rect 486938 700102 486950 700154
rect 486950 700102 486972 700154
rect 486996 700102 487002 700154
rect 487002 700102 487014 700154
rect 487014 700102 487052 700154
rect 487076 700102 487078 700154
rect 487078 700102 487130 700154
rect 487130 700102 487132 700154
rect 487156 700102 487194 700154
rect 487194 700102 487206 700154
rect 487206 700102 487212 700154
rect 487236 700102 487258 700154
rect 487258 700102 487270 700154
rect 487270 700102 487292 700154
rect 487316 700102 487322 700154
rect 487322 700102 487334 700154
rect 487334 700102 487372 700154
rect 486836 700100 486892 700102
rect 486916 700100 486972 700102
rect 486996 700100 487052 700102
rect 487076 700100 487132 700102
rect 487156 700100 487212 700102
rect 487236 700100 487292 700102
rect 487316 700100 487372 700102
rect 522836 700154 522892 700156
rect 522916 700154 522972 700156
rect 522996 700154 523052 700156
rect 523076 700154 523132 700156
rect 523156 700154 523212 700156
rect 523236 700154 523292 700156
rect 523316 700154 523372 700156
rect 522836 700102 522874 700154
rect 522874 700102 522886 700154
rect 522886 700102 522892 700154
rect 522916 700102 522938 700154
rect 522938 700102 522950 700154
rect 522950 700102 522972 700154
rect 522996 700102 523002 700154
rect 523002 700102 523014 700154
rect 523014 700102 523052 700154
rect 523076 700102 523078 700154
rect 523078 700102 523130 700154
rect 523130 700102 523132 700154
rect 523156 700102 523194 700154
rect 523194 700102 523206 700154
rect 523206 700102 523212 700154
rect 523236 700102 523258 700154
rect 523258 700102 523270 700154
rect 523270 700102 523292 700154
rect 523316 700102 523322 700154
rect 523322 700102 523334 700154
rect 523334 700102 523372 700154
rect 522836 700100 522892 700102
rect 522916 700100 522972 700102
rect 522996 700100 523052 700102
rect 523076 700100 523132 700102
rect 523156 700100 523212 700102
rect 523236 700100 523292 700102
rect 523316 700100 523372 700102
rect 558836 700154 558892 700156
rect 558916 700154 558972 700156
rect 558996 700154 559052 700156
rect 559076 700154 559132 700156
rect 559156 700154 559212 700156
rect 559236 700154 559292 700156
rect 559316 700154 559372 700156
rect 558836 700102 558874 700154
rect 558874 700102 558886 700154
rect 558886 700102 558892 700154
rect 558916 700102 558938 700154
rect 558938 700102 558950 700154
rect 558950 700102 558972 700154
rect 558996 700102 559002 700154
rect 559002 700102 559014 700154
rect 559014 700102 559052 700154
rect 559076 700102 559078 700154
rect 559078 700102 559130 700154
rect 559130 700102 559132 700154
rect 559156 700102 559194 700154
rect 559194 700102 559206 700154
rect 559206 700102 559212 700154
rect 559236 700102 559258 700154
rect 559258 700102 559270 700154
rect 559270 700102 559292 700154
rect 559316 700102 559322 700154
rect 559322 700102 559334 700154
rect 559334 700102 559372 700154
rect 558836 700100 558892 700102
rect 558916 700100 558972 700102
rect 558996 700100 559052 700102
rect 559076 700100 559132 700102
rect 559156 700100 559212 700102
rect 559236 700100 559292 700102
rect 559316 700100 559372 700102
rect 360836 699610 360892 699612
rect 360916 699610 360972 699612
rect 360996 699610 361052 699612
rect 361076 699610 361132 699612
rect 361156 699610 361212 699612
rect 361236 699610 361292 699612
rect 361316 699610 361372 699612
rect 360836 699558 360874 699610
rect 360874 699558 360886 699610
rect 360886 699558 360892 699610
rect 360916 699558 360938 699610
rect 360938 699558 360950 699610
rect 360950 699558 360972 699610
rect 360996 699558 361002 699610
rect 361002 699558 361014 699610
rect 361014 699558 361052 699610
rect 361076 699558 361078 699610
rect 361078 699558 361130 699610
rect 361130 699558 361132 699610
rect 361156 699558 361194 699610
rect 361194 699558 361206 699610
rect 361206 699558 361212 699610
rect 361236 699558 361258 699610
rect 361258 699558 361270 699610
rect 361270 699558 361292 699610
rect 361316 699558 361322 699610
rect 361322 699558 361334 699610
rect 361334 699558 361372 699610
rect 360836 699556 360892 699558
rect 360916 699556 360972 699558
rect 360996 699556 361052 699558
rect 361076 699556 361132 699558
rect 361156 699556 361212 699558
rect 361236 699556 361292 699558
rect 361316 699556 361372 699558
rect 396836 699610 396892 699612
rect 396916 699610 396972 699612
rect 396996 699610 397052 699612
rect 397076 699610 397132 699612
rect 397156 699610 397212 699612
rect 397236 699610 397292 699612
rect 397316 699610 397372 699612
rect 396836 699558 396874 699610
rect 396874 699558 396886 699610
rect 396886 699558 396892 699610
rect 396916 699558 396938 699610
rect 396938 699558 396950 699610
rect 396950 699558 396972 699610
rect 396996 699558 397002 699610
rect 397002 699558 397014 699610
rect 397014 699558 397052 699610
rect 397076 699558 397078 699610
rect 397078 699558 397130 699610
rect 397130 699558 397132 699610
rect 397156 699558 397194 699610
rect 397194 699558 397206 699610
rect 397206 699558 397212 699610
rect 397236 699558 397258 699610
rect 397258 699558 397270 699610
rect 397270 699558 397292 699610
rect 397316 699558 397322 699610
rect 397322 699558 397334 699610
rect 397334 699558 397372 699610
rect 396836 699556 396892 699558
rect 396916 699556 396972 699558
rect 396996 699556 397052 699558
rect 397076 699556 397132 699558
rect 397156 699556 397212 699558
rect 397236 699556 397292 699558
rect 397316 699556 397372 699558
rect 432836 699610 432892 699612
rect 432916 699610 432972 699612
rect 432996 699610 433052 699612
rect 433076 699610 433132 699612
rect 433156 699610 433212 699612
rect 433236 699610 433292 699612
rect 433316 699610 433372 699612
rect 432836 699558 432874 699610
rect 432874 699558 432886 699610
rect 432886 699558 432892 699610
rect 432916 699558 432938 699610
rect 432938 699558 432950 699610
rect 432950 699558 432972 699610
rect 432996 699558 433002 699610
rect 433002 699558 433014 699610
rect 433014 699558 433052 699610
rect 433076 699558 433078 699610
rect 433078 699558 433130 699610
rect 433130 699558 433132 699610
rect 433156 699558 433194 699610
rect 433194 699558 433206 699610
rect 433206 699558 433212 699610
rect 433236 699558 433258 699610
rect 433258 699558 433270 699610
rect 433270 699558 433292 699610
rect 433316 699558 433322 699610
rect 433322 699558 433334 699610
rect 433334 699558 433372 699610
rect 432836 699556 432892 699558
rect 432916 699556 432972 699558
rect 432996 699556 433052 699558
rect 433076 699556 433132 699558
rect 433156 699556 433212 699558
rect 433236 699556 433292 699558
rect 433316 699556 433372 699558
rect 468836 699610 468892 699612
rect 468916 699610 468972 699612
rect 468996 699610 469052 699612
rect 469076 699610 469132 699612
rect 469156 699610 469212 699612
rect 469236 699610 469292 699612
rect 469316 699610 469372 699612
rect 468836 699558 468874 699610
rect 468874 699558 468886 699610
rect 468886 699558 468892 699610
rect 468916 699558 468938 699610
rect 468938 699558 468950 699610
rect 468950 699558 468972 699610
rect 468996 699558 469002 699610
rect 469002 699558 469014 699610
rect 469014 699558 469052 699610
rect 469076 699558 469078 699610
rect 469078 699558 469130 699610
rect 469130 699558 469132 699610
rect 469156 699558 469194 699610
rect 469194 699558 469206 699610
rect 469206 699558 469212 699610
rect 469236 699558 469258 699610
rect 469258 699558 469270 699610
rect 469270 699558 469292 699610
rect 469316 699558 469322 699610
rect 469322 699558 469334 699610
rect 469334 699558 469372 699610
rect 468836 699556 468892 699558
rect 468916 699556 468972 699558
rect 468996 699556 469052 699558
rect 469076 699556 469132 699558
rect 469156 699556 469212 699558
rect 469236 699556 469292 699558
rect 469316 699556 469372 699558
rect 504836 699610 504892 699612
rect 504916 699610 504972 699612
rect 504996 699610 505052 699612
rect 505076 699610 505132 699612
rect 505156 699610 505212 699612
rect 505236 699610 505292 699612
rect 505316 699610 505372 699612
rect 504836 699558 504874 699610
rect 504874 699558 504886 699610
rect 504886 699558 504892 699610
rect 504916 699558 504938 699610
rect 504938 699558 504950 699610
rect 504950 699558 504972 699610
rect 504996 699558 505002 699610
rect 505002 699558 505014 699610
rect 505014 699558 505052 699610
rect 505076 699558 505078 699610
rect 505078 699558 505130 699610
rect 505130 699558 505132 699610
rect 505156 699558 505194 699610
rect 505194 699558 505206 699610
rect 505206 699558 505212 699610
rect 505236 699558 505258 699610
rect 505258 699558 505270 699610
rect 505270 699558 505292 699610
rect 505316 699558 505322 699610
rect 505322 699558 505334 699610
rect 505334 699558 505372 699610
rect 504836 699556 504892 699558
rect 504916 699556 504972 699558
rect 504996 699556 505052 699558
rect 505076 699556 505132 699558
rect 505156 699556 505212 699558
rect 505236 699556 505292 699558
rect 505316 699556 505372 699558
rect 540836 699610 540892 699612
rect 540916 699610 540972 699612
rect 540996 699610 541052 699612
rect 541076 699610 541132 699612
rect 541156 699610 541212 699612
rect 541236 699610 541292 699612
rect 541316 699610 541372 699612
rect 540836 699558 540874 699610
rect 540874 699558 540886 699610
rect 540886 699558 540892 699610
rect 540916 699558 540938 699610
rect 540938 699558 540950 699610
rect 540950 699558 540972 699610
rect 540996 699558 541002 699610
rect 541002 699558 541014 699610
rect 541014 699558 541052 699610
rect 541076 699558 541078 699610
rect 541078 699558 541130 699610
rect 541130 699558 541132 699610
rect 541156 699558 541194 699610
rect 541194 699558 541206 699610
rect 541206 699558 541212 699610
rect 541236 699558 541258 699610
rect 541258 699558 541270 699610
rect 541270 699558 541292 699610
rect 541316 699558 541322 699610
rect 541322 699558 541334 699610
rect 541334 699558 541372 699610
rect 540836 699556 540892 699558
rect 540916 699556 540972 699558
rect 540996 699556 541052 699558
rect 541076 699556 541132 699558
rect 541156 699556 541212 699558
rect 541236 699556 541292 699558
rect 541316 699556 541372 699558
rect 576836 699610 576892 699612
rect 576916 699610 576972 699612
rect 576996 699610 577052 699612
rect 577076 699610 577132 699612
rect 577156 699610 577212 699612
rect 577236 699610 577292 699612
rect 577316 699610 577372 699612
rect 576836 699558 576874 699610
rect 576874 699558 576886 699610
rect 576886 699558 576892 699610
rect 576916 699558 576938 699610
rect 576938 699558 576950 699610
rect 576950 699558 576972 699610
rect 576996 699558 577002 699610
rect 577002 699558 577014 699610
rect 577014 699558 577052 699610
rect 577076 699558 577078 699610
rect 577078 699558 577130 699610
rect 577130 699558 577132 699610
rect 577156 699558 577194 699610
rect 577194 699558 577206 699610
rect 577206 699558 577212 699610
rect 577236 699558 577258 699610
rect 577258 699558 577270 699610
rect 577270 699558 577292 699610
rect 577316 699558 577322 699610
rect 577322 699558 577334 699610
rect 577334 699558 577372 699610
rect 576836 699556 576892 699558
rect 576916 699556 576972 699558
rect 576996 699556 577052 699558
rect 577076 699556 577132 699558
rect 577156 699556 577212 699558
rect 577236 699556 577292 699558
rect 577316 699556 577372 699558
rect 364338 699236 364394 699272
rect 364338 699216 364340 699236
rect 364340 699216 364392 699236
rect 364392 699216 364394 699236
rect 373906 699236 373962 699272
rect 373906 699216 373908 699236
rect 373908 699216 373960 699236
rect 373960 699216 373962 699236
rect 374090 699216 374146 699272
rect 383566 699236 383622 699272
rect 383566 699216 383568 699236
rect 383568 699216 383620 699236
rect 383620 699216 383622 699236
rect 378836 699066 378892 699068
rect 378916 699066 378972 699068
rect 378996 699066 379052 699068
rect 379076 699066 379132 699068
rect 379156 699066 379212 699068
rect 379236 699066 379292 699068
rect 379316 699066 379372 699068
rect 378836 699014 378874 699066
rect 378874 699014 378886 699066
rect 378886 699014 378892 699066
rect 378916 699014 378938 699066
rect 378938 699014 378950 699066
rect 378950 699014 378972 699066
rect 378996 699014 379002 699066
rect 379002 699014 379014 699066
rect 379014 699014 379052 699066
rect 379076 699014 379078 699066
rect 379078 699014 379130 699066
rect 379130 699014 379132 699066
rect 379156 699014 379194 699066
rect 379194 699014 379206 699066
rect 379206 699014 379212 699066
rect 379236 699014 379258 699066
rect 379258 699014 379270 699066
rect 379270 699014 379292 699066
rect 379316 699014 379322 699066
rect 379322 699014 379334 699066
rect 379334 699014 379372 699066
rect 378836 699012 378892 699014
rect 378916 699012 378972 699014
rect 378996 699012 379052 699014
rect 379076 699012 379132 699014
rect 379156 699012 379212 699014
rect 379236 699012 379292 699014
rect 379316 699012 379372 699014
rect 360836 698522 360892 698524
rect 360916 698522 360972 698524
rect 360996 698522 361052 698524
rect 361076 698522 361132 698524
rect 361156 698522 361212 698524
rect 361236 698522 361292 698524
rect 361316 698522 361372 698524
rect 360836 698470 360874 698522
rect 360874 698470 360886 698522
rect 360886 698470 360892 698522
rect 360916 698470 360938 698522
rect 360938 698470 360950 698522
rect 360950 698470 360972 698522
rect 360996 698470 361002 698522
rect 361002 698470 361014 698522
rect 361014 698470 361052 698522
rect 361076 698470 361078 698522
rect 361078 698470 361130 698522
rect 361130 698470 361132 698522
rect 361156 698470 361194 698522
rect 361194 698470 361206 698522
rect 361206 698470 361212 698522
rect 361236 698470 361258 698522
rect 361258 698470 361270 698522
rect 361270 698470 361292 698522
rect 361316 698470 361322 698522
rect 361322 698470 361334 698522
rect 361334 698470 361372 698522
rect 360836 698468 360892 698470
rect 360916 698468 360972 698470
rect 360996 698468 361052 698470
rect 361076 698468 361132 698470
rect 361156 698468 361212 698470
rect 361236 698468 361292 698470
rect 361316 698468 361372 698470
rect 396836 698522 396892 698524
rect 396916 698522 396972 698524
rect 396996 698522 397052 698524
rect 397076 698522 397132 698524
rect 397156 698522 397212 698524
rect 397236 698522 397292 698524
rect 397316 698522 397372 698524
rect 396836 698470 396874 698522
rect 396874 698470 396886 698522
rect 396886 698470 396892 698522
rect 396916 698470 396938 698522
rect 396938 698470 396950 698522
rect 396950 698470 396972 698522
rect 396996 698470 397002 698522
rect 397002 698470 397014 698522
rect 397014 698470 397052 698522
rect 397076 698470 397078 698522
rect 397078 698470 397130 698522
rect 397130 698470 397132 698522
rect 397156 698470 397194 698522
rect 397194 698470 397206 698522
rect 397206 698470 397212 698522
rect 397236 698470 397258 698522
rect 397258 698470 397270 698522
rect 397270 698470 397292 698522
rect 397316 698470 397322 698522
rect 397322 698470 397334 698522
rect 397334 698470 397372 698522
rect 396836 698468 396892 698470
rect 396916 698468 396972 698470
rect 396996 698468 397052 698470
rect 397076 698468 397132 698470
rect 397156 698468 397212 698470
rect 397236 698468 397292 698470
rect 397316 698468 397372 698470
rect 350446 698164 350448 698184
rect 350448 698164 350500 698184
rect 350500 698164 350502 698184
rect 350446 698128 350502 698164
rect 350722 698128 350778 698184
rect 371882 695952 371938 696008
rect 414836 699066 414892 699068
rect 414916 699066 414972 699068
rect 414996 699066 415052 699068
rect 415076 699066 415132 699068
rect 415156 699066 415212 699068
rect 415236 699066 415292 699068
rect 415316 699066 415372 699068
rect 414836 699014 414874 699066
rect 414874 699014 414886 699066
rect 414886 699014 414892 699066
rect 414916 699014 414938 699066
rect 414938 699014 414950 699066
rect 414950 699014 414972 699066
rect 414996 699014 415002 699066
rect 415002 699014 415014 699066
rect 415014 699014 415052 699066
rect 415076 699014 415078 699066
rect 415078 699014 415130 699066
rect 415130 699014 415132 699066
rect 415156 699014 415194 699066
rect 415194 699014 415206 699066
rect 415206 699014 415212 699066
rect 415236 699014 415258 699066
rect 415258 699014 415270 699066
rect 415270 699014 415292 699066
rect 415316 699014 415322 699066
rect 415322 699014 415334 699066
rect 415334 699014 415372 699066
rect 414836 699012 414892 699014
rect 414916 699012 414972 699014
rect 414996 699012 415052 699014
rect 415076 699012 415132 699014
rect 415156 699012 415212 699014
rect 415236 699012 415292 699014
rect 415316 699012 415372 699014
rect 432836 698522 432892 698524
rect 432916 698522 432972 698524
rect 432996 698522 433052 698524
rect 433076 698522 433132 698524
rect 433156 698522 433212 698524
rect 433236 698522 433292 698524
rect 433316 698522 433372 698524
rect 432836 698470 432874 698522
rect 432874 698470 432886 698522
rect 432886 698470 432892 698522
rect 432916 698470 432938 698522
rect 432938 698470 432950 698522
rect 432950 698470 432972 698522
rect 432996 698470 433002 698522
rect 433002 698470 433014 698522
rect 433014 698470 433052 698522
rect 433076 698470 433078 698522
rect 433078 698470 433130 698522
rect 433130 698470 433132 698522
rect 433156 698470 433194 698522
rect 433194 698470 433206 698522
rect 433206 698470 433212 698522
rect 433236 698470 433258 698522
rect 433258 698470 433270 698522
rect 433270 698470 433292 698522
rect 433316 698470 433322 698522
rect 433322 698470 433334 698522
rect 433334 698470 433372 698522
rect 432836 698468 432892 698470
rect 432916 698468 432972 698470
rect 432996 698468 433052 698470
rect 433076 698468 433132 698470
rect 433156 698468 433212 698470
rect 433236 698468 433292 698470
rect 433316 698468 433372 698470
rect 292670 695816 292726 695872
rect 299386 695816 299442 695872
rect 253938 695680 253994 695736
rect 265622 695680 265678 695736
rect 292486 695680 292542 695736
rect 251086 695544 251142 695600
rect 253846 695544 253902 695600
rect 309230 695680 309286 695736
rect 299386 695544 299442 695600
rect 309138 695544 309194 695600
rect 331218 695680 331274 695736
rect 328366 695544 328422 695600
rect 331126 695544 331182 695600
rect 360290 695680 360346 695736
rect 422206 695816 422262 695872
rect 425058 695816 425114 695872
rect 384946 695680 385002 695736
rect 357438 695544 357494 695600
rect 357622 695544 357678 695600
rect 360106 695544 360162 695600
rect 371882 695544 371938 695600
rect 375378 695544 375434 695600
rect 386602 695680 386658 695736
rect 398746 695680 398802 695736
rect 403070 695680 403126 695736
rect 386510 695544 386566 695600
rect 398930 695544 398986 695600
rect 402978 695544 403034 695600
rect 215298 695408 215354 695464
rect 229006 695408 229062 695464
rect 15382 695272 15438 695328
rect 157062 695272 157118 695328
rect 526258 699216 526314 699272
rect 450836 699066 450892 699068
rect 450916 699066 450972 699068
rect 450996 699066 451052 699068
rect 451076 699066 451132 699068
rect 451156 699066 451212 699068
rect 451236 699066 451292 699068
rect 451316 699066 451372 699068
rect 450836 699014 450874 699066
rect 450874 699014 450886 699066
rect 450886 699014 450892 699066
rect 450916 699014 450938 699066
rect 450938 699014 450950 699066
rect 450950 699014 450972 699066
rect 450996 699014 451002 699066
rect 451002 699014 451014 699066
rect 451014 699014 451052 699066
rect 451076 699014 451078 699066
rect 451078 699014 451130 699066
rect 451130 699014 451132 699066
rect 451156 699014 451194 699066
rect 451194 699014 451206 699066
rect 451206 699014 451212 699066
rect 451236 699014 451258 699066
rect 451258 699014 451270 699066
rect 451270 699014 451292 699066
rect 451316 699014 451322 699066
rect 451322 699014 451334 699066
rect 451334 699014 451372 699066
rect 450836 699012 450892 699014
rect 450916 699012 450972 699014
rect 450996 699012 451052 699014
rect 451076 699012 451132 699014
rect 451156 699012 451212 699014
rect 451236 699012 451292 699014
rect 451316 699012 451372 699014
rect 486836 699066 486892 699068
rect 486916 699066 486972 699068
rect 486996 699066 487052 699068
rect 487076 699066 487132 699068
rect 487156 699066 487212 699068
rect 487236 699066 487292 699068
rect 487316 699066 487372 699068
rect 486836 699014 486874 699066
rect 486874 699014 486886 699066
rect 486886 699014 486892 699066
rect 486916 699014 486938 699066
rect 486938 699014 486950 699066
rect 486950 699014 486972 699066
rect 486996 699014 487002 699066
rect 487002 699014 487014 699066
rect 487014 699014 487052 699066
rect 487076 699014 487078 699066
rect 487078 699014 487130 699066
rect 487130 699014 487132 699066
rect 487156 699014 487194 699066
rect 487194 699014 487206 699066
rect 487206 699014 487212 699066
rect 487236 699014 487258 699066
rect 487258 699014 487270 699066
rect 487270 699014 487292 699066
rect 487316 699014 487322 699066
rect 487322 699014 487334 699066
rect 487334 699014 487372 699066
rect 486836 699012 486892 699014
rect 486916 699012 486972 699014
rect 486996 699012 487052 699014
rect 487076 699012 487132 699014
rect 487156 699012 487212 699014
rect 487236 699012 487292 699014
rect 487316 699012 487372 699014
rect 522836 699066 522892 699068
rect 522916 699066 522972 699068
rect 522996 699066 523052 699068
rect 523076 699066 523132 699068
rect 523156 699066 523212 699068
rect 523236 699066 523292 699068
rect 523316 699066 523372 699068
rect 522836 699014 522874 699066
rect 522874 699014 522886 699066
rect 522886 699014 522892 699066
rect 522916 699014 522938 699066
rect 522938 699014 522950 699066
rect 522950 699014 522972 699066
rect 522996 699014 523002 699066
rect 523002 699014 523014 699066
rect 523014 699014 523052 699066
rect 523076 699014 523078 699066
rect 523078 699014 523130 699066
rect 523130 699014 523132 699066
rect 523156 699014 523194 699066
rect 523194 699014 523206 699066
rect 523206 699014 523212 699066
rect 523236 699014 523258 699066
rect 523258 699014 523270 699066
rect 523270 699014 523292 699066
rect 523316 699014 523322 699066
rect 523322 699014 523334 699066
rect 523334 699014 523372 699066
rect 522836 699012 522892 699014
rect 522916 699012 522972 699014
rect 522996 699012 523052 699014
rect 523076 699012 523132 699014
rect 523156 699012 523212 699014
rect 523236 699012 523292 699014
rect 523316 699012 523372 699014
rect 468836 698522 468892 698524
rect 468916 698522 468972 698524
rect 468996 698522 469052 698524
rect 469076 698522 469132 698524
rect 469156 698522 469212 698524
rect 469236 698522 469292 698524
rect 469316 698522 469372 698524
rect 468836 698470 468874 698522
rect 468874 698470 468886 698522
rect 468886 698470 468892 698522
rect 468916 698470 468938 698522
rect 468938 698470 468950 698522
rect 468950 698470 468972 698522
rect 468996 698470 469002 698522
rect 469002 698470 469014 698522
rect 469014 698470 469052 698522
rect 469076 698470 469078 698522
rect 469078 698470 469130 698522
rect 469130 698470 469132 698522
rect 469156 698470 469194 698522
rect 469194 698470 469206 698522
rect 469206 698470 469212 698522
rect 469236 698470 469258 698522
rect 469258 698470 469270 698522
rect 469270 698470 469292 698522
rect 469316 698470 469322 698522
rect 469322 698470 469334 698522
rect 469334 698470 469372 698522
rect 468836 698468 468892 698470
rect 468916 698468 468972 698470
rect 468996 698468 469052 698470
rect 469076 698468 469132 698470
rect 469156 698468 469212 698470
rect 469236 698468 469292 698470
rect 469316 698468 469372 698470
rect 468482 695952 468538 696008
rect 516782 698672 516838 698728
rect 482926 695952 482982 696008
rect 504836 698522 504892 698524
rect 504916 698522 504972 698524
rect 504996 698522 505052 698524
rect 505076 698522 505132 698524
rect 505156 698522 505212 698524
rect 505236 698522 505292 698524
rect 505316 698522 505372 698524
rect 504836 698470 504874 698522
rect 504874 698470 504886 698522
rect 504886 698470 504892 698522
rect 504916 698470 504938 698522
rect 504938 698470 504950 698522
rect 504950 698470 504972 698522
rect 504996 698470 505002 698522
rect 505002 698470 505014 698522
rect 505014 698470 505052 698522
rect 505076 698470 505078 698522
rect 505078 698470 505130 698522
rect 505130 698470 505132 698522
rect 505156 698470 505194 698522
rect 505194 698470 505206 698522
rect 505206 698470 505212 698522
rect 505236 698470 505258 698522
rect 505258 698470 505270 698522
rect 505270 698470 505292 698522
rect 505316 698470 505322 698522
rect 505322 698470 505334 698522
rect 505334 698470 505372 698522
rect 504836 698468 504892 698470
rect 504916 698468 504972 698470
rect 504996 698468 505052 698470
rect 505076 698468 505132 698470
rect 505156 698468 505212 698470
rect 505236 698468 505292 698470
rect 505316 698468 505372 698470
rect 558836 699066 558892 699068
rect 558916 699066 558972 699068
rect 558996 699066 559052 699068
rect 559076 699066 559132 699068
rect 559156 699066 559212 699068
rect 559236 699066 559292 699068
rect 559316 699066 559372 699068
rect 558836 699014 558874 699066
rect 558874 699014 558886 699066
rect 558886 699014 558892 699066
rect 558916 699014 558938 699066
rect 558938 699014 558950 699066
rect 558950 699014 558972 699066
rect 558996 699014 559002 699066
rect 559002 699014 559014 699066
rect 559014 699014 559052 699066
rect 559076 699014 559078 699066
rect 559078 699014 559130 699066
rect 559130 699014 559132 699066
rect 559156 699014 559194 699066
rect 559194 699014 559206 699066
rect 559206 699014 559212 699066
rect 559236 699014 559258 699066
rect 559258 699014 559270 699066
rect 559270 699014 559292 699066
rect 559316 699014 559322 699066
rect 559322 699014 559334 699066
rect 559334 699014 559372 699066
rect 558836 699012 558892 699014
rect 558916 699012 558972 699014
rect 558996 699012 559052 699014
rect 559076 699012 559132 699014
rect 559156 699012 559212 699014
rect 559236 699012 559292 699014
rect 559316 699012 559372 699014
rect 545118 698808 545174 698864
rect 540836 698522 540892 698524
rect 540916 698522 540972 698524
rect 540996 698522 541052 698524
rect 541076 698522 541132 698524
rect 541156 698522 541212 698524
rect 541236 698522 541292 698524
rect 541316 698522 541372 698524
rect 540836 698470 540874 698522
rect 540874 698470 540886 698522
rect 540886 698470 540892 698522
rect 540916 698470 540938 698522
rect 540938 698470 540950 698522
rect 540950 698470 540972 698522
rect 540996 698470 541002 698522
rect 541002 698470 541014 698522
rect 541014 698470 541052 698522
rect 541076 698470 541078 698522
rect 541078 698470 541130 698522
rect 541130 698470 541132 698522
rect 541156 698470 541194 698522
rect 541194 698470 541206 698522
rect 541206 698470 541212 698522
rect 541236 698470 541258 698522
rect 541258 698470 541270 698522
rect 541270 698470 541292 698522
rect 541316 698470 541322 698522
rect 541322 698470 541334 698522
rect 541334 698470 541372 698522
rect 540836 698468 540892 698470
rect 540916 698468 540972 698470
rect 540996 698468 541052 698470
rect 541076 698468 541132 698470
rect 541156 698468 541212 698470
rect 541236 698468 541292 698470
rect 541316 698468 541372 698470
rect 540426 697040 540482 697096
rect 576836 698522 576892 698524
rect 576916 698522 576972 698524
rect 576996 698522 577052 698524
rect 577076 698522 577132 698524
rect 577156 698522 577212 698524
rect 577236 698522 577292 698524
rect 577316 698522 577372 698524
rect 576836 698470 576874 698522
rect 576874 698470 576886 698522
rect 576886 698470 576892 698522
rect 576916 698470 576938 698522
rect 576938 698470 576950 698522
rect 576950 698470 576972 698522
rect 576996 698470 577002 698522
rect 577002 698470 577014 698522
rect 577014 698470 577052 698522
rect 577076 698470 577078 698522
rect 577078 698470 577130 698522
rect 577130 698470 577132 698522
rect 577156 698470 577194 698522
rect 577194 698470 577206 698522
rect 577206 698470 577212 698522
rect 577236 698470 577258 698522
rect 577258 698470 577270 698522
rect 577270 698470 577292 698522
rect 577316 698470 577322 698522
rect 577322 698470 577334 698522
rect 577334 698470 577372 698522
rect 576836 698468 576892 698470
rect 576916 698468 576972 698470
rect 576996 698468 577052 698470
rect 577076 698468 577132 698470
rect 577156 698468 577212 698470
rect 577236 698468 577292 698470
rect 577316 698468 577372 698470
rect 437294 695816 437350 695872
rect 437478 695816 437534 695872
rect 452566 695680 452622 695736
rect 426530 695544 426586 695600
rect 426898 695544 426954 695600
rect 482926 695680 482982 695736
rect 485778 695680 485834 695736
rect 543830 695700 543886 695736
rect 543830 695680 543832 695700
rect 543832 695680 543884 695700
rect 543884 695680 543886 695700
rect 553214 695680 553270 695736
rect 553398 695680 553454 695736
rect 562322 695716 562324 695736
rect 562324 695716 562376 695736
rect 562376 695716 562378 695736
rect 562322 695680 562378 695716
rect 567106 695716 567108 695736
rect 567108 695716 567160 695736
rect 567160 695716 567162 695736
rect 567106 695680 567162 695716
rect 569314 695680 569370 695736
rect 468482 695544 468538 695600
rect 492586 695544 492642 695600
rect 540978 695544 541034 695600
rect 452566 695408 452622 695464
rect 422206 695272 422262 695328
rect 521382 695272 521438 695328
rect 568486 693776 568542 693832
rect 568486 693368 568542 693424
rect 574742 696904 574798 696960
rect 574650 627952 574706 628008
rect 576122 694320 576178 694376
rect 575478 627952 575534 628008
rect 577962 693912 578018 693968
rect 579618 698028 579620 698048
rect 579620 698028 579672 698048
rect 579672 698028 579674 698048
rect 579618 697992 579674 698028
rect 579434 693504 579490 693560
rect 580262 696088 580318 696144
rect 579802 674600 579858 674656
rect 579618 651072 579674 651128
rect 579802 627680 579858 627736
rect 579618 604152 579674 604208
rect 579526 592456 579582 592512
rect 580170 580760 580226 580816
rect 579618 557232 579674 557288
rect 579434 545536 579490 545592
rect 579802 533840 579858 533896
rect 580078 510312 580134 510368
rect 579342 498616 579398 498672
rect 580170 486784 580226 486840
rect 579250 451696 579306 451752
rect 579986 439864 580042 439920
rect 579618 416472 579674 416528
rect 579618 392944 579674 393000
rect 579158 357856 579214 357912
rect 580170 346024 580226 346080
rect 579066 310800 579122 310856
rect 580170 299104 580226 299160
rect 579618 275712 579674 275768
rect 578974 263880 579030 263936
rect 580170 252184 580226 252240
rect 578882 216960 578938 217016
rect 580170 205264 580226 205320
rect 579618 158344 579674 158400
rect 580170 134816 580226 134872
rect 580170 111424 580226 111480
rect 579894 87896 579950 87952
rect 580906 686296 580962 686352
rect 580906 639376 580962 639432
rect 580814 463392 580870 463448
rect 580722 404776 580778 404832
rect 580722 369552 580778 369608
rect 580630 322632 580686 322688
rect 580538 228792 580594 228848
rect 580446 181872 580502 181928
rect 580630 170040 580686 170096
rect 580354 123120 580410 123176
rect 580262 76200 580318 76256
rect 579802 64504 579858 64560
rect 580170 40976 580226 41032
rect 579618 29280 579674 29336
rect 580170 17584 580226 17640
rect 3146 7148 3148 7168
rect 3148 7148 3200 7168
rect 3200 7148 3202 7168
rect 3146 7112 3202 7148
rect 18836 6010 18892 6012
rect 18916 6010 18972 6012
rect 18996 6010 19052 6012
rect 19076 6010 19132 6012
rect 19156 6010 19212 6012
rect 19236 6010 19292 6012
rect 19316 6010 19372 6012
rect 18836 5958 18874 6010
rect 18874 5958 18886 6010
rect 18886 5958 18892 6010
rect 18916 5958 18938 6010
rect 18938 5958 18950 6010
rect 18950 5958 18972 6010
rect 18996 5958 19002 6010
rect 19002 5958 19014 6010
rect 19014 5958 19052 6010
rect 19076 5958 19078 6010
rect 19078 5958 19130 6010
rect 19130 5958 19132 6010
rect 19156 5958 19194 6010
rect 19194 5958 19206 6010
rect 19206 5958 19212 6010
rect 19236 5958 19258 6010
rect 19258 5958 19270 6010
rect 19270 5958 19292 6010
rect 19316 5958 19322 6010
rect 19322 5958 19334 6010
rect 19334 5958 19372 6010
rect 18836 5956 18892 5958
rect 18916 5956 18972 5958
rect 18996 5956 19052 5958
rect 19076 5956 19132 5958
rect 19156 5956 19212 5958
rect 19236 5956 19292 5958
rect 19316 5956 19372 5958
rect 18836 4922 18892 4924
rect 18916 4922 18972 4924
rect 18996 4922 19052 4924
rect 19076 4922 19132 4924
rect 19156 4922 19212 4924
rect 19236 4922 19292 4924
rect 19316 4922 19372 4924
rect 18836 4870 18874 4922
rect 18874 4870 18886 4922
rect 18886 4870 18892 4922
rect 18916 4870 18938 4922
rect 18938 4870 18950 4922
rect 18950 4870 18972 4922
rect 18996 4870 19002 4922
rect 19002 4870 19014 4922
rect 19014 4870 19052 4922
rect 19076 4870 19078 4922
rect 19078 4870 19130 4922
rect 19130 4870 19132 4922
rect 19156 4870 19194 4922
rect 19194 4870 19206 4922
rect 19206 4870 19212 4922
rect 19236 4870 19258 4922
rect 19258 4870 19270 4922
rect 19270 4870 19292 4922
rect 19316 4870 19322 4922
rect 19322 4870 19334 4922
rect 19334 4870 19372 4922
rect 18836 4868 18892 4870
rect 18916 4868 18972 4870
rect 18996 4868 19052 4870
rect 19076 4868 19132 4870
rect 19156 4868 19212 4870
rect 19236 4868 19292 4870
rect 19316 4868 19372 4870
rect 18836 3834 18892 3836
rect 18916 3834 18972 3836
rect 18996 3834 19052 3836
rect 19076 3834 19132 3836
rect 19156 3834 19212 3836
rect 19236 3834 19292 3836
rect 19316 3834 19372 3836
rect 18836 3782 18874 3834
rect 18874 3782 18886 3834
rect 18886 3782 18892 3834
rect 18916 3782 18938 3834
rect 18938 3782 18950 3834
rect 18950 3782 18972 3834
rect 18996 3782 19002 3834
rect 19002 3782 19014 3834
rect 19014 3782 19052 3834
rect 19076 3782 19078 3834
rect 19078 3782 19130 3834
rect 19130 3782 19132 3834
rect 19156 3782 19194 3834
rect 19194 3782 19206 3834
rect 19206 3782 19212 3834
rect 19236 3782 19258 3834
rect 19258 3782 19270 3834
rect 19270 3782 19292 3834
rect 19316 3782 19322 3834
rect 19322 3782 19334 3834
rect 19334 3782 19372 3834
rect 18836 3780 18892 3782
rect 18916 3780 18972 3782
rect 18996 3780 19052 3782
rect 19076 3780 19132 3782
rect 19156 3780 19212 3782
rect 19236 3780 19292 3782
rect 19316 3780 19372 3782
rect 18836 2746 18892 2748
rect 18916 2746 18972 2748
rect 18996 2746 19052 2748
rect 19076 2746 19132 2748
rect 19156 2746 19212 2748
rect 19236 2746 19292 2748
rect 19316 2746 19372 2748
rect 18836 2694 18874 2746
rect 18874 2694 18886 2746
rect 18886 2694 18892 2746
rect 18916 2694 18938 2746
rect 18938 2694 18950 2746
rect 18950 2694 18972 2746
rect 18996 2694 19002 2746
rect 19002 2694 19014 2746
rect 19014 2694 19052 2746
rect 19076 2694 19078 2746
rect 19078 2694 19130 2746
rect 19130 2694 19132 2746
rect 19156 2694 19194 2746
rect 19194 2694 19206 2746
rect 19206 2694 19212 2746
rect 19236 2694 19258 2746
rect 19258 2694 19270 2746
rect 19270 2694 19292 2746
rect 19316 2694 19322 2746
rect 19322 2694 19334 2746
rect 19334 2694 19372 2746
rect 18836 2692 18892 2694
rect 18916 2692 18972 2694
rect 18996 2692 19052 2694
rect 19076 2692 19132 2694
rect 19156 2692 19212 2694
rect 19236 2692 19292 2694
rect 19316 2692 19372 2694
rect 36836 5466 36892 5468
rect 36916 5466 36972 5468
rect 36996 5466 37052 5468
rect 37076 5466 37132 5468
rect 37156 5466 37212 5468
rect 37236 5466 37292 5468
rect 37316 5466 37372 5468
rect 36836 5414 36874 5466
rect 36874 5414 36886 5466
rect 36886 5414 36892 5466
rect 36916 5414 36938 5466
rect 36938 5414 36950 5466
rect 36950 5414 36972 5466
rect 36996 5414 37002 5466
rect 37002 5414 37014 5466
rect 37014 5414 37052 5466
rect 37076 5414 37078 5466
rect 37078 5414 37130 5466
rect 37130 5414 37132 5466
rect 37156 5414 37194 5466
rect 37194 5414 37206 5466
rect 37206 5414 37212 5466
rect 37236 5414 37258 5466
rect 37258 5414 37270 5466
rect 37270 5414 37292 5466
rect 37316 5414 37322 5466
rect 37322 5414 37334 5466
rect 37334 5414 37372 5466
rect 36836 5412 36892 5414
rect 36916 5412 36972 5414
rect 36996 5412 37052 5414
rect 37076 5412 37132 5414
rect 37156 5412 37212 5414
rect 37236 5412 37292 5414
rect 37316 5412 37372 5414
rect 36836 4378 36892 4380
rect 36916 4378 36972 4380
rect 36996 4378 37052 4380
rect 37076 4378 37132 4380
rect 37156 4378 37212 4380
rect 37236 4378 37292 4380
rect 37316 4378 37372 4380
rect 36836 4326 36874 4378
rect 36874 4326 36886 4378
rect 36886 4326 36892 4378
rect 36916 4326 36938 4378
rect 36938 4326 36950 4378
rect 36950 4326 36972 4378
rect 36996 4326 37002 4378
rect 37002 4326 37014 4378
rect 37014 4326 37052 4378
rect 37076 4326 37078 4378
rect 37078 4326 37130 4378
rect 37130 4326 37132 4378
rect 37156 4326 37194 4378
rect 37194 4326 37206 4378
rect 37206 4326 37212 4378
rect 37236 4326 37258 4378
rect 37258 4326 37270 4378
rect 37270 4326 37292 4378
rect 37316 4326 37322 4378
rect 37322 4326 37334 4378
rect 37334 4326 37372 4378
rect 36836 4324 36892 4326
rect 36916 4324 36972 4326
rect 36996 4324 37052 4326
rect 37076 4324 37132 4326
rect 37156 4324 37212 4326
rect 37236 4324 37292 4326
rect 37316 4324 37372 4326
rect 36836 3290 36892 3292
rect 36916 3290 36972 3292
rect 36996 3290 37052 3292
rect 37076 3290 37132 3292
rect 37156 3290 37212 3292
rect 37236 3290 37292 3292
rect 37316 3290 37372 3292
rect 36836 3238 36874 3290
rect 36874 3238 36886 3290
rect 36886 3238 36892 3290
rect 36916 3238 36938 3290
rect 36938 3238 36950 3290
rect 36950 3238 36972 3290
rect 36996 3238 37002 3290
rect 37002 3238 37014 3290
rect 37014 3238 37052 3290
rect 37076 3238 37078 3290
rect 37078 3238 37130 3290
rect 37130 3238 37132 3290
rect 37156 3238 37194 3290
rect 37194 3238 37206 3290
rect 37206 3238 37212 3290
rect 37236 3238 37258 3290
rect 37258 3238 37270 3290
rect 37270 3238 37292 3290
rect 37316 3238 37322 3290
rect 37322 3238 37334 3290
rect 37334 3238 37372 3290
rect 36836 3236 36892 3238
rect 36916 3236 36972 3238
rect 36996 3236 37052 3238
rect 37076 3236 37132 3238
rect 37156 3236 37212 3238
rect 37236 3236 37292 3238
rect 37316 3236 37372 3238
rect 36836 2202 36892 2204
rect 36916 2202 36972 2204
rect 36996 2202 37052 2204
rect 37076 2202 37132 2204
rect 37156 2202 37212 2204
rect 37236 2202 37292 2204
rect 37316 2202 37372 2204
rect 36836 2150 36874 2202
rect 36874 2150 36886 2202
rect 36886 2150 36892 2202
rect 36916 2150 36938 2202
rect 36938 2150 36950 2202
rect 36950 2150 36972 2202
rect 36996 2150 37002 2202
rect 37002 2150 37014 2202
rect 37014 2150 37052 2202
rect 37076 2150 37078 2202
rect 37078 2150 37130 2202
rect 37130 2150 37132 2202
rect 37156 2150 37194 2202
rect 37194 2150 37206 2202
rect 37206 2150 37212 2202
rect 37236 2150 37258 2202
rect 37258 2150 37270 2202
rect 37270 2150 37292 2202
rect 37316 2150 37322 2202
rect 37322 2150 37334 2202
rect 37334 2150 37372 2202
rect 36836 2148 36892 2150
rect 36916 2148 36972 2150
rect 36996 2148 37052 2150
rect 37076 2148 37132 2150
rect 37156 2148 37212 2150
rect 37236 2148 37292 2150
rect 37316 2148 37372 2150
rect 54836 6010 54892 6012
rect 54916 6010 54972 6012
rect 54996 6010 55052 6012
rect 55076 6010 55132 6012
rect 55156 6010 55212 6012
rect 55236 6010 55292 6012
rect 55316 6010 55372 6012
rect 54836 5958 54874 6010
rect 54874 5958 54886 6010
rect 54886 5958 54892 6010
rect 54916 5958 54938 6010
rect 54938 5958 54950 6010
rect 54950 5958 54972 6010
rect 54996 5958 55002 6010
rect 55002 5958 55014 6010
rect 55014 5958 55052 6010
rect 55076 5958 55078 6010
rect 55078 5958 55130 6010
rect 55130 5958 55132 6010
rect 55156 5958 55194 6010
rect 55194 5958 55206 6010
rect 55206 5958 55212 6010
rect 55236 5958 55258 6010
rect 55258 5958 55270 6010
rect 55270 5958 55292 6010
rect 55316 5958 55322 6010
rect 55322 5958 55334 6010
rect 55334 5958 55372 6010
rect 54836 5956 54892 5958
rect 54916 5956 54972 5958
rect 54996 5956 55052 5958
rect 55076 5956 55132 5958
rect 55156 5956 55212 5958
rect 55236 5956 55292 5958
rect 55316 5956 55372 5958
rect 54836 4922 54892 4924
rect 54916 4922 54972 4924
rect 54996 4922 55052 4924
rect 55076 4922 55132 4924
rect 55156 4922 55212 4924
rect 55236 4922 55292 4924
rect 55316 4922 55372 4924
rect 54836 4870 54874 4922
rect 54874 4870 54886 4922
rect 54886 4870 54892 4922
rect 54916 4870 54938 4922
rect 54938 4870 54950 4922
rect 54950 4870 54972 4922
rect 54996 4870 55002 4922
rect 55002 4870 55014 4922
rect 55014 4870 55052 4922
rect 55076 4870 55078 4922
rect 55078 4870 55130 4922
rect 55130 4870 55132 4922
rect 55156 4870 55194 4922
rect 55194 4870 55206 4922
rect 55206 4870 55212 4922
rect 55236 4870 55258 4922
rect 55258 4870 55270 4922
rect 55270 4870 55292 4922
rect 55316 4870 55322 4922
rect 55322 4870 55334 4922
rect 55334 4870 55372 4922
rect 54836 4868 54892 4870
rect 54916 4868 54972 4870
rect 54996 4868 55052 4870
rect 55076 4868 55132 4870
rect 55156 4868 55212 4870
rect 55236 4868 55292 4870
rect 55316 4868 55372 4870
rect 54836 3834 54892 3836
rect 54916 3834 54972 3836
rect 54996 3834 55052 3836
rect 55076 3834 55132 3836
rect 55156 3834 55212 3836
rect 55236 3834 55292 3836
rect 55316 3834 55372 3836
rect 54836 3782 54874 3834
rect 54874 3782 54886 3834
rect 54886 3782 54892 3834
rect 54916 3782 54938 3834
rect 54938 3782 54950 3834
rect 54950 3782 54972 3834
rect 54996 3782 55002 3834
rect 55002 3782 55014 3834
rect 55014 3782 55052 3834
rect 55076 3782 55078 3834
rect 55078 3782 55130 3834
rect 55130 3782 55132 3834
rect 55156 3782 55194 3834
rect 55194 3782 55206 3834
rect 55206 3782 55212 3834
rect 55236 3782 55258 3834
rect 55258 3782 55270 3834
rect 55270 3782 55292 3834
rect 55316 3782 55322 3834
rect 55322 3782 55334 3834
rect 55334 3782 55372 3834
rect 54836 3780 54892 3782
rect 54916 3780 54972 3782
rect 54996 3780 55052 3782
rect 55076 3780 55132 3782
rect 55156 3780 55212 3782
rect 55236 3780 55292 3782
rect 55316 3780 55372 3782
rect 54836 2746 54892 2748
rect 54916 2746 54972 2748
rect 54996 2746 55052 2748
rect 55076 2746 55132 2748
rect 55156 2746 55212 2748
rect 55236 2746 55292 2748
rect 55316 2746 55372 2748
rect 54836 2694 54874 2746
rect 54874 2694 54886 2746
rect 54886 2694 54892 2746
rect 54916 2694 54938 2746
rect 54938 2694 54950 2746
rect 54950 2694 54972 2746
rect 54996 2694 55002 2746
rect 55002 2694 55014 2746
rect 55014 2694 55052 2746
rect 55076 2694 55078 2746
rect 55078 2694 55130 2746
rect 55130 2694 55132 2746
rect 55156 2694 55194 2746
rect 55194 2694 55206 2746
rect 55206 2694 55212 2746
rect 55236 2694 55258 2746
rect 55258 2694 55270 2746
rect 55270 2694 55292 2746
rect 55316 2694 55322 2746
rect 55322 2694 55334 2746
rect 55334 2694 55372 2746
rect 54836 2692 54892 2694
rect 54916 2692 54972 2694
rect 54996 2692 55052 2694
rect 55076 2692 55132 2694
rect 55156 2692 55212 2694
rect 55236 2692 55292 2694
rect 55316 2692 55372 2694
rect 72836 5466 72892 5468
rect 72916 5466 72972 5468
rect 72996 5466 73052 5468
rect 73076 5466 73132 5468
rect 73156 5466 73212 5468
rect 73236 5466 73292 5468
rect 73316 5466 73372 5468
rect 72836 5414 72874 5466
rect 72874 5414 72886 5466
rect 72886 5414 72892 5466
rect 72916 5414 72938 5466
rect 72938 5414 72950 5466
rect 72950 5414 72972 5466
rect 72996 5414 73002 5466
rect 73002 5414 73014 5466
rect 73014 5414 73052 5466
rect 73076 5414 73078 5466
rect 73078 5414 73130 5466
rect 73130 5414 73132 5466
rect 73156 5414 73194 5466
rect 73194 5414 73206 5466
rect 73206 5414 73212 5466
rect 73236 5414 73258 5466
rect 73258 5414 73270 5466
rect 73270 5414 73292 5466
rect 73316 5414 73322 5466
rect 73322 5414 73334 5466
rect 73334 5414 73372 5466
rect 72836 5412 72892 5414
rect 72916 5412 72972 5414
rect 72996 5412 73052 5414
rect 73076 5412 73132 5414
rect 73156 5412 73212 5414
rect 73236 5412 73292 5414
rect 73316 5412 73372 5414
rect 72836 4378 72892 4380
rect 72916 4378 72972 4380
rect 72996 4378 73052 4380
rect 73076 4378 73132 4380
rect 73156 4378 73212 4380
rect 73236 4378 73292 4380
rect 73316 4378 73372 4380
rect 72836 4326 72874 4378
rect 72874 4326 72886 4378
rect 72886 4326 72892 4378
rect 72916 4326 72938 4378
rect 72938 4326 72950 4378
rect 72950 4326 72972 4378
rect 72996 4326 73002 4378
rect 73002 4326 73014 4378
rect 73014 4326 73052 4378
rect 73076 4326 73078 4378
rect 73078 4326 73130 4378
rect 73130 4326 73132 4378
rect 73156 4326 73194 4378
rect 73194 4326 73206 4378
rect 73206 4326 73212 4378
rect 73236 4326 73258 4378
rect 73258 4326 73270 4378
rect 73270 4326 73292 4378
rect 73316 4326 73322 4378
rect 73322 4326 73334 4378
rect 73334 4326 73372 4378
rect 72836 4324 72892 4326
rect 72916 4324 72972 4326
rect 72996 4324 73052 4326
rect 73076 4324 73132 4326
rect 73156 4324 73212 4326
rect 73236 4324 73292 4326
rect 73316 4324 73372 4326
rect 72836 3290 72892 3292
rect 72916 3290 72972 3292
rect 72996 3290 73052 3292
rect 73076 3290 73132 3292
rect 73156 3290 73212 3292
rect 73236 3290 73292 3292
rect 73316 3290 73372 3292
rect 72836 3238 72874 3290
rect 72874 3238 72886 3290
rect 72886 3238 72892 3290
rect 72916 3238 72938 3290
rect 72938 3238 72950 3290
rect 72950 3238 72972 3290
rect 72996 3238 73002 3290
rect 73002 3238 73014 3290
rect 73014 3238 73052 3290
rect 73076 3238 73078 3290
rect 73078 3238 73130 3290
rect 73130 3238 73132 3290
rect 73156 3238 73194 3290
rect 73194 3238 73206 3290
rect 73206 3238 73212 3290
rect 73236 3238 73258 3290
rect 73258 3238 73270 3290
rect 73270 3238 73292 3290
rect 73316 3238 73322 3290
rect 73322 3238 73334 3290
rect 73334 3238 73372 3290
rect 72836 3236 72892 3238
rect 72916 3236 72972 3238
rect 72996 3236 73052 3238
rect 73076 3236 73132 3238
rect 73156 3236 73212 3238
rect 73236 3236 73292 3238
rect 73316 3236 73372 3238
rect 72836 2202 72892 2204
rect 72916 2202 72972 2204
rect 72996 2202 73052 2204
rect 73076 2202 73132 2204
rect 73156 2202 73212 2204
rect 73236 2202 73292 2204
rect 73316 2202 73372 2204
rect 72836 2150 72874 2202
rect 72874 2150 72886 2202
rect 72886 2150 72892 2202
rect 72916 2150 72938 2202
rect 72938 2150 72950 2202
rect 72950 2150 72972 2202
rect 72996 2150 73002 2202
rect 73002 2150 73014 2202
rect 73014 2150 73052 2202
rect 73076 2150 73078 2202
rect 73078 2150 73130 2202
rect 73130 2150 73132 2202
rect 73156 2150 73194 2202
rect 73194 2150 73206 2202
rect 73206 2150 73212 2202
rect 73236 2150 73258 2202
rect 73258 2150 73270 2202
rect 73270 2150 73292 2202
rect 73316 2150 73322 2202
rect 73322 2150 73334 2202
rect 73334 2150 73372 2202
rect 72836 2148 72892 2150
rect 72916 2148 72972 2150
rect 72996 2148 73052 2150
rect 73076 2148 73132 2150
rect 73156 2148 73212 2150
rect 73236 2148 73292 2150
rect 73316 2148 73372 2150
rect 90836 6010 90892 6012
rect 90916 6010 90972 6012
rect 90996 6010 91052 6012
rect 91076 6010 91132 6012
rect 91156 6010 91212 6012
rect 91236 6010 91292 6012
rect 91316 6010 91372 6012
rect 90836 5958 90874 6010
rect 90874 5958 90886 6010
rect 90886 5958 90892 6010
rect 90916 5958 90938 6010
rect 90938 5958 90950 6010
rect 90950 5958 90972 6010
rect 90996 5958 91002 6010
rect 91002 5958 91014 6010
rect 91014 5958 91052 6010
rect 91076 5958 91078 6010
rect 91078 5958 91130 6010
rect 91130 5958 91132 6010
rect 91156 5958 91194 6010
rect 91194 5958 91206 6010
rect 91206 5958 91212 6010
rect 91236 5958 91258 6010
rect 91258 5958 91270 6010
rect 91270 5958 91292 6010
rect 91316 5958 91322 6010
rect 91322 5958 91334 6010
rect 91334 5958 91372 6010
rect 90836 5956 90892 5958
rect 90916 5956 90972 5958
rect 90996 5956 91052 5958
rect 91076 5956 91132 5958
rect 91156 5956 91212 5958
rect 91236 5956 91292 5958
rect 91316 5956 91372 5958
rect 90836 4922 90892 4924
rect 90916 4922 90972 4924
rect 90996 4922 91052 4924
rect 91076 4922 91132 4924
rect 91156 4922 91212 4924
rect 91236 4922 91292 4924
rect 91316 4922 91372 4924
rect 90836 4870 90874 4922
rect 90874 4870 90886 4922
rect 90886 4870 90892 4922
rect 90916 4870 90938 4922
rect 90938 4870 90950 4922
rect 90950 4870 90972 4922
rect 90996 4870 91002 4922
rect 91002 4870 91014 4922
rect 91014 4870 91052 4922
rect 91076 4870 91078 4922
rect 91078 4870 91130 4922
rect 91130 4870 91132 4922
rect 91156 4870 91194 4922
rect 91194 4870 91206 4922
rect 91206 4870 91212 4922
rect 91236 4870 91258 4922
rect 91258 4870 91270 4922
rect 91270 4870 91292 4922
rect 91316 4870 91322 4922
rect 91322 4870 91334 4922
rect 91334 4870 91372 4922
rect 90836 4868 90892 4870
rect 90916 4868 90972 4870
rect 90996 4868 91052 4870
rect 91076 4868 91132 4870
rect 91156 4868 91212 4870
rect 91236 4868 91292 4870
rect 91316 4868 91372 4870
rect 90836 3834 90892 3836
rect 90916 3834 90972 3836
rect 90996 3834 91052 3836
rect 91076 3834 91132 3836
rect 91156 3834 91212 3836
rect 91236 3834 91292 3836
rect 91316 3834 91372 3836
rect 90836 3782 90874 3834
rect 90874 3782 90886 3834
rect 90886 3782 90892 3834
rect 90916 3782 90938 3834
rect 90938 3782 90950 3834
rect 90950 3782 90972 3834
rect 90996 3782 91002 3834
rect 91002 3782 91014 3834
rect 91014 3782 91052 3834
rect 91076 3782 91078 3834
rect 91078 3782 91130 3834
rect 91130 3782 91132 3834
rect 91156 3782 91194 3834
rect 91194 3782 91206 3834
rect 91206 3782 91212 3834
rect 91236 3782 91258 3834
rect 91258 3782 91270 3834
rect 91270 3782 91292 3834
rect 91316 3782 91322 3834
rect 91322 3782 91334 3834
rect 91334 3782 91372 3834
rect 90836 3780 90892 3782
rect 90916 3780 90972 3782
rect 90996 3780 91052 3782
rect 91076 3780 91132 3782
rect 91156 3780 91212 3782
rect 91236 3780 91292 3782
rect 91316 3780 91372 3782
rect 90836 2746 90892 2748
rect 90916 2746 90972 2748
rect 90996 2746 91052 2748
rect 91076 2746 91132 2748
rect 91156 2746 91212 2748
rect 91236 2746 91292 2748
rect 91316 2746 91372 2748
rect 90836 2694 90874 2746
rect 90874 2694 90886 2746
rect 90886 2694 90892 2746
rect 90916 2694 90938 2746
rect 90938 2694 90950 2746
rect 90950 2694 90972 2746
rect 90996 2694 91002 2746
rect 91002 2694 91014 2746
rect 91014 2694 91052 2746
rect 91076 2694 91078 2746
rect 91078 2694 91130 2746
rect 91130 2694 91132 2746
rect 91156 2694 91194 2746
rect 91194 2694 91206 2746
rect 91206 2694 91212 2746
rect 91236 2694 91258 2746
rect 91258 2694 91270 2746
rect 91270 2694 91292 2746
rect 91316 2694 91322 2746
rect 91322 2694 91334 2746
rect 91334 2694 91372 2746
rect 90836 2692 90892 2694
rect 90916 2692 90972 2694
rect 90996 2692 91052 2694
rect 91076 2692 91132 2694
rect 91156 2692 91212 2694
rect 91236 2692 91292 2694
rect 91316 2692 91372 2694
rect 108836 5466 108892 5468
rect 108916 5466 108972 5468
rect 108996 5466 109052 5468
rect 109076 5466 109132 5468
rect 109156 5466 109212 5468
rect 109236 5466 109292 5468
rect 109316 5466 109372 5468
rect 108836 5414 108874 5466
rect 108874 5414 108886 5466
rect 108886 5414 108892 5466
rect 108916 5414 108938 5466
rect 108938 5414 108950 5466
rect 108950 5414 108972 5466
rect 108996 5414 109002 5466
rect 109002 5414 109014 5466
rect 109014 5414 109052 5466
rect 109076 5414 109078 5466
rect 109078 5414 109130 5466
rect 109130 5414 109132 5466
rect 109156 5414 109194 5466
rect 109194 5414 109206 5466
rect 109206 5414 109212 5466
rect 109236 5414 109258 5466
rect 109258 5414 109270 5466
rect 109270 5414 109292 5466
rect 109316 5414 109322 5466
rect 109322 5414 109334 5466
rect 109334 5414 109372 5466
rect 108836 5412 108892 5414
rect 108916 5412 108972 5414
rect 108996 5412 109052 5414
rect 109076 5412 109132 5414
rect 109156 5412 109212 5414
rect 109236 5412 109292 5414
rect 109316 5412 109372 5414
rect 108836 4378 108892 4380
rect 108916 4378 108972 4380
rect 108996 4378 109052 4380
rect 109076 4378 109132 4380
rect 109156 4378 109212 4380
rect 109236 4378 109292 4380
rect 109316 4378 109372 4380
rect 108836 4326 108874 4378
rect 108874 4326 108886 4378
rect 108886 4326 108892 4378
rect 108916 4326 108938 4378
rect 108938 4326 108950 4378
rect 108950 4326 108972 4378
rect 108996 4326 109002 4378
rect 109002 4326 109014 4378
rect 109014 4326 109052 4378
rect 109076 4326 109078 4378
rect 109078 4326 109130 4378
rect 109130 4326 109132 4378
rect 109156 4326 109194 4378
rect 109194 4326 109206 4378
rect 109206 4326 109212 4378
rect 109236 4326 109258 4378
rect 109258 4326 109270 4378
rect 109270 4326 109292 4378
rect 109316 4326 109322 4378
rect 109322 4326 109334 4378
rect 109334 4326 109372 4378
rect 108836 4324 108892 4326
rect 108916 4324 108972 4326
rect 108996 4324 109052 4326
rect 109076 4324 109132 4326
rect 109156 4324 109212 4326
rect 109236 4324 109292 4326
rect 109316 4324 109372 4326
rect 108836 3290 108892 3292
rect 108916 3290 108972 3292
rect 108996 3290 109052 3292
rect 109076 3290 109132 3292
rect 109156 3290 109212 3292
rect 109236 3290 109292 3292
rect 109316 3290 109372 3292
rect 108836 3238 108874 3290
rect 108874 3238 108886 3290
rect 108886 3238 108892 3290
rect 108916 3238 108938 3290
rect 108938 3238 108950 3290
rect 108950 3238 108972 3290
rect 108996 3238 109002 3290
rect 109002 3238 109014 3290
rect 109014 3238 109052 3290
rect 109076 3238 109078 3290
rect 109078 3238 109130 3290
rect 109130 3238 109132 3290
rect 109156 3238 109194 3290
rect 109194 3238 109206 3290
rect 109206 3238 109212 3290
rect 109236 3238 109258 3290
rect 109258 3238 109270 3290
rect 109270 3238 109292 3290
rect 109316 3238 109322 3290
rect 109322 3238 109334 3290
rect 109334 3238 109372 3290
rect 108836 3236 108892 3238
rect 108916 3236 108972 3238
rect 108996 3236 109052 3238
rect 109076 3236 109132 3238
rect 109156 3236 109212 3238
rect 109236 3236 109292 3238
rect 109316 3236 109372 3238
rect 108836 2202 108892 2204
rect 108916 2202 108972 2204
rect 108996 2202 109052 2204
rect 109076 2202 109132 2204
rect 109156 2202 109212 2204
rect 109236 2202 109292 2204
rect 109316 2202 109372 2204
rect 108836 2150 108874 2202
rect 108874 2150 108886 2202
rect 108886 2150 108892 2202
rect 108916 2150 108938 2202
rect 108938 2150 108950 2202
rect 108950 2150 108972 2202
rect 108996 2150 109002 2202
rect 109002 2150 109014 2202
rect 109014 2150 109052 2202
rect 109076 2150 109078 2202
rect 109078 2150 109130 2202
rect 109130 2150 109132 2202
rect 109156 2150 109194 2202
rect 109194 2150 109206 2202
rect 109206 2150 109212 2202
rect 109236 2150 109258 2202
rect 109258 2150 109270 2202
rect 109270 2150 109292 2202
rect 109316 2150 109322 2202
rect 109322 2150 109334 2202
rect 109334 2150 109372 2202
rect 108836 2148 108892 2150
rect 108916 2148 108972 2150
rect 108996 2148 109052 2150
rect 109076 2148 109132 2150
rect 109156 2148 109212 2150
rect 109236 2148 109292 2150
rect 109316 2148 109372 2150
rect 126836 6010 126892 6012
rect 126916 6010 126972 6012
rect 126996 6010 127052 6012
rect 127076 6010 127132 6012
rect 127156 6010 127212 6012
rect 127236 6010 127292 6012
rect 127316 6010 127372 6012
rect 126836 5958 126874 6010
rect 126874 5958 126886 6010
rect 126886 5958 126892 6010
rect 126916 5958 126938 6010
rect 126938 5958 126950 6010
rect 126950 5958 126972 6010
rect 126996 5958 127002 6010
rect 127002 5958 127014 6010
rect 127014 5958 127052 6010
rect 127076 5958 127078 6010
rect 127078 5958 127130 6010
rect 127130 5958 127132 6010
rect 127156 5958 127194 6010
rect 127194 5958 127206 6010
rect 127206 5958 127212 6010
rect 127236 5958 127258 6010
rect 127258 5958 127270 6010
rect 127270 5958 127292 6010
rect 127316 5958 127322 6010
rect 127322 5958 127334 6010
rect 127334 5958 127372 6010
rect 126836 5956 126892 5958
rect 126916 5956 126972 5958
rect 126996 5956 127052 5958
rect 127076 5956 127132 5958
rect 127156 5956 127212 5958
rect 127236 5956 127292 5958
rect 127316 5956 127372 5958
rect 126836 4922 126892 4924
rect 126916 4922 126972 4924
rect 126996 4922 127052 4924
rect 127076 4922 127132 4924
rect 127156 4922 127212 4924
rect 127236 4922 127292 4924
rect 127316 4922 127372 4924
rect 126836 4870 126874 4922
rect 126874 4870 126886 4922
rect 126886 4870 126892 4922
rect 126916 4870 126938 4922
rect 126938 4870 126950 4922
rect 126950 4870 126972 4922
rect 126996 4870 127002 4922
rect 127002 4870 127014 4922
rect 127014 4870 127052 4922
rect 127076 4870 127078 4922
rect 127078 4870 127130 4922
rect 127130 4870 127132 4922
rect 127156 4870 127194 4922
rect 127194 4870 127206 4922
rect 127206 4870 127212 4922
rect 127236 4870 127258 4922
rect 127258 4870 127270 4922
rect 127270 4870 127292 4922
rect 127316 4870 127322 4922
rect 127322 4870 127334 4922
rect 127334 4870 127372 4922
rect 126836 4868 126892 4870
rect 126916 4868 126972 4870
rect 126996 4868 127052 4870
rect 127076 4868 127132 4870
rect 127156 4868 127212 4870
rect 127236 4868 127292 4870
rect 127316 4868 127372 4870
rect 126836 3834 126892 3836
rect 126916 3834 126972 3836
rect 126996 3834 127052 3836
rect 127076 3834 127132 3836
rect 127156 3834 127212 3836
rect 127236 3834 127292 3836
rect 127316 3834 127372 3836
rect 126836 3782 126874 3834
rect 126874 3782 126886 3834
rect 126886 3782 126892 3834
rect 126916 3782 126938 3834
rect 126938 3782 126950 3834
rect 126950 3782 126972 3834
rect 126996 3782 127002 3834
rect 127002 3782 127014 3834
rect 127014 3782 127052 3834
rect 127076 3782 127078 3834
rect 127078 3782 127130 3834
rect 127130 3782 127132 3834
rect 127156 3782 127194 3834
rect 127194 3782 127206 3834
rect 127206 3782 127212 3834
rect 127236 3782 127258 3834
rect 127258 3782 127270 3834
rect 127270 3782 127292 3834
rect 127316 3782 127322 3834
rect 127322 3782 127334 3834
rect 127334 3782 127372 3834
rect 126836 3780 126892 3782
rect 126916 3780 126972 3782
rect 126996 3780 127052 3782
rect 127076 3780 127132 3782
rect 127156 3780 127212 3782
rect 127236 3780 127292 3782
rect 127316 3780 127372 3782
rect 126836 2746 126892 2748
rect 126916 2746 126972 2748
rect 126996 2746 127052 2748
rect 127076 2746 127132 2748
rect 127156 2746 127212 2748
rect 127236 2746 127292 2748
rect 127316 2746 127372 2748
rect 126836 2694 126874 2746
rect 126874 2694 126886 2746
rect 126886 2694 126892 2746
rect 126916 2694 126938 2746
rect 126938 2694 126950 2746
rect 126950 2694 126972 2746
rect 126996 2694 127002 2746
rect 127002 2694 127014 2746
rect 127014 2694 127052 2746
rect 127076 2694 127078 2746
rect 127078 2694 127130 2746
rect 127130 2694 127132 2746
rect 127156 2694 127194 2746
rect 127194 2694 127206 2746
rect 127206 2694 127212 2746
rect 127236 2694 127258 2746
rect 127258 2694 127270 2746
rect 127270 2694 127292 2746
rect 127316 2694 127322 2746
rect 127322 2694 127334 2746
rect 127334 2694 127372 2746
rect 126836 2692 126892 2694
rect 126916 2692 126972 2694
rect 126996 2692 127052 2694
rect 127076 2692 127132 2694
rect 127156 2692 127212 2694
rect 127236 2692 127292 2694
rect 127316 2692 127372 2694
rect 144836 5466 144892 5468
rect 144916 5466 144972 5468
rect 144996 5466 145052 5468
rect 145076 5466 145132 5468
rect 145156 5466 145212 5468
rect 145236 5466 145292 5468
rect 145316 5466 145372 5468
rect 144836 5414 144874 5466
rect 144874 5414 144886 5466
rect 144886 5414 144892 5466
rect 144916 5414 144938 5466
rect 144938 5414 144950 5466
rect 144950 5414 144972 5466
rect 144996 5414 145002 5466
rect 145002 5414 145014 5466
rect 145014 5414 145052 5466
rect 145076 5414 145078 5466
rect 145078 5414 145130 5466
rect 145130 5414 145132 5466
rect 145156 5414 145194 5466
rect 145194 5414 145206 5466
rect 145206 5414 145212 5466
rect 145236 5414 145258 5466
rect 145258 5414 145270 5466
rect 145270 5414 145292 5466
rect 145316 5414 145322 5466
rect 145322 5414 145334 5466
rect 145334 5414 145372 5466
rect 144836 5412 144892 5414
rect 144916 5412 144972 5414
rect 144996 5412 145052 5414
rect 145076 5412 145132 5414
rect 145156 5412 145212 5414
rect 145236 5412 145292 5414
rect 145316 5412 145372 5414
rect 144836 4378 144892 4380
rect 144916 4378 144972 4380
rect 144996 4378 145052 4380
rect 145076 4378 145132 4380
rect 145156 4378 145212 4380
rect 145236 4378 145292 4380
rect 145316 4378 145372 4380
rect 144836 4326 144874 4378
rect 144874 4326 144886 4378
rect 144886 4326 144892 4378
rect 144916 4326 144938 4378
rect 144938 4326 144950 4378
rect 144950 4326 144972 4378
rect 144996 4326 145002 4378
rect 145002 4326 145014 4378
rect 145014 4326 145052 4378
rect 145076 4326 145078 4378
rect 145078 4326 145130 4378
rect 145130 4326 145132 4378
rect 145156 4326 145194 4378
rect 145194 4326 145206 4378
rect 145206 4326 145212 4378
rect 145236 4326 145258 4378
rect 145258 4326 145270 4378
rect 145270 4326 145292 4378
rect 145316 4326 145322 4378
rect 145322 4326 145334 4378
rect 145334 4326 145372 4378
rect 144836 4324 144892 4326
rect 144916 4324 144972 4326
rect 144996 4324 145052 4326
rect 145076 4324 145132 4326
rect 145156 4324 145212 4326
rect 145236 4324 145292 4326
rect 145316 4324 145372 4326
rect 144836 3290 144892 3292
rect 144916 3290 144972 3292
rect 144996 3290 145052 3292
rect 145076 3290 145132 3292
rect 145156 3290 145212 3292
rect 145236 3290 145292 3292
rect 145316 3290 145372 3292
rect 144836 3238 144874 3290
rect 144874 3238 144886 3290
rect 144886 3238 144892 3290
rect 144916 3238 144938 3290
rect 144938 3238 144950 3290
rect 144950 3238 144972 3290
rect 144996 3238 145002 3290
rect 145002 3238 145014 3290
rect 145014 3238 145052 3290
rect 145076 3238 145078 3290
rect 145078 3238 145130 3290
rect 145130 3238 145132 3290
rect 145156 3238 145194 3290
rect 145194 3238 145206 3290
rect 145206 3238 145212 3290
rect 145236 3238 145258 3290
rect 145258 3238 145270 3290
rect 145270 3238 145292 3290
rect 145316 3238 145322 3290
rect 145322 3238 145334 3290
rect 145334 3238 145372 3290
rect 144836 3236 144892 3238
rect 144916 3236 144972 3238
rect 144996 3236 145052 3238
rect 145076 3236 145132 3238
rect 145156 3236 145212 3238
rect 145236 3236 145292 3238
rect 145316 3236 145372 3238
rect 144836 2202 144892 2204
rect 144916 2202 144972 2204
rect 144996 2202 145052 2204
rect 145076 2202 145132 2204
rect 145156 2202 145212 2204
rect 145236 2202 145292 2204
rect 145316 2202 145372 2204
rect 144836 2150 144874 2202
rect 144874 2150 144886 2202
rect 144886 2150 144892 2202
rect 144916 2150 144938 2202
rect 144938 2150 144950 2202
rect 144950 2150 144972 2202
rect 144996 2150 145002 2202
rect 145002 2150 145014 2202
rect 145014 2150 145052 2202
rect 145076 2150 145078 2202
rect 145078 2150 145130 2202
rect 145130 2150 145132 2202
rect 145156 2150 145194 2202
rect 145194 2150 145206 2202
rect 145206 2150 145212 2202
rect 145236 2150 145258 2202
rect 145258 2150 145270 2202
rect 145270 2150 145292 2202
rect 145316 2150 145322 2202
rect 145322 2150 145334 2202
rect 145334 2150 145372 2202
rect 144836 2148 144892 2150
rect 144916 2148 144972 2150
rect 144996 2148 145052 2150
rect 145076 2148 145132 2150
rect 145156 2148 145212 2150
rect 145236 2148 145292 2150
rect 145316 2148 145372 2150
rect 162836 6010 162892 6012
rect 162916 6010 162972 6012
rect 162996 6010 163052 6012
rect 163076 6010 163132 6012
rect 163156 6010 163212 6012
rect 163236 6010 163292 6012
rect 163316 6010 163372 6012
rect 162836 5958 162874 6010
rect 162874 5958 162886 6010
rect 162886 5958 162892 6010
rect 162916 5958 162938 6010
rect 162938 5958 162950 6010
rect 162950 5958 162972 6010
rect 162996 5958 163002 6010
rect 163002 5958 163014 6010
rect 163014 5958 163052 6010
rect 163076 5958 163078 6010
rect 163078 5958 163130 6010
rect 163130 5958 163132 6010
rect 163156 5958 163194 6010
rect 163194 5958 163206 6010
rect 163206 5958 163212 6010
rect 163236 5958 163258 6010
rect 163258 5958 163270 6010
rect 163270 5958 163292 6010
rect 163316 5958 163322 6010
rect 163322 5958 163334 6010
rect 163334 5958 163372 6010
rect 162836 5956 162892 5958
rect 162916 5956 162972 5958
rect 162996 5956 163052 5958
rect 163076 5956 163132 5958
rect 163156 5956 163212 5958
rect 163236 5956 163292 5958
rect 163316 5956 163372 5958
rect 162836 4922 162892 4924
rect 162916 4922 162972 4924
rect 162996 4922 163052 4924
rect 163076 4922 163132 4924
rect 163156 4922 163212 4924
rect 163236 4922 163292 4924
rect 163316 4922 163372 4924
rect 162836 4870 162874 4922
rect 162874 4870 162886 4922
rect 162886 4870 162892 4922
rect 162916 4870 162938 4922
rect 162938 4870 162950 4922
rect 162950 4870 162972 4922
rect 162996 4870 163002 4922
rect 163002 4870 163014 4922
rect 163014 4870 163052 4922
rect 163076 4870 163078 4922
rect 163078 4870 163130 4922
rect 163130 4870 163132 4922
rect 163156 4870 163194 4922
rect 163194 4870 163206 4922
rect 163206 4870 163212 4922
rect 163236 4870 163258 4922
rect 163258 4870 163270 4922
rect 163270 4870 163292 4922
rect 163316 4870 163322 4922
rect 163322 4870 163334 4922
rect 163334 4870 163372 4922
rect 162836 4868 162892 4870
rect 162916 4868 162972 4870
rect 162996 4868 163052 4870
rect 163076 4868 163132 4870
rect 163156 4868 163212 4870
rect 163236 4868 163292 4870
rect 163316 4868 163372 4870
rect 162836 3834 162892 3836
rect 162916 3834 162972 3836
rect 162996 3834 163052 3836
rect 163076 3834 163132 3836
rect 163156 3834 163212 3836
rect 163236 3834 163292 3836
rect 163316 3834 163372 3836
rect 162836 3782 162874 3834
rect 162874 3782 162886 3834
rect 162886 3782 162892 3834
rect 162916 3782 162938 3834
rect 162938 3782 162950 3834
rect 162950 3782 162972 3834
rect 162996 3782 163002 3834
rect 163002 3782 163014 3834
rect 163014 3782 163052 3834
rect 163076 3782 163078 3834
rect 163078 3782 163130 3834
rect 163130 3782 163132 3834
rect 163156 3782 163194 3834
rect 163194 3782 163206 3834
rect 163206 3782 163212 3834
rect 163236 3782 163258 3834
rect 163258 3782 163270 3834
rect 163270 3782 163292 3834
rect 163316 3782 163322 3834
rect 163322 3782 163334 3834
rect 163334 3782 163372 3834
rect 162836 3780 162892 3782
rect 162916 3780 162972 3782
rect 162996 3780 163052 3782
rect 163076 3780 163132 3782
rect 163156 3780 163212 3782
rect 163236 3780 163292 3782
rect 163316 3780 163372 3782
rect 162836 2746 162892 2748
rect 162916 2746 162972 2748
rect 162996 2746 163052 2748
rect 163076 2746 163132 2748
rect 163156 2746 163212 2748
rect 163236 2746 163292 2748
rect 163316 2746 163372 2748
rect 162836 2694 162874 2746
rect 162874 2694 162886 2746
rect 162886 2694 162892 2746
rect 162916 2694 162938 2746
rect 162938 2694 162950 2746
rect 162950 2694 162972 2746
rect 162996 2694 163002 2746
rect 163002 2694 163014 2746
rect 163014 2694 163052 2746
rect 163076 2694 163078 2746
rect 163078 2694 163130 2746
rect 163130 2694 163132 2746
rect 163156 2694 163194 2746
rect 163194 2694 163206 2746
rect 163206 2694 163212 2746
rect 163236 2694 163258 2746
rect 163258 2694 163270 2746
rect 163270 2694 163292 2746
rect 163316 2694 163322 2746
rect 163322 2694 163334 2746
rect 163334 2694 163372 2746
rect 162836 2692 162892 2694
rect 162916 2692 162972 2694
rect 162996 2692 163052 2694
rect 163076 2692 163132 2694
rect 163156 2692 163212 2694
rect 163236 2692 163292 2694
rect 163316 2692 163372 2694
rect 180836 5466 180892 5468
rect 180916 5466 180972 5468
rect 180996 5466 181052 5468
rect 181076 5466 181132 5468
rect 181156 5466 181212 5468
rect 181236 5466 181292 5468
rect 181316 5466 181372 5468
rect 180836 5414 180874 5466
rect 180874 5414 180886 5466
rect 180886 5414 180892 5466
rect 180916 5414 180938 5466
rect 180938 5414 180950 5466
rect 180950 5414 180972 5466
rect 180996 5414 181002 5466
rect 181002 5414 181014 5466
rect 181014 5414 181052 5466
rect 181076 5414 181078 5466
rect 181078 5414 181130 5466
rect 181130 5414 181132 5466
rect 181156 5414 181194 5466
rect 181194 5414 181206 5466
rect 181206 5414 181212 5466
rect 181236 5414 181258 5466
rect 181258 5414 181270 5466
rect 181270 5414 181292 5466
rect 181316 5414 181322 5466
rect 181322 5414 181334 5466
rect 181334 5414 181372 5466
rect 180836 5412 180892 5414
rect 180916 5412 180972 5414
rect 180996 5412 181052 5414
rect 181076 5412 181132 5414
rect 181156 5412 181212 5414
rect 181236 5412 181292 5414
rect 181316 5412 181372 5414
rect 180836 4378 180892 4380
rect 180916 4378 180972 4380
rect 180996 4378 181052 4380
rect 181076 4378 181132 4380
rect 181156 4378 181212 4380
rect 181236 4378 181292 4380
rect 181316 4378 181372 4380
rect 180836 4326 180874 4378
rect 180874 4326 180886 4378
rect 180886 4326 180892 4378
rect 180916 4326 180938 4378
rect 180938 4326 180950 4378
rect 180950 4326 180972 4378
rect 180996 4326 181002 4378
rect 181002 4326 181014 4378
rect 181014 4326 181052 4378
rect 181076 4326 181078 4378
rect 181078 4326 181130 4378
rect 181130 4326 181132 4378
rect 181156 4326 181194 4378
rect 181194 4326 181206 4378
rect 181206 4326 181212 4378
rect 181236 4326 181258 4378
rect 181258 4326 181270 4378
rect 181270 4326 181292 4378
rect 181316 4326 181322 4378
rect 181322 4326 181334 4378
rect 181334 4326 181372 4378
rect 180836 4324 180892 4326
rect 180916 4324 180972 4326
rect 180996 4324 181052 4326
rect 181076 4324 181132 4326
rect 181156 4324 181212 4326
rect 181236 4324 181292 4326
rect 181316 4324 181372 4326
rect 180836 3290 180892 3292
rect 180916 3290 180972 3292
rect 180996 3290 181052 3292
rect 181076 3290 181132 3292
rect 181156 3290 181212 3292
rect 181236 3290 181292 3292
rect 181316 3290 181372 3292
rect 180836 3238 180874 3290
rect 180874 3238 180886 3290
rect 180886 3238 180892 3290
rect 180916 3238 180938 3290
rect 180938 3238 180950 3290
rect 180950 3238 180972 3290
rect 180996 3238 181002 3290
rect 181002 3238 181014 3290
rect 181014 3238 181052 3290
rect 181076 3238 181078 3290
rect 181078 3238 181130 3290
rect 181130 3238 181132 3290
rect 181156 3238 181194 3290
rect 181194 3238 181206 3290
rect 181206 3238 181212 3290
rect 181236 3238 181258 3290
rect 181258 3238 181270 3290
rect 181270 3238 181292 3290
rect 181316 3238 181322 3290
rect 181322 3238 181334 3290
rect 181334 3238 181372 3290
rect 180836 3236 180892 3238
rect 180916 3236 180972 3238
rect 180996 3236 181052 3238
rect 181076 3236 181132 3238
rect 181156 3236 181212 3238
rect 181236 3236 181292 3238
rect 181316 3236 181372 3238
rect 180836 2202 180892 2204
rect 180916 2202 180972 2204
rect 180996 2202 181052 2204
rect 181076 2202 181132 2204
rect 181156 2202 181212 2204
rect 181236 2202 181292 2204
rect 181316 2202 181372 2204
rect 180836 2150 180874 2202
rect 180874 2150 180886 2202
rect 180886 2150 180892 2202
rect 180916 2150 180938 2202
rect 180938 2150 180950 2202
rect 180950 2150 180972 2202
rect 180996 2150 181002 2202
rect 181002 2150 181014 2202
rect 181014 2150 181052 2202
rect 181076 2150 181078 2202
rect 181078 2150 181130 2202
rect 181130 2150 181132 2202
rect 181156 2150 181194 2202
rect 181194 2150 181206 2202
rect 181206 2150 181212 2202
rect 181236 2150 181258 2202
rect 181258 2150 181270 2202
rect 181270 2150 181292 2202
rect 181316 2150 181322 2202
rect 181322 2150 181334 2202
rect 181334 2150 181372 2202
rect 180836 2148 180892 2150
rect 180916 2148 180972 2150
rect 180996 2148 181052 2150
rect 181076 2148 181132 2150
rect 181156 2148 181212 2150
rect 181236 2148 181292 2150
rect 181316 2148 181372 2150
rect 198836 6010 198892 6012
rect 198916 6010 198972 6012
rect 198996 6010 199052 6012
rect 199076 6010 199132 6012
rect 199156 6010 199212 6012
rect 199236 6010 199292 6012
rect 199316 6010 199372 6012
rect 198836 5958 198874 6010
rect 198874 5958 198886 6010
rect 198886 5958 198892 6010
rect 198916 5958 198938 6010
rect 198938 5958 198950 6010
rect 198950 5958 198972 6010
rect 198996 5958 199002 6010
rect 199002 5958 199014 6010
rect 199014 5958 199052 6010
rect 199076 5958 199078 6010
rect 199078 5958 199130 6010
rect 199130 5958 199132 6010
rect 199156 5958 199194 6010
rect 199194 5958 199206 6010
rect 199206 5958 199212 6010
rect 199236 5958 199258 6010
rect 199258 5958 199270 6010
rect 199270 5958 199292 6010
rect 199316 5958 199322 6010
rect 199322 5958 199334 6010
rect 199334 5958 199372 6010
rect 198836 5956 198892 5958
rect 198916 5956 198972 5958
rect 198996 5956 199052 5958
rect 199076 5956 199132 5958
rect 199156 5956 199212 5958
rect 199236 5956 199292 5958
rect 199316 5956 199372 5958
rect 198836 4922 198892 4924
rect 198916 4922 198972 4924
rect 198996 4922 199052 4924
rect 199076 4922 199132 4924
rect 199156 4922 199212 4924
rect 199236 4922 199292 4924
rect 199316 4922 199372 4924
rect 198836 4870 198874 4922
rect 198874 4870 198886 4922
rect 198886 4870 198892 4922
rect 198916 4870 198938 4922
rect 198938 4870 198950 4922
rect 198950 4870 198972 4922
rect 198996 4870 199002 4922
rect 199002 4870 199014 4922
rect 199014 4870 199052 4922
rect 199076 4870 199078 4922
rect 199078 4870 199130 4922
rect 199130 4870 199132 4922
rect 199156 4870 199194 4922
rect 199194 4870 199206 4922
rect 199206 4870 199212 4922
rect 199236 4870 199258 4922
rect 199258 4870 199270 4922
rect 199270 4870 199292 4922
rect 199316 4870 199322 4922
rect 199322 4870 199334 4922
rect 199334 4870 199372 4922
rect 198836 4868 198892 4870
rect 198916 4868 198972 4870
rect 198996 4868 199052 4870
rect 199076 4868 199132 4870
rect 199156 4868 199212 4870
rect 199236 4868 199292 4870
rect 199316 4868 199372 4870
rect 198836 3834 198892 3836
rect 198916 3834 198972 3836
rect 198996 3834 199052 3836
rect 199076 3834 199132 3836
rect 199156 3834 199212 3836
rect 199236 3834 199292 3836
rect 199316 3834 199372 3836
rect 198836 3782 198874 3834
rect 198874 3782 198886 3834
rect 198886 3782 198892 3834
rect 198916 3782 198938 3834
rect 198938 3782 198950 3834
rect 198950 3782 198972 3834
rect 198996 3782 199002 3834
rect 199002 3782 199014 3834
rect 199014 3782 199052 3834
rect 199076 3782 199078 3834
rect 199078 3782 199130 3834
rect 199130 3782 199132 3834
rect 199156 3782 199194 3834
rect 199194 3782 199206 3834
rect 199206 3782 199212 3834
rect 199236 3782 199258 3834
rect 199258 3782 199270 3834
rect 199270 3782 199292 3834
rect 199316 3782 199322 3834
rect 199322 3782 199334 3834
rect 199334 3782 199372 3834
rect 198836 3780 198892 3782
rect 198916 3780 198972 3782
rect 198996 3780 199052 3782
rect 199076 3780 199132 3782
rect 199156 3780 199212 3782
rect 199236 3780 199292 3782
rect 199316 3780 199372 3782
rect 198836 2746 198892 2748
rect 198916 2746 198972 2748
rect 198996 2746 199052 2748
rect 199076 2746 199132 2748
rect 199156 2746 199212 2748
rect 199236 2746 199292 2748
rect 199316 2746 199372 2748
rect 198836 2694 198874 2746
rect 198874 2694 198886 2746
rect 198886 2694 198892 2746
rect 198916 2694 198938 2746
rect 198938 2694 198950 2746
rect 198950 2694 198972 2746
rect 198996 2694 199002 2746
rect 199002 2694 199014 2746
rect 199014 2694 199052 2746
rect 199076 2694 199078 2746
rect 199078 2694 199130 2746
rect 199130 2694 199132 2746
rect 199156 2694 199194 2746
rect 199194 2694 199206 2746
rect 199206 2694 199212 2746
rect 199236 2694 199258 2746
rect 199258 2694 199270 2746
rect 199270 2694 199292 2746
rect 199316 2694 199322 2746
rect 199322 2694 199334 2746
rect 199334 2694 199372 2746
rect 198836 2692 198892 2694
rect 198916 2692 198972 2694
rect 198996 2692 199052 2694
rect 199076 2692 199132 2694
rect 199156 2692 199212 2694
rect 199236 2692 199292 2694
rect 199316 2692 199372 2694
rect 216836 5466 216892 5468
rect 216916 5466 216972 5468
rect 216996 5466 217052 5468
rect 217076 5466 217132 5468
rect 217156 5466 217212 5468
rect 217236 5466 217292 5468
rect 217316 5466 217372 5468
rect 216836 5414 216874 5466
rect 216874 5414 216886 5466
rect 216886 5414 216892 5466
rect 216916 5414 216938 5466
rect 216938 5414 216950 5466
rect 216950 5414 216972 5466
rect 216996 5414 217002 5466
rect 217002 5414 217014 5466
rect 217014 5414 217052 5466
rect 217076 5414 217078 5466
rect 217078 5414 217130 5466
rect 217130 5414 217132 5466
rect 217156 5414 217194 5466
rect 217194 5414 217206 5466
rect 217206 5414 217212 5466
rect 217236 5414 217258 5466
rect 217258 5414 217270 5466
rect 217270 5414 217292 5466
rect 217316 5414 217322 5466
rect 217322 5414 217334 5466
rect 217334 5414 217372 5466
rect 216836 5412 216892 5414
rect 216916 5412 216972 5414
rect 216996 5412 217052 5414
rect 217076 5412 217132 5414
rect 217156 5412 217212 5414
rect 217236 5412 217292 5414
rect 217316 5412 217372 5414
rect 216836 4378 216892 4380
rect 216916 4378 216972 4380
rect 216996 4378 217052 4380
rect 217076 4378 217132 4380
rect 217156 4378 217212 4380
rect 217236 4378 217292 4380
rect 217316 4378 217372 4380
rect 216836 4326 216874 4378
rect 216874 4326 216886 4378
rect 216886 4326 216892 4378
rect 216916 4326 216938 4378
rect 216938 4326 216950 4378
rect 216950 4326 216972 4378
rect 216996 4326 217002 4378
rect 217002 4326 217014 4378
rect 217014 4326 217052 4378
rect 217076 4326 217078 4378
rect 217078 4326 217130 4378
rect 217130 4326 217132 4378
rect 217156 4326 217194 4378
rect 217194 4326 217206 4378
rect 217206 4326 217212 4378
rect 217236 4326 217258 4378
rect 217258 4326 217270 4378
rect 217270 4326 217292 4378
rect 217316 4326 217322 4378
rect 217322 4326 217334 4378
rect 217334 4326 217372 4378
rect 216836 4324 216892 4326
rect 216916 4324 216972 4326
rect 216996 4324 217052 4326
rect 217076 4324 217132 4326
rect 217156 4324 217212 4326
rect 217236 4324 217292 4326
rect 217316 4324 217372 4326
rect 216836 3290 216892 3292
rect 216916 3290 216972 3292
rect 216996 3290 217052 3292
rect 217076 3290 217132 3292
rect 217156 3290 217212 3292
rect 217236 3290 217292 3292
rect 217316 3290 217372 3292
rect 216836 3238 216874 3290
rect 216874 3238 216886 3290
rect 216886 3238 216892 3290
rect 216916 3238 216938 3290
rect 216938 3238 216950 3290
rect 216950 3238 216972 3290
rect 216996 3238 217002 3290
rect 217002 3238 217014 3290
rect 217014 3238 217052 3290
rect 217076 3238 217078 3290
rect 217078 3238 217130 3290
rect 217130 3238 217132 3290
rect 217156 3238 217194 3290
rect 217194 3238 217206 3290
rect 217206 3238 217212 3290
rect 217236 3238 217258 3290
rect 217258 3238 217270 3290
rect 217270 3238 217292 3290
rect 217316 3238 217322 3290
rect 217322 3238 217334 3290
rect 217334 3238 217372 3290
rect 216836 3236 216892 3238
rect 216916 3236 216972 3238
rect 216996 3236 217052 3238
rect 217076 3236 217132 3238
rect 217156 3236 217212 3238
rect 217236 3236 217292 3238
rect 217316 3236 217372 3238
rect 216836 2202 216892 2204
rect 216916 2202 216972 2204
rect 216996 2202 217052 2204
rect 217076 2202 217132 2204
rect 217156 2202 217212 2204
rect 217236 2202 217292 2204
rect 217316 2202 217372 2204
rect 216836 2150 216874 2202
rect 216874 2150 216886 2202
rect 216886 2150 216892 2202
rect 216916 2150 216938 2202
rect 216938 2150 216950 2202
rect 216950 2150 216972 2202
rect 216996 2150 217002 2202
rect 217002 2150 217014 2202
rect 217014 2150 217052 2202
rect 217076 2150 217078 2202
rect 217078 2150 217130 2202
rect 217130 2150 217132 2202
rect 217156 2150 217194 2202
rect 217194 2150 217206 2202
rect 217206 2150 217212 2202
rect 217236 2150 217258 2202
rect 217258 2150 217270 2202
rect 217270 2150 217292 2202
rect 217316 2150 217322 2202
rect 217322 2150 217334 2202
rect 217334 2150 217372 2202
rect 216836 2148 216892 2150
rect 216916 2148 216972 2150
rect 216996 2148 217052 2150
rect 217076 2148 217132 2150
rect 217156 2148 217212 2150
rect 217236 2148 217292 2150
rect 217316 2148 217372 2150
rect 234836 6010 234892 6012
rect 234916 6010 234972 6012
rect 234996 6010 235052 6012
rect 235076 6010 235132 6012
rect 235156 6010 235212 6012
rect 235236 6010 235292 6012
rect 235316 6010 235372 6012
rect 234836 5958 234874 6010
rect 234874 5958 234886 6010
rect 234886 5958 234892 6010
rect 234916 5958 234938 6010
rect 234938 5958 234950 6010
rect 234950 5958 234972 6010
rect 234996 5958 235002 6010
rect 235002 5958 235014 6010
rect 235014 5958 235052 6010
rect 235076 5958 235078 6010
rect 235078 5958 235130 6010
rect 235130 5958 235132 6010
rect 235156 5958 235194 6010
rect 235194 5958 235206 6010
rect 235206 5958 235212 6010
rect 235236 5958 235258 6010
rect 235258 5958 235270 6010
rect 235270 5958 235292 6010
rect 235316 5958 235322 6010
rect 235322 5958 235334 6010
rect 235334 5958 235372 6010
rect 234836 5956 234892 5958
rect 234916 5956 234972 5958
rect 234996 5956 235052 5958
rect 235076 5956 235132 5958
rect 235156 5956 235212 5958
rect 235236 5956 235292 5958
rect 235316 5956 235372 5958
rect 234836 4922 234892 4924
rect 234916 4922 234972 4924
rect 234996 4922 235052 4924
rect 235076 4922 235132 4924
rect 235156 4922 235212 4924
rect 235236 4922 235292 4924
rect 235316 4922 235372 4924
rect 234836 4870 234874 4922
rect 234874 4870 234886 4922
rect 234886 4870 234892 4922
rect 234916 4870 234938 4922
rect 234938 4870 234950 4922
rect 234950 4870 234972 4922
rect 234996 4870 235002 4922
rect 235002 4870 235014 4922
rect 235014 4870 235052 4922
rect 235076 4870 235078 4922
rect 235078 4870 235130 4922
rect 235130 4870 235132 4922
rect 235156 4870 235194 4922
rect 235194 4870 235206 4922
rect 235206 4870 235212 4922
rect 235236 4870 235258 4922
rect 235258 4870 235270 4922
rect 235270 4870 235292 4922
rect 235316 4870 235322 4922
rect 235322 4870 235334 4922
rect 235334 4870 235372 4922
rect 234836 4868 234892 4870
rect 234916 4868 234972 4870
rect 234996 4868 235052 4870
rect 235076 4868 235132 4870
rect 235156 4868 235212 4870
rect 235236 4868 235292 4870
rect 235316 4868 235372 4870
rect 234836 3834 234892 3836
rect 234916 3834 234972 3836
rect 234996 3834 235052 3836
rect 235076 3834 235132 3836
rect 235156 3834 235212 3836
rect 235236 3834 235292 3836
rect 235316 3834 235372 3836
rect 234836 3782 234874 3834
rect 234874 3782 234886 3834
rect 234886 3782 234892 3834
rect 234916 3782 234938 3834
rect 234938 3782 234950 3834
rect 234950 3782 234972 3834
rect 234996 3782 235002 3834
rect 235002 3782 235014 3834
rect 235014 3782 235052 3834
rect 235076 3782 235078 3834
rect 235078 3782 235130 3834
rect 235130 3782 235132 3834
rect 235156 3782 235194 3834
rect 235194 3782 235206 3834
rect 235206 3782 235212 3834
rect 235236 3782 235258 3834
rect 235258 3782 235270 3834
rect 235270 3782 235292 3834
rect 235316 3782 235322 3834
rect 235322 3782 235334 3834
rect 235334 3782 235372 3834
rect 234836 3780 234892 3782
rect 234916 3780 234972 3782
rect 234996 3780 235052 3782
rect 235076 3780 235132 3782
rect 235156 3780 235212 3782
rect 235236 3780 235292 3782
rect 235316 3780 235372 3782
rect 234836 2746 234892 2748
rect 234916 2746 234972 2748
rect 234996 2746 235052 2748
rect 235076 2746 235132 2748
rect 235156 2746 235212 2748
rect 235236 2746 235292 2748
rect 235316 2746 235372 2748
rect 234836 2694 234874 2746
rect 234874 2694 234886 2746
rect 234886 2694 234892 2746
rect 234916 2694 234938 2746
rect 234938 2694 234950 2746
rect 234950 2694 234972 2746
rect 234996 2694 235002 2746
rect 235002 2694 235014 2746
rect 235014 2694 235052 2746
rect 235076 2694 235078 2746
rect 235078 2694 235130 2746
rect 235130 2694 235132 2746
rect 235156 2694 235194 2746
rect 235194 2694 235206 2746
rect 235206 2694 235212 2746
rect 235236 2694 235258 2746
rect 235258 2694 235270 2746
rect 235270 2694 235292 2746
rect 235316 2694 235322 2746
rect 235322 2694 235334 2746
rect 235334 2694 235372 2746
rect 234836 2692 234892 2694
rect 234916 2692 234972 2694
rect 234996 2692 235052 2694
rect 235076 2692 235132 2694
rect 235156 2692 235212 2694
rect 235236 2692 235292 2694
rect 235316 2692 235372 2694
rect 252836 5466 252892 5468
rect 252916 5466 252972 5468
rect 252996 5466 253052 5468
rect 253076 5466 253132 5468
rect 253156 5466 253212 5468
rect 253236 5466 253292 5468
rect 253316 5466 253372 5468
rect 252836 5414 252874 5466
rect 252874 5414 252886 5466
rect 252886 5414 252892 5466
rect 252916 5414 252938 5466
rect 252938 5414 252950 5466
rect 252950 5414 252972 5466
rect 252996 5414 253002 5466
rect 253002 5414 253014 5466
rect 253014 5414 253052 5466
rect 253076 5414 253078 5466
rect 253078 5414 253130 5466
rect 253130 5414 253132 5466
rect 253156 5414 253194 5466
rect 253194 5414 253206 5466
rect 253206 5414 253212 5466
rect 253236 5414 253258 5466
rect 253258 5414 253270 5466
rect 253270 5414 253292 5466
rect 253316 5414 253322 5466
rect 253322 5414 253334 5466
rect 253334 5414 253372 5466
rect 252836 5412 252892 5414
rect 252916 5412 252972 5414
rect 252996 5412 253052 5414
rect 253076 5412 253132 5414
rect 253156 5412 253212 5414
rect 253236 5412 253292 5414
rect 253316 5412 253372 5414
rect 252836 4378 252892 4380
rect 252916 4378 252972 4380
rect 252996 4378 253052 4380
rect 253076 4378 253132 4380
rect 253156 4378 253212 4380
rect 253236 4378 253292 4380
rect 253316 4378 253372 4380
rect 252836 4326 252874 4378
rect 252874 4326 252886 4378
rect 252886 4326 252892 4378
rect 252916 4326 252938 4378
rect 252938 4326 252950 4378
rect 252950 4326 252972 4378
rect 252996 4326 253002 4378
rect 253002 4326 253014 4378
rect 253014 4326 253052 4378
rect 253076 4326 253078 4378
rect 253078 4326 253130 4378
rect 253130 4326 253132 4378
rect 253156 4326 253194 4378
rect 253194 4326 253206 4378
rect 253206 4326 253212 4378
rect 253236 4326 253258 4378
rect 253258 4326 253270 4378
rect 253270 4326 253292 4378
rect 253316 4326 253322 4378
rect 253322 4326 253334 4378
rect 253334 4326 253372 4378
rect 252836 4324 252892 4326
rect 252916 4324 252972 4326
rect 252996 4324 253052 4326
rect 253076 4324 253132 4326
rect 253156 4324 253212 4326
rect 253236 4324 253292 4326
rect 253316 4324 253372 4326
rect 252836 3290 252892 3292
rect 252916 3290 252972 3292
rect 252996 3290 253052 3292
rect 253076 3290 253132 3292
rect 253156 3290 253212 3292
rect 253236 3290 253292 3292
rect 253316 3290 253372 3292
rect 252836 3238 252874 3290
rect 252874 3238 252886 3290
rect 252886 3238 252892 3290
rect 252916 3238 252938 3290
rect 252938 3238 252950 3290
rect 252950 3238 252972 3290
rect 252996 3238 253002 3290
rect 253002 3238 253014 3290
rect 253014 3238 253052 3290
rect 253076 3238 253078 3290
rect 253078 3238 253130 3290
rect 253130 3238 253132 3290
rect 253156 3238 253194 3290
rect 253194 3238 253206 3290
rect 253206 3238 253212 3290
rect 253236 3238 253258 3290
rect 253258 3238 253270 3290
rect 253270 3238 253292 3290
rect 253316 3238 253322 3290
rect 253322 3238 253334 3290
rect 253334 3238 253372 3290
rect 252836 3236 252892 3238
rect 252916 3236 252972 3238
rect 252996 3236 253052 3238
rect 253076 3236 253132 3238
rect 253156 3236 253212 3238
rect 253236 3236 253292 3238
rect 253316 3236 253372 3238
rect 252836 2202 252892 2204
rect 252916 2202 252972 2204
rect 252996 2202 253052 2204
rect 253076 2202 253132 2204
rect 253156 2202 253212 2204
rect 253236 2202 253292 2204
rect 253316 2202 253372 2204
rect 252836 2150 252874 2202
rect 252874 2150 252886 2202
rect 252886 2150 252892 2202
rect 252916 2150 252938 2202
rect 252938 2150 252950 2202
rect 252950 2150 252972 2202
rect 252996 2150 253002 2202
rect 253002 2150 253014 2202
rect 253014 2150 253052 2202
rect 253076 2150 253078 2202
rect 253078 2150 253130 2202
rect 253130 2150 253132 2202
rect 253156 2150 253194 2202
rect 253194 2150 253206 2202
rect 253206 2150 253212 2202
rect 253236 2150 253258 2202
rect 253258 2150 253270 2202
rect 253270 2150 253292 2202
rect 253316 2150 253322 2202
rect 253322 2150 253334 2202
rect 253334 2150 253372 2202
rect 252836 2148 252892 2150
rect 252916 2148 252972 2150
rect 252996 2148 253052 2150
rect 253076 2148 253132 2150
rect 253156 2148 253212 2150
rect 253236 2148 253292 2150
rect 253316 2148 253372 2150
rect 270836 6010 270892 6012
rect 270916 6010 270972 6012
rect 270996 6010 271052 6012
rect 271076 6010 271132 6012
rect 271156 6010 271212 6012
rect 271236 6010 271292 6012
rect 271316 6010 271372 6012
rect 270836 5958 270874 6010
rect 270874 5958 270886 6010
rect 270886 5958 270892 6010
rect 270916 5958 270938 6010
rect 270938 5958 270950 6010
rect 270950 5958 270972 6010
rect 270996 5958 271002 6010
rect 271002 5958 271014 6010
rect 271014 5958 271052 6010
rect 271076 5958 271078 6010
rect 271078 5958 271130 6010
rect 271130 5958 271132 6010
rect 271156 5958 271194 6010
rect 271194 5958 271206 6010
rect 271206 5958 271212 6010
rect 271236 5958 271258 6010
rect 271258 5958 271270 6010
rect 271270 5958 271292 6010
rect 271316 5958 271322 6010
rect 271322 5958 271334 6010
rect 271334 5958 271372 6010
rect 270836 5956 270892 5958
rect 270916 5956 270972 5958
rect 270996 5956 271052 5958
rect 271076 5956 271132 5958
rect 271156 5956 271212 5958
rect 271236 5956 271292 5958
rect 271316 5956 271372 5958
rect 270836 4922 270892 4924
rect 270916 4922 270972 4924
rect 270996 4922 271052 4924
rect 271076 4922 271132 4924
rect 271156 4922 271212 4924
rect 271236 4922 271292 4924
rect 271316 4922 271372 4924
rect 270836 4870 270874 4922
rect 270874 4870 270886 4922
rect 270886 4870 270892 4922
rect 270916 4870 270938 4922
rect 270938 4870 270950 4922
rect 270950 4870 270972 4922
rect 270996 4870 271002 4922
rect 271002 4870 271014 4922
rect 271014 4870 271052 4922
rect 271076 4870 271078 4922
rect 271078 4870 271130 4922
rect 271130 4870 271132 4922
rect 271156 4870 271194 4922
rect 271194 4870 271206 4922
rect 271206 4870 271212 4922
rect 271236 4870 271258 4922
rect 271258 4870 271270 4922
rect 271270 4870 271292 4922
rect 271316 4870 271322 4922
rect 271322 4870 271334 4922
rect 271334 4870 271372 4922
rect 270836 4868 270892 4870
rect 270916 4868 270972 4870
rect 270996 4868 271052 4870
rect 271076 4868 271132 4870
rect 271156 4868 271212 4870
rect 271236 4868 271292 4870
rect 271316 4868 271372 4870
rect 270836 3834 270892 3836
rect 270916 3834 270972 3836
rect 270996 3834 271052 3836
rect 271076 3834 271132 3836
rect 271156 3834 271212 3836
rect 271236 3834 271292 3836
rect 271316 3834 271372 3836
rect 270836 3782 270874 3834
rect 270874 3782 270886 3834
rect 270886 3782 270892 3834
rect 270916 3782 270938 3834
rect 270938 3782 270950 3834
rect 270950 3782 270972 3834
rect 270996 3782 271002 3834
rect 271002 3782 271014 3834
rect 271014 3782 271052 3834
rect 271076 3782 271078 3834
rect 271078 3782 271130 3834
rect 271130 3782 271132 3834
rect 271156 3782 271194 3834
rect 271194 3782 271206 3834
rect 271206 3782 271212 3834
rect 271236 3782 271258 3834
rect 271258 3782 271270 3834
rect 271270 3782 271292 3834
rect 271316 3782 271322 3834
rect 271322 3782 271334 3834
rect 271334 3782 271372 3834
rect 270836 3780 270892 3782
rect 270916 3780 270972 3782
rect 270996 3780 271052 3782
rect 271076 3780 271132 3782
rect 271156 3780 271212 3782
rect 271236 3780 271292 3782
rect 271316 3780 271372 3782
rect 270836 2746 270892 2748
rect 270916 2746 270972 2748
rect 270996 2746 271052 2748
rect 271076 2746 271132 2748
rect 271156 2746 271212 2748
rect 271236 2746 271292 2748
rect 271316 2746 271372 2748
rect 270836 2694 270874 2746
rect 270874 2694 270886 2746
rect 270886 2694 270892 2746
rect 270916 2694 270938 2746
rect 270938 2694 270950 2746
rect 270950 2694 270972 2746
rect 270996 2694 271002 2746
rect 271002 2694 271014 2746
rect 271014 2694 271052 2746
rect 271076 2694 271078 2746
rect 271078 2694 271130 2746
rect 271130 2694 271132 2746
rect 271156 2694 271194 2746
rect 271194 2694 271206 2746
rect 271206 2694 271212 2746
rect 271236 2694 271258 2746
rect 271258 2694 271270 2746
rect 271270 2694 271292 2746
rect 271316 2694 271322 2746
rect 271322 2694 271334 2746
rect 271334 2694 271372 2746
rect 270836 2692 270892 2694
rect 270916 2692 270972 2694
rect 270996 2692 271052 2694
rect 271076 2692 271132 2694
rect 271156 2692 271212 2694
rect 271236 2692 271292 2694
rect 271316 2692 271372 2694
rect 288836 5466 288892 5468
rect 288916 5466 288972 5468
rect 288996 5466 289052 5468
rect 289076 5466 289132 5468
rect 289156 5466 289212 5468
rect 289236 5466 289292 5468
rect 289316 5466 289372 5468
rect 288836 5414 288874 5466
rect 288874 5414 288886 5466
rect 288886 5414 288892 5466
rect 288916 5414 288938 5466
rect 288938 5414 288950 5466
rect 288950 5414 288972 5466
rect 288996 5414 289002 5466
rect 289002 5414 289014 5466
rect 289014 5414 289052 5466
rect 289076 5414 289078 5466
rect 289078 5414 289130 5466
rect 289130 5414 289132 5466
rect 289156 5414 289194 5466
rect 289194 5414 289206 5466
rect 289206 5414 289212 5466
rect 289236 5414 289258 5466
rect 289258 5414 289270 5466
rect 289270 5414 289292 5466
rect 289316 5414 289322 5466
rect 289322 5414 289334 5466
rect 289334 5414 289372 5466
rect 288836 5412 288892 5414
rect 288916 5412 288972 5414
rect 288996 5412 289052 5414
rect 289076 5412 289132 5414
rect 289156 5412 289212 5414
rect 289236 5412 289292 5414
rect 289316 5412 289372 5414
rect 288836 4378 288892 4380
rect 288916 4378 288972 4380
rect 288996 4378 289052 4380
rect 289076 4378 289132 4380
rect 289156 4378 289212 4380
rect 289236 4378 289292 4380
rect 289316 4378 289372 4380
rect 288836 4326 288874 4378
rect 288874 4326 288886 4378
rect 288886 4326 288892 4378
rect 288916 4326 288938 4378
rect 288938 4326 288950 4378
rect 288950 4326 288972 4378
rect 288996 4326 289002 4378
rect 289002 4326 289014 4378
rect 289014 4326 289052 4378
rect 289076 4326 289078 4378
rect 289078 4326 289130 4378
rect 289130 4326 289132 4378
rect 289156 4326 289194 4378
rect 289194 4326 289206 4378
rect 289206 4326 289212 4378
rect 289236 4326 289258 4378
rect 289258 4326 289270 4378
rect 289270 4326 289292 4378
rect 289316 4326 289322 4378
rect 289322 4326 289334 4378
rect 289334 4326 289372 4378
rect 288836 4324 288892 4326
rect 288916 4324 288972 4326
rect 288996 4324 289052 4326
rect 289076 4324 289132 4326
rect 289156 4324 289212 4326
rect 289236 4324 289292 4326
rect 289316 4324 289372 4326
rect 288836 3290 288892 3292
rect 288916 3290 288972 3292
rect 288996 3290 289052 3292
rect 289076 3290 289132 3292
rect 289156 3290 289212 3292
rect 289236 3290 289292 3292
rect 289316 3290 289372 3292
rect 288836 3238 288874 3290
rect 288874 3238 288886 3290
rect 288886 3238 288892 3290
rect 288916 3238 288938 3290
rect 288938 3238 288950 3290
rect 288950 3238 288972 3290
rect 288996 3238 289002 3290
rect 289002 3238 289014 3290
rect 289014 3238 289052 3290
rect 289076 3238 289078 3290
rect 289078 3238 289130 3290
rect 289130 3238 289132 3290
rect 289156 3238 289194 3290
rect 289194 3238 289206 3290
rect 289206 3238 289212 3290
rect 289236 3238 289258 3290
rect 289258 3238 289270 3290
rect 289270 3238 289292 3290
rect 289316 3238 289322 3290
rect 289322 3238 289334 3290
rect 289334 3238 289372 3290
rect 288836 3236 288892 3238
rect 288916 3236 288972 3238
rect 288996 3236 289052 3238
rect 289076 3236 289132 3238
rect 289156 3236 289212 3238
rect 289236 3236 289292 3238
rect 289316 3236 289372 3238
rect 288836 2202 288892 2204
rect 288916 2202 288972 2204
rect 288996 2202 289052 2204
rect 289076 2202 289132 2204
rect 289156 2202 289212 2204
rect 289236 2202 289292 2204
rect 289316 2202 289372 2204
rect 288836 2150 288874 2202
rect 288874 2150 288886 2202
rect 288886 2150 288892 2202
rect 288916 2150 288938 2202
rect 288938 2150 288950 2202
rect 288950 2150 288972 2202
rect 288996 2150 289002 2202
rect 289002 2150 289014 2202
rect 289014 2150 289052 2202
rect 289076 2150 289078 2202
rect 289078 2150 289130 2202
rect 289130 2150 289132 2202
rect 289156 2150 289194 2202
rect 289194 2150 289206 2202
rect 289206 2150 289212 2202
rect 289236 2150 289258 2202
rect 289258 2150 289270 2202
rect 289270 2150 289292 2202
rect 289316 2150 289322 2202
rect 289322 2150 289334 2202
rect 289334 2150 289372 2202
rect 288836 2148 288892 2150
rect 288916 2148 288972 2150
rect 288996 2148 289052 2150
rect 289076 2148 289132 2150
rect 289156 2148 289212 2150
rect 289236 2148 289292 2150
rect 289316 2148 289372 2150
rect 306836 6010 306892 6012
rect 306916 6010 306972 6012
rect 306996 6010 307052 6012
rect 307076 6010 307132 6012
rect 307156 6010 307212 6012
rect 307236 6010 307292 6012
rect 307316 6010 307372 6012
rect 306836 5958 306874 6010
rect 306874 5958 306886 6010
rect 306886 5958 306892 6010
rect 306916 5958 306938 6010
rect 306938 5958 306950 6010
rect 306950 5958 306972 6010
rect 306996 5958 307002 6010
rect 307002 5958 307014 6010
rect 307014 5958 307052 6010
rect 307076 5958 307078 6010
rect 307078 5958 307130 6010
rect 307130 5958 307132 6010
rect 307156 5958 307194 6010
rect 307194 5958 307206 6010
rect 307206 5958 307212 6010
rect 307236 5958 307258 6010
rect 307258 5958 307270 6010
rect 307270 5958 307292 6010
rect 307316 5958 307322 6010
rect 307322 5958 307334 6010
rect 307334 5958 307372 6010
rect 306836 5956 306892 5958
rect 306916 5956 306972 5958
rect 306996 5956 307052 5958
rect 307076 5956 307132 5958
rect 307156 5956 307212 5958
rect 307236 5956 307292 5958
rect 307316 5956 307372 5958
rect 306836 4922 306892 4924
rect 306916 4922 306972 4924
rect 306996 4922 307052 4924
rect 307076 4922 307132 4924
rect 307156 4922 307212 4924
rect 307236 4922 307292 4924
rect 307316 4922 307372 4924
rect 306836 4870 306874 4922
rect 306874 4870 306886 4922
rect 306886 4870 306892 4922
rect 306916 4870 306938 4922
rect 306938 4870 306950 4922
rect 306950 4870 306972 4922
rect 306996 4870 307002 4922
rect 307002 4870 307014 4922
rect 307014 4870 307052 4922
rect 307076 4870 307078 4922
rect 307078 4870 307130 4922
rect 307130 4870 307132 4922
rect 307156 4870 307194 4922
rect 307194 4870 307206 4922
rect 307206 4870 307212 4922
rect 307236 4870 307258 4922
rect 307258 4870 307270 4922
rect 307270 4870 307292 4922
rect 307316 4870 307322 4922
rect 307322 4870 307334 4922
rect 307334 4870 307372 4922
rect 306836 4868 306892 4870
rect 306916 4868 306972 4870
rect 306996 4868 307052 4870
rect 307076 4868 307132 4870
rect 307156 4868 307212 4870
rect 307236 4868 307292 4870
rect 307316 4868 307372 4870
rect 306836 3834 306892 3836
rect 306916 3834 306972 3836
rect 306996 3834 307052 3836
rect 307076 3834 307132 3836
rect 307156 3834 307212 3836
rect 307236 3834 307292 3836
rect 307316 3834 307372 3836
rect 306836 3782 306874 3834
rect 306874 3782 306886 3834
rect 306886 3782 306892 3834
rect 306916 3782 306938 3834
rect 306938 3782 306950 3834
rect 306950 3782 306972 3834
rect 306996 3782 307002 3834
rect 307002 3782 307014 3834
rect 307014 3782 307052 3834
rect 307076 3782 307078 3834
rect 307078 3782 307130 3834
rect 307130 3782 307132 3834
rect 307156 3782 307194 3834
rect 307194 3782 307206 3834
rect 307206 3782 307212 3834
rect 307236 3782 307258 3834
rect 307258 3782 307270 3834
rect 307270 3782 307292 3834
rect 307316 3782 307322 3834
rect 307322 3782 307334 3834
rect 307334 3782 307372 3834
rect 306836 3780 306892 3782
rect 306916 3780 306972 3782
rect 306996 3780 307052 3782
rect 307076 3780 307132 3782
rect 307156 3780 307212 3782
rect 307236 3780 307292 3782
rect 307316 3780 307372 3782
rect 306836 2746 306892 2748
rect 306916 2746 306972 2748
rect 306996 2746 307052 2748
rect 307076 2746 307132 2748
rect 307156 2746 307212 2748
rect 307236 2746 307292 2748
rect 307316 2746 307372 2748
rect 306836 2694 306874 2746
rect 306874 2694 306886 2746
rect 306886 2694 306892 2746
rect 306916 2694 306938 2746
rect 306938 2694 306950 2746
rect 306950 2694 306972 2746
rect 306996 2694 307002 2746
rect 307002 2694 307014 2746
rect 307014 2694 307052 2746
rect 307076 2694 307078 2746
rect 307078 2694 307130 2746
rect 307130 2694 307132 2746
rect 307156 2694 307194 2746
rect 307194 2694 307206 2746
rect 307206 2694 307212 2746
rect 307236 2694 307258 2746
rect 307258 2694 307270 2746
rect 307270 2694 307292 2746
rect 307316 2694 307322 2746
rect 307322 2694 307334 2746
rect 307334 2694 307372 2746
rect 306836 2692 306892 2694
rect 306916 2692 306972 2694
rect 306996 2692 307052 2694
rect 307076 2692 307132 2694
rect 307156 2692 307212 2694
rect 307236 2692 307292 2694
rect 307316 2692 307372 2694
rect 324836 5466 324892 5468
rect 324916 5466 324972 5468
rect 324996 5466 325052 5468
rect 325076 5466 325132 5468
rect 325156 5466 325212 5468
rect 325236 5466 325292 5468
rect 325316 5466 325372 5468
rect 324836 5414 324874 5466
rect 324874 5414 324886 5466
rect 324886 5414 324892 5466
rect 324916 5414 324938 5466
rect 324938 5414 324950 5466
rect 324950 5414 324972 5466
rect 324996 5414 325002 5466
rect 325002 5414 325014 5466
rect 325014 5414 325052 5466
rect 325076 5414 325078 5466
rect 325078 5414 325130 5466
rect 325130 5414 325132 5466
rect 325156 5414 325194 5466
rect 325194 5414 325206 5466
rect 325206 5414 325212 5466
rect 325236 5414 325258 5466
rect 325258 5414 325270 5466
rect 325270 5414 325292 5466
rect 325316 5414 325322 5466
rect 325322 5414 325334 5466
rect 325334 5414 325372 5466
rect 324836 5412 324892 5414
rect 324916 5412 324972 5414
rect 324996 5412 325052 5414
rect 325076 5412 325132 5414
rect 325156 5412 325212 5414
rect 325236 5412 325292 5414
rect 325316 5412 325372 5414
rect 324836 4378 324892 4380
rect 324916 4378 324972 4380
rect 324996 4378 325052 4380
rect 325076 4378 325132 4380
rect 325156 4378 325212 4380
rect 325236 4378 325292 4380
rect 325316 4378 325372 4380
rect 324836 4326 324874 4378
rect 324874 4326 324886 4378
rect 324886 4326 324892 4378
rect 324916 4326 324938 4378
rect 324938 4326 324950 4378
rect 324950 4326 324972 4378
rect 324996 4326 325002 4378
rect 325002 4326 325014 4378
rect 325014 4326 325052 4378
rect 325076 4326 325078 4378
rect 325078 4326 325130 4378
rect 325130 4326 325132 4378
rect 325156 4326 325194 4378
rect 325194 4326 325206 4378
rect 325206 4326 325212 4378
rect 325236 4326 325258 4378
rect 325258 4326 325270 4378
rect 325270 4326 325292 4378
rect 325316 4326 325322 4378
rect 325322 4326 325334 4378
rect 325334 4326 325372 4378
rect 324836 4324 324892 4326
rect 324916 4324 324972 4326
rect 324996 4324 325052 4326
rect 325076 4324 325132 4326
rect 325156 4324 325212 4326
rect 325236 4324 325292 4326
rect 325316 4324 325372 4326
rect 324836 3290 324892 3292
rect 324916 3290 324972 3292
rect 324996 3290 325052 3292
rect 325076 3290 325132 3292
rect 325156 3290 325212 3292
rect 325236 3290 325292 3292
rect 325316 3290 325372 3292
rect 324836 3238 324874 3290
rect 324874 3238 324886 3290
rect 324886 3238 324892 3290
rect 324916 3238 324938 3290
rect 324938 3238 324950 3290
rect 324950 3238 324972 3290
rect 324996 3238 325002 3290
rect 325002 3238 325014 3290
rect 325014 3238 325052 3290
rect 325076 3238 325078 3290
rect 325078 3238 325130 3290
rect 325130 3238 325132 3290
rect 325156 3238 325194 3290
rect 325194 3238 325206 3290
rect 325206 3238 325212 3290
rect 325236 3238 325258 3290
rect 325258 3238 325270 3290
rect 325270 3238 325292 3290
rect 325316 3238 325322 3290
rect 325322 3238 325334 3290
rect 325334 3238 325372 3290
rect 324836 3236 324892 3238
rect 324916 3236 324972 3238
rect 324996 3236 325052 3238
rect 325076 3236 325132 3238
rect 325156 3236 325212 3238
rect 325236 3236 325292 3238
rect 325316 3236 325372 3238
rect 324836 2202 324892 2204
rect 324916 2202 324972 2204
rect 324996 2202 325052 2204
rect 325076 2202 325132 2204
rect 325156 2202 325212 2204
rect 325236 2202 325292 2204
rect 325316 2202 325372 2204
rect 324836 2150 324874 2202
rect 324874 2150 324886 2202
rect 324886 2150 324892 2202
rect 324916 2150 324938 2202
rect 324938 2150 324950 2202
rect 324950 2150 324972 2202
rect 324996 2150 325002 2202
rect 325002 2150 325014 2202
rect 325014 2150 325052 2202
rect 325076 2150 325078 2202
rect 325078 2150 325130 2202
rect 325130 2150 325132 2202
rect 325156 2150 325194 2202
rect 325194 2150 325206 2202
rect 325206 2150 325212 2202
rect 325236 2150 325258 2202
rect 325258 2150 325270 2202
rect 325270 2150 325292 2202
rect 325316 2150 325322 2202
rect 325322 2150 325334 2202
rect 325334 2150 325372 2202
rect 324836 2148 324892 2150
rect 324916 2148 324972 2150
rect 324996 2148 325052 2150
rect 325076 2148 325132 2150
rect 325156 2148 325212 2150
rect 325236 2148 325292 2150
rect 325316 2148 325372 2150
rect 342836 6010 342892 6012
rect 342916 6010 342972 6012
rect 342996 6010 343052 6012
rect 343076 6010 343132 6012
rect 343156 6010 343212 6012
rect 343236 6010 343292 6012
rect 343316 6010 343372 6012
rect 342836 5958 342874 6010
rect 342874 5958 342886 6010
rect 342886 5958 342892 6010
rect 342916 5958 342938 6010
rect 342938 5958 342950 6010
rect 342950 5958 342972 6010
rect 342996 5958 343002 6010
rect 343002 5958 343014 6010
rect 343014 5958 343052 6010
rect 343076 5958 343078 6010
rect 343078 5958 343130 6010
rect 343130 5958 343132 6010
rect 343156 5958 343194 6010
rect 343194 5958 343206 6010
rect 343206 5958 343212 6010
rect 343236 5958 343258 6010
rect 343258 5958 343270 6010
rect 343270 5958 343292 6010
rect 343316 5958 343322 6010
rect 343322 5958 343334 6010
rect 343334 5958 343372 6010
rect 342836 5956 342892 5958
rect 342916 5956 342972 5958
rect 342996 5956 343052 5958
rect 343076 5956 343132 5958
rect 343156 5956 343212 5958
rect 343236 5956 343292 5958
rect 343316 5956 343372 5958
rect 342836 4922 342892 4924
rect 342916 4922 342972 4924
rect 342996 4922 343052 4924
rect 343076 4922 343132 4924
rect 343156 4922 343212 4924
rect 343236 4922 343292 4924
rect 343316 4922 343372 4924
rect 342836 4870 342874 4922
rect 342874 4870 342886 4922
rect 342886 4870 342892 4922
rect 342916 4870 342938 4922
rect 342938 4870 342950 4922
rect 342950 4870 342972 4922
rect 342996 4870 343002 4922
rect 343002 4870 343014 4922
rect 343014 4870 343052 4922
rect 343076 4870 343078 4922
rect 343078 4870 343130 4922
rect 343130 4870 343132 4922
rect 343156 4870 343194 4922
rect 343194 4870 343206 4922
rect 343206 4870 343212 4922
rect 343236 4870 343258 4922
rect 343258 4870 343270 4922
rect 343270 4870 343292 4922
rect 343316 4870 343322 4922
rect 343322 4870 343334 4922
rect 343334 4870 343372 4922
rect 342836 4868 342892 4870
rect 342916 4868 342972 4870
rect 342996 4868 343052 4870
rect 343076 4868 343132 4870
rect 343156 4868 343212 4870
rect 343236 4868 343292 4870
rect 343316 4868 343372 4870
rect 342836 3834 342892 3836
rect 342916 3834 342972 3836
rect 342996 3834 343052 3836
rect 343076 3834 343132 3836
rect 343156 3834 343212 3836
rect 343236 3834 343292 3836
rect 343316 3834 343372 3836
rect 342836 3782 342874 3834
rect 342874 3782 342886 3834
rect 342886 3782 342892 3834
rect 342916 3782 342938 3834
rect 342938 3782 342950 3834
rect 342950 3782 342972 3834
rect 342996 3782 343002 3834
rect 343002 3782 343014 3834
rect 343014 3782 343052 3834
rect 343076 3782 343078 3834
rect 343078 3782 343130 3834
rect 343130 3782 343132 3834
rect 343156 3782 343194 3834
rect 343194 3782 343206 3834
rect 343206 3782 343212 3834
rect 343236 3782 343258 3834
rect 343258 3782 343270 3834
rect 343270 3782 343292 3834
rect 343316 3782 343322 3834
rect 343322 3782 343334 3834
rect 343334 3782 343372 3834
rect 342836 3780 342892 3782
rect 342916 3780 342972 3782
rect 342996 3780 343052 3782
rect 343076 3780 343132 3782
rect 343156 3780 343212 3782
rect 343236 3780 343292 3782
rect 343316 3780 343372 3782
rect 342836 2746 342892 2748
rect 342916 2746 342972 2748
rect 342996 2746 343052 2748
rect 343076 2746 343132 2748
rect 343156 2746 343212 2748
rect 343236 2746 343292 2748
rect 343316 2746 343372 2748
rect 342836 2694 342874 2746
rect 342874 2694 342886 2746
rect 342886 2694 342892 2746
rect 342916 2694 342938 2746
rect 342938 2694 342950 2746
rect 342950 2694 342972 2746
rect 342996 2694 343002 2746
rect 343002 2694 343014 2746
rect 343014 2694 343052 2746
rect 343076 2694 343078 2746
rect 343078 2694 343130 2746
rect 343130 2694 343132 2746
rect 343156 2694 343194 2746
rect 343194 2694 343206 2746
rect 343206 2694 343212 2746
rect 343236 2694 343258 2746
rect 343258 2694 343270 2746
rect 343270 2694 343292 2746
rect 343316 2694 343322 2746
rect 343322 2694 343334 2746
rect 343334 2694 343372 2746
rect 342836 2692 342892 2694
rect 342916 2692 342972 2694
rect 342996 2692 343052 2694
rect 343076 2692 343132 2694
rect 343156 2692 343212 2694
rect 343236 2692 343292 2694
rect 343316 2692 343372 2694
rect 360836 5466 360892 5468
rect 360916 5466 360972 5468
rect 360996 5466 361052 5468
rect 361076 5466 361132 5468
rect 361156 5466 361212 5468
rect 361236 5466 361292 5468
rect 361316 5466 361372 5468
rect 360836 5414 360874 5466
rect 360874 5414 360886 5466
rect 360886 5414 360892 5466
rect 360916 5414 360938 5466
rect 360938 5414 360950 5466
rect 360950 5414 360972 5466
rect 360996 5414 361002 5466
rect 361002 5414 361014 5466
rect 361014 5414 361052 5466
rect 361076 5414 361078 5466
rect 361078 5414 361130 5466
rect 361130 5414 361132 5466
rect 361156 5414 361194 5466
rect 361194 5414 361206 5466
rect 361206 5414 361212 5466
rect 361236 5414 361258 5466
rect 361258 5414 361270 5466
rect 361270 5414 361292 5466
rect 361316 5414 361322 5466
rect 361322 5414 361334 5466
rect 361334 5414 361372 5466
rect 360836 5412 360892 5414
rect 360916 5412 360972 5414
rect 360996 5412 361052 5414
rect 361076 5412 361132 5414
rect 361156 5412 361212 5414
rect 361236 5412 361292 5414
rect 361316 5412 361372 5414
rect 360836 4378 360892 4380
rect 360916 4378 360972 4380
rect 360996 4378 361052 4380
rect 361076 4378 361132 4380
rect 361156 4378 361212 4380
rect 361236 4378 361292 4380
rect 361316 4378 361372 4380
rect 360836 4326 360874 4378
rect 360874 4326 360886 4378
rect 360886 4326 360892 4378
rect 360916 4326 360938 4378
rect 360938 4326 360950 4378
rect 360950 4326 360972 4378
rect 360996 4326 361002 4378
rect 361002 4326 361014 4378
rect 361014 4326 361052 4378
rect 361076 4326 361078 4378
rect 361078 4326 361130 4378
rect 361130 4326 361132 4378
rect 361156 4326 361194 4378
rect 361194 4326 361206 4378
rect 361206 4326 361212 4378
rect 361236 4326 361258 4378
rect 361258 4326 361270 4378
rect 361270 4326 361292 4378
rect 361316 4326 361322 4378
rect 361322 4326 361334 4378
rect 361334 4326 361372 4378
rect 360836 4324 360892 4326
rect 360916 4324 360972 4326
rect 360996 4324 361052 4326
rect 361076 4324 361132 4326
rect 361156 4324 361212 4326
rect 361236 4324 361292 4326
rect 361316 4324 361372 4326
rect 360836 3290 360892 3292
rect 360916 3290 360972 3292
rect 360996 3290 361052 3292
rect 361076 3290 361132 3292
rect 361156 3290 361212 3292
rect 361236 3290 361292 3292
rect 361316 3290 361372 3292
rect 360836 3238 360874 3290
rect 360874 3238 360886 3290
rect 360886 3238 360892 3290
rect 360916 3238 360938 3290
rect 360938 3238 360950 3290
rect 360950 3238 360972 3290
rect 360996 3238 361002 3290
rect 361002 3238 361014 3290
rect 361014 3238 361052 3290
rect 361076 3238 361078 3290
rect 361078 3238 361130 3290
rect 361130 3238 361132 3290
rect 361156 3238 361194 3290
rect 361194 3238 361206 3290
rect 361206 3238 361212 3290
rect 361236 3238 361258 3290
rect 361258 3238 361270 3290
rect 361270 3238 361292 3290
rect 361316 3238 361322 3290
rect 361322 3238 361334 3290
rect 361334 3238 361372 3290
rect 360836 3236 360892 3238
rect 360916 3236 360972 3238
rect 360996 3236 361052 3238
rect 361076 3236 361132 3238
rect 361156 3236 361212 3238
rect 361236 3236 361292 3238
rect 361316 3236 361372 3238
rect 360836 2202 360892 2204
rect 360916 2202 360972 2204
rect 360996 2202 361052 2204
rect 361076 2202 361132 2204
rect 361156 2202 361212 2204
rect 361236 2202 361292 2204
rect 361316 2202 361372 2204
rect 360836 2150 360874 2202
rect 360874 2150 360886 2202
rect 360886 2150 360892 2202
rect 360916 2150 360938 2202
rect 360938 2150 360950 2202
rect 360950 2150 360972 2202
rect 360996 2150 361002 2202
rect 361002 2150 361014 2202
rect 361014 2150 361052 2202
rect 361076 2150 361078 2202
rect 361078 2150 361130 2202
rect 361130 2150 361132 2202
rect 361156 2150 361194 2202
rect 361194 2150 361206 2202
rect 361206 2150 361212 2202
rect 361236 2150 361258 2202
rect 361258 2150 361270 2202
rect 361270 2150 361292 2202
rect 361316 2150 361322 2202
rect 361322 2150 361334 2202
rect 361334 2150 361372 2202
rect 360836 2148 360892 2150
rect 360916 2148 360972 2150
rect 360996 2148 361052 2150
rect 361076 2148 361132 2150
rect 361156 2148 361212 2150
rect 361236 2148 361292 2150
rect 361316 2148 361372 2150
rect 378836 6010 378892 6012
rect 378916 6010 378972 6012
rect 378996 6010 379052 6012
rect 379076 6010 379132 6012
rect 379156 6010 379212 6012
rect 379236 6010 379292 6012
rect 379316 6010 379372 6012
rect 378836 5958 378874 6010
rect 378874 5958 378886 6010
rect 378886 5958 378892 6010
rect 378916 5958 378938 6010
rect 378938 5958 378950 6010
rect 378950 5958 378972 6010
rect 378996 5958 379002 6010
rect 379002 5958 379014 6010
rect 379014 5958 379052 6010
rect 379076 5958 379078 6010
rect 379078 5958 379130 6010
rect 379130 5958 379132 6010
rect 379156 5958 379194 6010
rect 379194 5958 379206 6010
rect 379206 5958 379212 6010
rect 379236 5958 379258 6010
rect 379258 5958 379270 6010
rect 379270 5958 379292 6010
rect 379316 5958 379322 6010
rect 379322 5958 379334 6010
rect 379334 5958 379372 6010
rect 378836 5956 378892 5958
rect 378916 5956 378972 5958
rect 378996 5956 379052 5958
rect 379076 5956 379132 5958
rect 379156 5956 379212 5958
rect 379236 5956 379292 5958
rect 379316 5956 379372 5958
rect 378836 4922 378892 4924
rect 378916 4922 378972 4924
rect 378996 4922 379052 4924
rect 379076 4922 379132 4924
rect 379156 4922 379212 4924
rect 379236 4922 379292 4924
rect 379316 4922 379372 4924
rect 378836 4870 378874 4922
rect 378874 4870 378886 4922
rect 378886 4870 378892 4922
rect 378916 4870 378938 4922
rect 378938 4870 378950 4922
rect 378950 4870 378972 4922
rect 378996 4870 379002 4922
rect 379002 4870 379014 4922
rect 379014 4870 379052 4922
rect 379076 4870 379078 4922
rect 379078 4870 379130 4922
rect 379130 4870 379132 4922
rect 379156 4870 379194 4922
rect 379194 4870 379206 4922
rect 379206 4870 379212 4922
rect 379236 4870 379258 4922
rect 379258 4870 379270 4922
rect 379270 4870 379292 4922
rect 379316 4870 379322 4922
rect 379322 4870 379334 4922
rect 379334 4870 379372 4922
rect 378836 4868 378892 4870
rect 378916 4868 378972 4870
rect 378996 4868 379052 4870
rect 379076 4868 379132 4870
rect 379156 4868 379212 4870
rect 379236 4868 379292 4870
rect 379316 4868 379372 4870
rect 378836 3834 378892 3836
rect 378916 3834 378972 3836
rect 378996 3834 379052 3836
rect 379076 3834 379132 3836
rect 379156 3834 379212 3836
rect 379236 3834 379292 3836
rect 379316 3834 379372 3836
rect 378836 3782 378874 3834
rect 378874 3782 378886 3834
rect 378886 3782 378892 3834
rect 378916 3782 378938 3834
rect 378938 3782 378950 3834
rect 378950 3782 378972 3834
rect 378996 3782 379002 3834
rect 379002 3782 379014 3834
rect 379014 3782 379052 3834
rect 379076 3782 379078 3834
rect 379078 3782 379130 3834
rect 379130 3782 379132 3834
rect 379156 3782 379194 3834
rect 379194 3782 379206 3834
rect 379206 3782 379212 3834
rect 379236 3782 379258 3834
rect 379258 3782 379270 3834
rect 379270 3782 379292 3834
rect 379316 3782 379322 3834
rect 379322 3782 379334 3834
rect 379334 3782 379372 3834
rect 378836 3780 378892 3782
rect 378916 3780 378972 3782
rect 378996 3780 379052 3782
rect 379076 3780 379132 3782
rect 379156 3780 379212 3782
rect 379236 3780 379292 3782
rect 379316 3780 379372 3782
rect 378836 2746 378892 2748
rect 378916 2746 378972 2748
rect 378996 2746 379052 2748
rect 379076 2746 379132 2748
rect 379156 2746 379212 2748
rect 379236 2746 379292 2748
rect 379316 2746 379372 2748
rect 378836 2694 378874 2746
rect 378874 2694 378886 2746
rect 378886 2694 378892 2746
rect 378916 2694 378938 2746
rect 378938 2694 378950 2746
rect 378950 2694 378972 2746
rect 378996 2694 379002 2746
rect 379002 2694 379014 2746
rect 379014 2694 379052 2746
rect 379076 2694 379078 2746
rect 379078 2694 379130 2746
rect 379130 2694 379132 2746
rect 379156 2694 379194 2746
rect 379194 2694 379206 2746
rect 379206 2694 379212 2746
rect 379236 2694 379258 2746
rect 379258 2694 379270 2746
rect 379270 2694 379292 2746
rect 379316 2694 379322 2746
rect 379322 2694 379334 2746
rect 379334 2694 379372 2746
rect 378836 2692 378892 2694
rect 378916 2692 378972 2694
rect 378996 2692 379052 2694
rect 379076 2692 379132 2694
rect 379156 2692 379212 2694
rect 379236 2692 379292 2694
rect 379316 2692 379372 2694
rect 396836 5466 396892 5468
rect 396916 5466 396972 5468
rect 396996 5466 397052 5468
rect 397076 5466 397132 5468
rect 397156 5466 397212 5468
rect 397236 5466 397292 5468
rect 397316 5466 397372 5468
rect 396836 5414 396874 5466
rect 396874 5414 396886 5466
rect 396886 5414 396892 5466
rect 396916 5414 396938 5466
rect 396938 5414 396950 5466
rect 396950 5414 396972 5466
rect 396996 5414 397002 5466
rect 397002 5414 397014 5466
rect 397014 5414 397052 5466
rect 397076 5414 397078 5466
rect 397078 5414 397130 5466
rect 397130 5414 397132 5466
rect 397156 5414 397194 5466
rect 397194 5414 397206 5466
rect 397206 5414 397212 5466
rect 397236 5414 397258 5466
rect 397258 5414 397270 5466
rect 397270 5414 397292 5466
rect 397316 5414 397322 5466
rect 397322 5414 397334 5466
rect 397334 5414 397372 5466
rect 396836 5412 396892 5414
rect 396916 5412 396972 5414
rect 396996 5412 397052 5414
rect 397076 5412 397132 5414
rect 397156 5412 397212 5414
rect 397236 5412 397292 5414
rect 397316 5412 397372 5414
rect 396836 4378 396892 4380
rect 396916 4378 396972 4380
rect 396996 4378 397052 4380
rect 397076 4378 397132 4380
rect 397156 4378 397212 4380
rect 397236 4378 397292 4380
rect 397316 4378 397372 4380
rect 396836 4326 396874 4378
rect 396874 4326 396886 4378
rect 396886 4326 396892 4378
rect 396916 4326 396938 4378
rect 396938 4326 396950 4378
rect 396950 4326 396972 4378
rect 396996 4326 397002 4378
rect 397002 4326 397014 4378
rect 397014 4326 397052 4378
rect 397076 4326 397078 4378
rect 397078 4326 397130 4378
rect 397130 4326 397132 4378
rect 397156 4326 397194 4378
rect 397194 4326 397206 4378
rect 397206 4326 397212 4378
rect 397236 4326 397258 4378
rect 397258 4326 397270 4378
rect 397270 4326 397292 4378
rect 397316 4326 397322 4378
rect 397322 4326 397334 4378
rect 397334 4326 397372 4378
rect 396836 4324 396892 4326
rect 396916 4324 396972 4326
rect 396996 4324 397052 4326
rect 397076 4324 397132 4326
rect 397156 4324 397212 4326
rect 397236 4324 397292 4326
rect 397316 4324 397372 4326
rect 396836 3290 396892 3292
rect 396916 3290 396972 3292
rect 396996 3290 397052 3292
rect 397076 3290 397132 3292
rect 397156 3290 397212 3292
rect 397236 3290 397292 3292
rect 397316 3290 397372 3292
rect 396836 3238 396874 3290
rect 396874 3238 396886 3290
rect 396886 3238 396892 3290
rect 396916 3238 396938 3290
rect 396938 3238 396950 3290
rect 396950 3238 396972 3290
rect 396996 3238 397002 3290
rect 397002 3238 397014 3290
rect 397014 3238 397052 3290
rect 397076 3238 397078 3290
rect 397078 3238 397130 3290
rect 397130 3238 397132 3290
rect 397156 3238 397194 3290
rect 397194 3238 397206 3290
rect 397206 3238 397212 3290
rect 397236 3238 397258 3290
rect 397258 3238 397270 3290
rect 397270 3238 397292 3290
rect 397316 3238 397322 3290
rect 397322 3238 397334 3290
rect 397334 3238 397372 3290
rect 396836 3236 396892 3238
rect 396916 3236 396972 3238
rect 396996 3236 397052 3238
rect 397076 3236 397132 3238
rect 397156 3236 397212 3238
rect 397236 3236 397292 3238
rect 397316 3236 397372 3238
rect 396836 2202 396892 2204
rect 396916 2202 396972 2204
rect 396996 2202 397052 2204
rect 397076 2202 397132 2204
rect 397156 2202 397212 2204
rect 397236 2202 397292 2204
rect 397316 2202 397372 2204
rect 396836 2150 396874 2202
rect 396874 2150 396886 2202
rect 396886 2150 396892 2202
rect 396916 2150 396938 2202
rect 396938 2150 396950 2202
rect 396950 2150 396972 2202
rect 396996 2150 397002 2202
rect 397002 2150 397014 2202
rect 397014 2150 397052 2202
rect 397076 2150 397078 2202
rect 397078 2150 397130 2202
rect 397130 2150 397132 2202
rect 397156 2150 397194 2202
rect 397194 2150 397206 2202
rect 397206 2150 397212 2202
rect 397236 2150 397258 2202
rect 397258 2150 397270 2202
rect 397270 2150 397292 2202
rect 397316 2150 397322 2202
rect 397322 2150 397334 2202
rect 397334 2150 397372 2202
rect 396836 2148 396892 2150
rect 396916 2148 396972 2150
rect 396996 2148 397052 2150
rect 397076 2148 397132 2150
rect 397156 2148 397212 2150
rect 397236 2148 397292 2150
rect 397316 2148 397372 2150
rect 414836 6010 414892 6012
rect 414916 6010 414972 6012
rect 414996 6010 415052 6012
rect 415076 6010 415132 6012
rect 415156 6010 415212 6012
rect 415236 6010 415292 6012
rect 415316 6010 415372 6012
rect 414836 5958 414874 6010
rect 414874 5958 414886 6010
rect 414886 5958 414892 6010
rect 414916 5958 414938 6010
rect 414938 5958 414950 6010
rect 414950 5958 414972 6010
rect 414996 5958 415002 6010
rect 415002 5958 415014 6010
rect 415014 5958 415052 6010
rect 415076 5958 415078 6010
rect 415078 5958 415130 6010
rect 415130 5958 415132 6010
rect 415156 5958 415194 6010
rect 415194 5958 415206 6010
rect 415206 5958 415212 6010
rect 415236 5958 415258 6010
rect 415258 5958 415270 6010
rect 415270 5958 415292 6010
rect 415316 5958 415322 6010
rect 415322 5958 415334 6010
rect 415334 5958 415372 6010
rect 414836 5956 414892 5958
rect 414916 5956 414972 5958
rect 414996 5956 415052 5958
rect 415076 5956 415132 5958
rect 415156 5956 415212 5958
rect 415236 5956 415292 5958
rect 415316 5956 415372 5958
rect 414836 4922 414892 4924
rect 414916 4922 414972 4924
rect 414996 4922 415052 4924
rect 415076 4922 415132 4924
rect 415156 4922 415212 4924
rect 415236 4922 415292 4924
rect 415316 4922 415372 4924
rect 414836 4870 414874 4922
rect 414874 4870 414886 4922
rect 414886 4870 414892 4922
rect 414916 4870 414938 4922
rect 414938 4870 414950 4922
rect 414950 4870 414972 4922
rect 414996 4870 415002 4922
rect 415002 4870 415014 4922
rect 415014 4870 415052 4922
rect 415076 4870 415078 4922
rect 415078 4870 415130 4922
rect 415130 4870 415132 4922
rect 415156 4870 415194 4922
rect 415194 4870 415206 4922
rect 415206 4870 415212 4922
rect 415236 4870 415258 4922
rect 415258 4870 415270 4922
rect 415270 4870 415292 4922
rect 415316 4870 415322 4922
rect 415322 4870 415334 4922
rect 415334 4870 415372 4922
rect 414836 4868 414892 4870
rect 414916 4868 414972 4870
rect 414996 4868 415052 4870
rect 415076 4868 415132 4870
rect 415156 4868 415212 4870
rect 415236 4868 415292 4870
rect 415316 4868 415372 4870
rect 414836 3834 414892 3836
rect 414916 3834 414972 3836
rect 414996 3834 415052 3836
rect 415076 3834 415132 3836
rect 415156 3834 415212 3836
rect 415236 3834 415292 3836
rect 415316 3834 415372 3836
rect 414836 3782 414874 3834
rect 414874 3782 414886 3834
rect 414886 3782 414892 3834
rect 414916 3782 414938 3834
rect 414938 3782 414950 3834
rect 414950 3782 414972 3834
rect 414996 3782 415002 3834
rect 415002 3782 415014 3834
rect 415014 3782 415052 3834
rect 415076 3782 415078 3834
rect 415078 3782 415130 3834
rect 415130 3782 415132 3834
rect 415156 3782 415194 3834
rect 415194 3782 415206 3834
rect 415206 3782 415212 3834
rect 415236 3782 415258 3834
rect 415258 3782 415270 3834
rect 415270 3782 415292 3834
rect 415316 3782 415322 3834
rect 415322 3782 415334 3834
rect 415334 3782 415372 3834
rect 414836 3780 414892 3782
rect 414916 3780 414972 3782
rect 414996 3780 415052 3782
rect 415076 3780 415132 3782
rect 415156 3780 415212 3782
rect 415236 3780 415292 3782
rect 415316 3780 415372 3782
rect 414836 2746 414892 2748
rect 414916 2746 414972 2748
rect 414996 2746 415052 2748
rect 415076 2746 415132 2748
rect 415156 2746 415212 2748
rect 415236 2746 415292 2748
rect 415316 2746 415372 2748
rect 414836 2694 414874 2746
rect 414874 2694 414886 2746
rect 414886 2694 414892 2746
rect 414916 2694 414938 2746
rect 414938 2694 414950 2746
rect 414950 2694 414972 2746
rect 414996 2694 415002 2746
rect 415002 2694 415014 2746
rect 415014 2694 415052 2746
rect 415076 2694 415078 2746
rect 415078 2694 415130 2746
rect 415130 2694 415132 2746
rect 415156 2694 415194 2746
rect 415194 2694 415206 2746
rect 415206 2694 415212 2746
rect 415236 2694 415258 2746
rect 415258 2694 415270 2746
rect 415270 2694 415292 2746
rect 415316 2694 415322 2746
rect 415322 2694 415334 2746
rect 415334 2694 415372 2746
rect 414836 2692 414892 2694
rect 414916 2692 414972 2694
rect 414996 2692 415052 2694
rect 415076 2692 415132 2694
rect 415156 2692 415212 2694
rect 415236 2692 415292 2694
rect 415316 2692 415372 2694
rect 432836 5466 432892 5468
rect 432916 5466 432972 5468
rect 432996 5466 433052 5468
rect 433076 5466 433132 5468
rect 433156 5466 433212 5468
rect 433236 5466 433292 5468
rect 433316 5466 433372 5468
rect 432836 5414 432874 5466
rect 432874 5414 432886 5466
rect 432886 5414 432892 5466
rect 432916 5414 432938 5466
rect 432938 5414 432950 5466
rect 432950 5414 432972 5466
rect 432996 5414 433002 5466
rect 433002 5414 433014 5466
rect 433014 5414 433052 5466
rect 433076 5414 433078 5466
rect 433078 5414 433130 5466
rect 433130 5414 433132 5466
rect 433156 5414 433194 5466
rect 433194 5414 433206 5466
rect 433206 5414 433212 5466
rect 433236 5414 433258 5466
rect 433258 5414 433270 5466
rect 433270 5414 433292 5466
rect 433316 5414 433322 5466
rect 433322 5414 433334 5466
rect 433334 5414 433372 5466
rect 432836 5412 432892 5414
rect 432916 5412 432972 5414
rect 432996 5412 433052 5414
rect 433076 5412 433132 5414
rect 433156 5412 433212 5414
rect 433236 5412 433292 5414
rect 433316 5412 433372 5414
rect 432836 4378 432892 4380
rect 432916 4378 432972 4380
rect 432996 4378 433052 4380
rect 433076 4378 433132 4380
rect 433156 4378 433212 4380
rect 433236 4378 433292 4380
rect 433316 4378 433372 4380
rect 432836 4326 432874 4378
rect 432874 4326 432886 4378
rect 432886 4326 432892 4378
rect 432916 4326 432938 4378
rect 432938 4326 432950 4378
rect 432950 4326 432972 4378
rect 432996 4326 433002 4378
rect 433002 4326 433014 4378
rect 433014 4326 433052 4378
rect 433076 4326 433078 4378
rect 433078 4326 433130 4378
rect 433130 4326 433132 4378
rect 433156 4326 433194 4378
rect 433194 4326 433206 4378
rect 433206 4326 433212 4378
rect 433236 4326 433258 4378
rect 433258 4326 433270 4378
rect 433270 4326 433292 4378
rect 433316 4326 433322 4378
rect 433322 4326 433334 4378
rect 433334 4326 433372 4378
rect 432836 4324 432892 4326
rect 432916 4324 432972 4326
rect 432996 4324 433052 4326
rect 433076 4324 433132 4326
rect 433156 4324 433212 4326
rect 433236 4324 433292 4326
rect 433316 4324 433372 4326
rect 432836 3290 432892 3292
rect 432916 3290 432972 3292
rect 432996 3290 433052 3292
rect 433076 3290 433132 3292
rect 433156 3290 433212 3292
rect 433236 3290 433292 3292
rect 433316 3290 433372 3292
rect 432836 3238 432874 3290
rect 432874 3238 432886 3290
rect 432886 3238 432892 3290
rect 432916 3238 432938 3290
rect 432938 3238 432950 3290
rect 432950 3238 432972 3290
rect 432996 3238 433002 3290
rect 433002 3238 433014 3290
rect 433014 3238 433052 3290
rect 433076 3238 433078 3290
rect 433078 3238 433130 3290
rect 433130 3238 433132 3290
rect 433156 3238 433194 3290
rect 433194 3238 433206 3290
rect 433206 3238 433212 3290
rect 433236 3238 433258 3290
rect 433258 3238 433270 3290
rect 433270 3238 433292 3290
rect 433316 3238 433322 3290
rect 433322 3238 433334 3290
rect 433334 3238 433372 3290
rect 432836 3236 432892 3238
rect 432916 3236 432972 3238
rect 432996 3236 433052 3238
rect 433076 3236 433132 3238
rect 433156 3236 433212 3238
rect 433236 3236 433292 3238
rect 433316 3236 433372 3238
rect 432836 2202 432892 2204
rect 432916 2202 432972 2204
rect 432996 2202 433052 2204
rect 433076 2202 433132 2204
rect 433156 2202 433212 2204
rect 433236 2202 433292 2204
rect 433316 2202 433372 2204
rect 432836 2150 432874 2202
rect 432874 2150 432886 2202
rect 432886 2150 432892 2202
rect 432916 2150 432938 2202
rect 432938 2150 432950 2202
rect 432950 2150 432972 2202
rect 432996 2150 433002 2202
rect 433002 2150 433014 2202
rect 433014 2150 433052 2202
rect 433076 2150 433078 2202
rect 433078 2150 433130 2202
rect 433130 2150 433132 2202
rect 433156 2150 433194 2202
rect 433194 2150 433206 2202
rect 433206 2150 433212 2202
rect 433236 2150 433258 2202
rect 433258 2150 433270 2202
rect 433270 2150 433292 2202
rect 433316 2150 433322 2202
rect 433322 2150 433334 2202
rect 433334 2150 433372 2202
rect 432836 2148 432892 2150
rect 432916 2148 432972 2150
rect 432996 2148 433052 2150
rect 433076 2148 433132 2150
rect 433156 2148 433212 2150
rect 433236 2148 433292 2150
rect 433316 2148 433372 2150
rect 450836 6010 450892 6012
rect 450916 6010 450972 6012
rect 450996 6010 451052 6012
rect 451076 6010 451132 6012
rect 451156 6010 451212 6012
rect 451236 6010 451292 6012
rect 451316 6010 451372 6012
rect 450836 5958 450874 6010
rect 450874 5958 450886 6010
rect 450886 5958 450892 6010
rect 450916 5958 450938 6010
rect 450938 5958 450950 6010
rect 450950 5958 450972 6010
rect 450996 5958 451002 6010
rect 451002 5958 451014 6010
rect 451014 5958 451052 6010
rect 451076 5958 451078 6010
rect 451078 5958 451130 6010
rect 451130 5958 451132 6010
rect 451156 5958 451194 6010
rect 451194 5958 451206 6010
rect 451206 5958 451212 6010
rect 451236 5958 451258 6010
rect 451258 5958 451270 6010
rect 451270 5958 451292 6010
rect 451316 5958 451322 6010
rect 451322 5958 451334 6010
rect 451334 5958 451372 6010
rect 450836 5956 450892 5958
rect 450916 5956 450972 5958
rect 450996 5956 451052 5958
rect 451076 5956 451132 5958
rect 451156 5956 451212 5958
rect 451236 5956 451292 5958
rect 451316 5956 451372 5958
rect 450836 4922 450892 4924
rect 450916 4922 450972 4924
rect 450996 4922 451052 4924
rect 451076 4922 451132 4924
rect 451156 4922 451212 4924
rect 451236 4922 451292 4924
rect 451316 4922 451372 4924
rect 450836 4870 450874 4922
rect 450874 4870 450886 4922
rect 450886 4870 450892 4922
rect 450916 4870 450938 4922
rect 450938 4870 450950 4922
rect 450950 4870 450972 4922
rect 450996 4870 451002 4922
rect 451002 4870 451014 4922
rect 451014 4870 451052 4922
rect 451076 4870 451078 4922
rect 451078 4870 451130 4922
rect 451130 4870 451132 4922
rect 451156 4870 451194 4922
rect 451194 4870 451206 4922
rect 451206 4870 451212 4922
rect 451236 4870 451258 4922
rect 451258 4870 451270 4922
rect 451270 4870 451292 4922
rect 451316 4870 451322 4922
rect 451322 4870 451334 4922
rect 451334 4870 451372 4922
rect 450836 4868 450892 4870
rect 450916 4868 450972 4870
rect 450996 4868 451052 4870
rect 451076 4868 451132 4870
rect 451156 4868 451212 4870
rect 451236 4868 451292 4870
rect 451316 4868 451372 4870
rect 450836 3834 450892 3836
rect 450916 3834 450972 3836
rect 450996 3834 451052 3836
rect 451076 3834 451132 3836
rect 451156 3834 451212 3836
rect 451236 3834 451292 3836
rect 451316 3834 451372 3836
rect 450836 3782 450874 3834
rect 450874 3782 450886 3834
rect 450886 3782 450892 3834
rect 450916 3782 450938 3834
rect 450938 3782 450950 3834
rect 450950 3782 450972 3834
rect 450996 3782 451002 3834
rect 451002 3782 451014 3834
rect 451014 3782 451052 3834
rect 451076 3782 451078 3834
rect 451078 3782 451130 3834
rect 451130 3782 451132 3834
rect 451156 3782 451194 3834
rect 451194 3782 451206 3834
rect 451206 3782 451212 3834
rect 451236 3782 451258 3834
rect 451258 3782 451270 3834
rect 451270 3782 451292 3834
rect 451316 3782 451322 3834
rect 451322 3782 451334 3834
rect 451334 3782 451372 3834
rect 450836 3780 450892 3782
rect 450916 3780 450972 3782
rect 450996 3780 451052 3782
rect 451076 3780 451132 3782
rect 451156 3780 451212 3782
rect 451236 3780 451292 3782
rect 451316 3780 451372 3782
rect 450836 2746 450892 2748
rect 450916 2746 450972 2748
rect 450996 2746 451052 2748
rect 451076 2746 451132 2748
rect 451156 2746 451212 2748
rect 451236 2746 451292 2748
rect 451316 2746 451372 2748
rect 450836 2694 450874 2746
rect 450874 2694 450886 2746
rect 450886 2694 450892 2746
rect 450916 2694 450938 2746
rect 450938 2694 450950 2746
rect 450950 2694 450972 2746
rect 450996 2694 451002 2746
rect 451002 2694 451014 2746
rect 451014 2694 451052 2746
rect 451076 2694 451078 2746
rect 451078 2694 451130 2746
rect 451130 2694 451132 2746
rect 451156 2694 451194 2746
rect 451194 2694 451206 2746
rect 451206 2694 451212 2746
rect 451236 2694 451258 2746
rect 451258 2694 451270 2746
rect 451270 2694 451292 2746
rect 451316 2694 451322 2746
rect 451322 2694 451334 2746
rect 451334 2694 451372 2746
rect 450836 2692 450892 2694
rect 450916 2692 450972 2694
rect 450996 2692 451052 2694
rect 451076 2692 451132 2694
rect 451156 2692 451212 2694
rect 451236 2692 451292 2694
rect 451316 2692 451372 2694
rect 468836 5466 468892 5468
rect 468916 5466 468972 5468
rect 468996 5466 469052 5468
rect 469076 5466 469132 5468
rect 469156 5466 469212 5468
rect 469236 5466 469292 5468
rect 469316 5466 469372 5468
rect 468836 5414 468874 5466
rect 468874 5414 468886 5466
rect 468886 5414 468892 5466
rect 468916 5414 468938 5466
rect 468938 5414 468950 5466
rect 468950 5414 468972 5466
rect 468996 5414 469002 5466
rect 469002 5414 469014 5466
rect 469014 5414 469052 5466
rect 469076 5414 469078 5466
rect 469078 5414 469130 5466
rect 469130 5414 469132 5466
rect 469156 5414 469194 5466
rect 469194 5414 469206 5466
rect 469206 5414 469212 5466
rect 469236 5414 469258 5466
rect 469258 5414 469270 5466
rect 469270 5414 469292 5466
rect 469316 5414 469322 5466
rect 469322 5414 469334 5466
rect 469334 5414 469372 5466
rect 468836 5412 468892 5414
rect 468916 5412 468972 5414
rect 468996 5412 469052 5414
rect 469076 5412 469132 5414
rect 469156 5412 469212 5414
rect 469236 5412 469292 5414
rect 469316 5412 469372 5414
rect 468836 4378 468892 4380
rect 468916 4378 468972 4380
rect 468996 4378 469052 4380
rect 469076 4378 469132 4380
rect 469156 4378 469212 4380
rect 469236 4378 469292 4380
rect 469316 4378 469372 4380
rect 468836 4326 468874 4378
rect 468874 4326 468886 4378
rect 468886 4326 468892 4378
rect 468916 4326 468938 4378
rect 468938 4326 468950 4378
rect 468950 4326 468972 4378
rect 468996 4326 469002 4378
rect 469002 4326 469014 4378
rect 469014 4326 469052 4378
rect 469076 4326 469078 4378
rect 469078 4326 469130 4378
rect 469130 4326 469132 4378
rect 469156 4326 469194 4378
rect 469194 4326 469206 4378
rect 469206 4326 469212 4378
rect 469236 4326 469258 4378
rect 469258 4326 469270 4378
rect 469270 4326 469292 4378
rect 469316 4326 469322 4378
rect 469322 4326 469334 4378
rect 469334 4326 469372 4378
rect 468836 4324 468892 4326
rect 468916 4324 468972 4326
rect 468996 4324 469052 4326
rect 469076 4324 469132 4326
rect 469156 4324 469212 4326
rect 469236 4324 469292 4326
rect 469316 4324 469372 4326
rect 468836 3290 468892 3292
rect 468916 3290 468972 3292
rect 468996 3290 469052 3292
rect 469076 3290 469132 3292
rect 469156 3290 469212 3292
rect 469236 3290 469292 3292
rect 469316 3290 469372 3292
rect 468836 3238 468874 3290
rect 468874 3238 468886 3290
rect 468886 3238 468892 3290
rect 468916 3238 468938 3290
rect 468938 3238 468950 3290
rect 468950 3238 468972 3290
rect 468996 3238 469002 3290
rect 469002 3238 469014 3290
rect 469014 3238 469052 3290
rect 469076 3238 469078 3290
rect 469078 3238 469130 3290
rect 469130 3238 469132 3290
rect 469156 3238 469194 3290
rect 469194 3238 469206 3290
rect 469206 3238 469212 3290
rect 469236 3238 469258 3290
rect 469258 3238 469270 3290
rect 469270 3238 469292 3290
rect 469316 3238 469322 3290
rect 469322 3238 469334 3290
rect 469334 3238 469372 3290
rect 468836 3236 468892 3238
rect 468916 3236 468972 3238
rect 468996 3236 469052 3238
rect 469076 3236 469132 3238
rect 469156 3236 469212 3238
rect 469236 3236 469292 3238
rect 469316 3236 469372 3238
rect 468836 2202 468892 2204
rect 468916 2202 468972 2204
rect 468996 2202 469052 2204
rect 469076 2202 469132 2204
rect 469156 2202 469212 2204
rect 469236 2202 469292 2204
rect 469316 2202 469372 2204
rect 468836 2150 468874 2202
rect 468874 2150 468886 2202
rect 468886 2150 468892 2202
rect 468916 2150 468938 2202
rect 468938 2150 468950 2202
rect 468950 2150 468972 2202
rect 468996 2150 469002 2202
rect 469002 2150 469014 2202
rect 469014 2150 469052 2202
rect 469076 2150 469078 2202
rect 469078 2150 469130 2202
rect 469130 2150 469132 2202
rect 469156 2150 469194 2202
rect 469194 2150 469206 2202
rect 469206 2150 469212 2202
rect 469236 2150 469258 2202
rect 469258 2150 469270 2202
rect 469270 2150 469292 2202
rect 469316 2150 469322 2202
rect 469322 2150 469334 2202
rect 469334 2150 469372 2202
rect 468836 2148 468892 2150
rect 468916 2148 468972 2150
rect 468996 2148 469052 2150
rect 469076 2148 469132 2150
rect 469156 2148 469212 2150
rect 469236 2148 469292 2150
rect 469316 2148 469372 2150
rect 486836 6010 486892 6012
rect 486916 6010 486972 6012
rect 486996 6010 487052 6012
rect 487076 6010 487132 6012
rect 487156 6010 487212 6012
rect 487236 6010 487292 6012
rect 487316 6010 487372 6012
rect 486836 5958 486874 6010
rect 486874 5958 486886 6010
rect 486886 5958 486892 6010
rect 486916 5958 486938 6010
rect 486938 5958 486950 6010
rect 486950 5958 486972 6010
rect 486996 5958 487002 6010
rect 487002 5958 487014 6010
rect 487014 5958 487052 6010
rect 487076 5958 487078 6010
rect 487078 5958 487130 6010
rect 487130 5958 487132 6010
rect 487156 5958 487194 6010
rect 487194 5958 487206 6010
rect 487206 5958 487212 6010
rect 487236 5958 487258 6010
rect 487258 5958 487270 6010
rect 487270 5958 487292 6010
rect 487316 5958 487322 6010
rect 487322 5958 487334 6010
rect 487334 5958 487372 6010
rect 486836 5956 486892 5958
rect 486916 5956 486972 5958
rect 486996 5956 487052 5958
rect 487076 5956 487132 5958
rect 487156 5956 487212 5958
rect 487236 5956 487292 5958
rect 487316 5956 487372 5958
rect 486836 4922 486892 4924
rect 486916 4922 486972 4924
rect 486996 4922 487052 4924
rect 487076 4922 487132 4924
rect 487156 4922 487212 4924
rect 487236 4922 487292 4924
rect 487316 4922 487372 4924
rect 486836 4870 486874 4922
rect 486874 4870 486886 4922
rect 486886 4870 486892 4922
rect 486916 4870 486938 4922
rect 486938 4870 486950 4922
rect 486950 4870 486972 4922
rect 486996 4870 487002 4922
rect 487002 4870 487014 4922
rect 487014 4870 487052 4922
rect 487076 4870 487078 4922
rect 487078 4870 487130 4922
rect 487130 4870 487132 4922
rect 487156 4870 487194 4922
rect 487194 4870 487206 4922
rect 487206 4870 487212 4922
rect 487236 4870 487258 4922
rect 487258 4870 487270 4922
rect 487270 4870 487292 4922
rect 487316 4870 487322 4922
rect 487322 4870 487334 4922
rect 487334 4870 487372 4922
rect 486836 4868 486892 4870
rect 486916 4868 486972 4870
rect 486996 4868 487052 4870
rect 487076 4868 487132 4870
rect 487156 4868 487212 4870
rect 487236 4868 487292 4870
rect 487316 4868 487372 4870
rect 486836 3834 486892 3836
rect 486916 3834 486972 3836
rect 486996 3834 487052 3836
rect 487076 3834 487132 3836
rect 487156 3834 487212 3836
rect 487236 3834 487292 3836
rect 487316 3834 487372 3836
rect 486836 3782 486874 3834
rect 486874 3782 486886 3834
rect 486886 3782 486892 3834
rect 486916 3782 486938 3834
rect 486938 3782 486950 3834
rect 486950 3782 486972 3834
rect 486996 3782 487002 3834
rect 487002 3782 487014 3834
rect 487014 3782 487052 3834
rect 487076 3782 487078 3834
rect 487078 3782 487130 3834
rect 487130 3782 487132 3834
rect 487156 3782 487194 3834
rect 487194 3782 487206 3834
rect 487206 3782 487212 3834
rect 487236 3782 487258 3834
rect 487258 3782 487270 3834
rect 487270 3782 487292 3834
rect 487316 3782 487322 3834
rect 487322 3782 487334 3834
rect 487334 3782 487372 3834
rect 486836 3780 486892 3782
rect 486916 3780 486972 3782
rect 486996 3780 487052 3782
rect 487076 3780 487132 3782
rect 487156 3780 487212 3782
rect 487236 3780 487292 3782
rect 487316 3780 487372 3782
rect 486836 2746 486892 2748
rect 486916 2746 486972 2748
rect 486996 2746 487052 2748
rect 487076 2746 487132 2748
rect 487156 2746 487212 2748
rect 487236 2746 487292 2748
rect 487316 2746 487372 2748
rect 486836 2694 486874 2746
rect 486874 2694 486886 2746
rect 486886 2694 486892 2746
rect 486916 2694 486938 2746
rect 486938 2694 486950 2746
rect 486950 2694 486972 2746
rect 486996 2694 487002 2746
rect 487002 2694 487014 2746
rect 487014 2694 487052 2746
rect 487076 2694 487078 2746
rect 487078 2694 487130 2746
rect 487130 2694 487132 2746
rect 487156 2694 487194 2746
rect 487194 2694 487206 2746
rect 487206 2694 487212 2746
rect 487236 2694 487258 2746
rect 487258 2694 487270 2746
rect 487270 2694 487292 2746
rect 487316 2694 487322 2746
rect 487322 2694 487334 2746
rect 487334 2694 487372 2746
rect 486836 2692 486892 2694
rect 486916 2692 486972 2694
rect 486996 2692 487052 2694
rect 487076 2692 487132 2694
rect 487156 2692 487212 2694
rect 487236 2692 487292 2694
rect 487316 2692 487372 2694
rect 504836 5466 504892 5468
rect 504916 5466 504972 5468
rect 504996 5466 505052 5468
rect 505076 5466 505132 5468
rect 505156 5466 505212 5468
rect 505236 5466 505292 5468
rect 505316 5466 505372 5468
rect 504836 5414 504874 5466
rect 504874 5414 504886 5466
rect 504886 5414 504892 5466
rect 504916 5414 504938 5466
rect 504938 5414 504950 5466
rect 504950 5414 504972 5466
rect 504996 5414 505002 5466
rect 505002 5414 505014 5466
rect 505014 5414 505052 5466
rect 505076 5414 505078 5466
rect 505078 5414 505130 5466
rect 505130 5414 505132 5466
rect 505156 5414 505194 5466
rect 505194 5414 505206 5466
rect 505206 5414 505212 5466
rect 505236 5414 505258 5466
rect 505258 5414 505270 5466
rect 505270 5414 505292 5466
rect 505316 5414 505322 5466
rect 505322 5414 505334 5466
rect 505334 5414 505372 5466
rect 504836 5412 504892 5414
rect 504916 5412 504972 5414
rect 504996 5412 505052 5414
rect 505076 5412 505132 5414
rect 505156 5412 505212 5414
rect 505236 5412 505292 5414
rect 505316 5412 505372 5414
rect 504836 4378 504892 4380
rect 504916 4378 504972 4380
rect 504996 4378 505052 4380
rect 505076 4378 505132 4380
rect 505156 4378 505212 4380
rect 505236 4378 505292 4380
rect 505316 4378 505372 4380
rect 504836 4326 504874 4378
rect 504874 4326 504886 4378
rect 504886 4326 504892 4378
rect 504916 4326 504938 4378
rect 504938 4326 504950 4378
rect 504950 4326 504972 4378
rect 504996 4326 505002 4378
rect 505002 4326 505014 4378
rect 505014 4326 505052 4378
rect 505076 4326 505078 4378
rect 505078 4326 505130 4378
rect 505130 4326 505132 4378
rect 505156 4326 505194 4378
rect 505194 4326 505206 4378
rect 505206 4326 505212 4378
rect 505236 4326 505258 4378
rect 505258 4326 505270 4378
rect 505270 4326 505292 4378
rect 505316 4326 505322 4378
rect 505322 4326 505334 4378
rect 505334 4326 505372 4378
rect 504836 4324 504892 4326
rect 504916 4324 504972 4326
rect 504996 4324 505052 4326
rect 505076 4324 505132 4326
rect 505156 4324 505212 4326
rect 505236 4324 505292 4326
rect 505316 4324 505372 4326
rect 504836 3290 504892 3292
rect 504916 3290 504972 3292
rect 504996 3290 505052 3292
rect 505076 3290 505132 3292
rect 505156 3290 505212 3292
rect 505236 3290 505292 3292
rect 505316 3290 505372 3292
rect 504836 3238 504874 3290
rect 504874 3238 504886 3290
rect 504886 3238 504892 3290
rect 504916 3238 504938 3290
rect 504938 3238 504950 3290
rect 504950 3238 504972 3290
rect 504996 3238 505002 3290
rect 505002 3238 505014 3290
rect 505014 3238 505052 3290
rect 505076 3238 505078 3290
rect 505078 3238 505130 3290
rect 505130 3238 505132 3290
rect 505156 3238 505194 3290
rect 505194 3238 505206 3290
rect 505206 3238 505212 3290
rect 505236 3238 505258 3290
rect 505258 3238 505270 3290
rect 505270 3238 505292 3290
rect 505316 3238 505322 3290
rect 505322 3238 505334 3290
rect 505334 3238 505372 3290
rect 504836 3236 504892 3238
rect 504916 3236 504972 3238
rect 504996 3236 505052 3238
rect 505076 3236 505132 3238
rect 505156 3236 505212 3238
rect 505236 3236 505292 3238
rect 505316 3236 505372 3238
rect 504836 2202 504892 2204
rect 504916 2202 504972 2204
rect 504996 2202 505052 2204
rect 505076 2202 505132 2204
rect 505156 2202 505212 2204
rect 505236 2202 505292 2204
rect 505316 2202 505372 2204
rect 504836 2150 504874 2202
rect 504874 2150 504886 2202
rect 504886 2150 504892 2202
rect 504916 2150 504938 2202
rect 504938 2150 504950 2202
rect 504950 2150 504972 2202
rect 504996 2150 505002 2202
rect 505002 2150 505014 2202
rect 505014 2150 505052 2202
rect 505076 2150 505078 2202
rect 505078 2150 505130 2202
rect 505130 2150 505132 2202
rect 505156 2150 505194 2202
rect 505194 2150 505206 2202
rect 505206 2150 505212 2202
rect 505236 2150 505258 2202
rect 505258 2150 505270 2202
rect 505270 2150 505292 2202
rect 505316 2150 505322 2202
rect 505322 2150 505334 2202
rect 505334 2150 505372 2202
rect 504836 2148 504892 2150
rect 504916 2148 504972 2150
rect 504996 2148 505052 2150
rect 505076 2148 505132 2150
rect 505156 2148 505212 2150
rect 505236 2148 505292 2150
rect 505316 2148 505372 2150
rect 522836 6010 522892 6012
rect 522916 6010 522972 6012
rect 522996 6010 523052 6012
rect 523076 6010 523132 6012
rect 523156 6010 523212 6012
rect 523236 6010 523292 6012
rect 523316 6010 523372 6012
rect 522836 5958 522874 6010
rect 522874 5958 522886 6010
rect 522886 5958 522892 6010
rect 522916 5958 522938 6010
rect 522938 5958 522950 6010
rect 522950 5958 522972 6010
rect 522996 5958 523002 6010
rect 523002 5958 523014 6010
rect 523014 5958 523052 6010
rect 523076 5958 523078 6010
rect 523078 5958 523130 6010
rect 523130 5958 523132 6010
rect 523156 5958 523194 6010
rect 523194 5958 523206 6010
rect 523206 5958 523212 6010
rect 523236 5958 523258 6010
rect 523258 5958 523270 6010
rect 523270 5958 523292 6010
rect 523316 5958 523322 6010
rect 523322 5958 523334 6010
rect 523334 5958 523372 6010
rect 522836 5956 522892 5958
rect 522916 5956 522972 5958
rect 522996 5956 523052 5958
rect 523076 5956 523132 5958
rect 523156 5956 523212 5958
rect 523236 5956 523292 5958
rect 523316 5956 523372 5958
rect 522836 4922 522892 4924
rect 522916 4922 522972 4924
rect 522996 4922 523052 4924
rect 523076 4922 523132 4924
rect 523156 4922 523212 4924
rect 523236 4922 523292 4924
rect 523316 4922 523372 4924
rect 522836 4870 522874 4922
rect 522874 4870 522886 4922
rect 522886 4870 522892 4922
rect 522916 4870 522938 4922
rect 522938 4870 522950 4922
rect 522950 4870 522972 4922
rect 522996 4870 523002 4922
rect 523002 4870 523014 4922
rect 523014 4870 523052 4922
rect 523076 4870 523078 4922
rect 523078 4870 523130 4922
rect 523130 4870 523132 4922
rect 523156 4870 523194 4922
rect 523194 4870 523206 4922
rect 523206 4870 523212 4922
rect 523236 4870 523258 4922
rect 523258 4870 523270 4922
rect 523270 4870 523292 4922
rect 523316 4870 523322 4922
rect 523322 4870 523334 4922
rect 523334 4870 523372 4922
rect 522836 4868 522892 4870
rect 522916 4868 522972 4870
rect 522996 4868 523052 4870
rect 523076 4868 523132 4870
rect 523156 4868 523212 4870
rect 523236 4868 523292 4870
rect 523316 4868 523372 4870
rect 522836 3834 522892 3836
rect 522916 3834 522972 3836
rect 522996 3834 523052 3836
rect 523076 3834 523132 3836
rect 523156 3834 523212 3836
rect 523236 3834 523292 3836
rect 523316 3834 523372 3836
rect 522836 3782 522874 3834
rect 522874 3782 522886 3834
rect 522886 3782 522892 3834
rect 522916 3782 522938 3834
rect 522938 3782 522950 3834
rect 522950 3782 522972 3834
rect 522996 3782 523002 3834
rect 523002 3782 523014 3834
rect 523014 3782 523052 3834
rect 523076 3782 523078 3834
rect 523078 3782 523130 3834
rect 523130 3782 523132 3834
rect 523156 3782 523194 3834
rect 523194 3782 523206 3834
rect 523206 3782 523212 3834
rect 523236 3782 523258 3834
rect 523258 3782 523270 3834
rect 523270 3782 523292 3834
rect 523316 3782 523322 3834
rect 523322 3782 523334 3834
rect 523334 3782 523372 3834
rect 522836 3780 522892 3782
rect 522916 3780 522972 3782
rect 522996 3780 523052 3782
rect 523076 3780 523132 3782
rect 523156 3780 523212 3782
rect 523236 3780 523292 3782
rect 523316 3780 523372 3782
rect 522836 2746 522892 2748
rect 522916 2746 522972 2748
rect 522996 2746 523052 2748
rect 523076 2746 523132 2748
rect 523156 2746 523212 2748
rect 523236 2746 523292 2748
rect 523316 2746 523372 2748
rect 522836 2694 522874 2746
rect 522874 2694 522886 2746
rect 522886 2694 522892 2746
rect 522916 2694 522938 2746
rect 522938 2694 522950 2746
rect 522950 2694 522972 2746
rect 522996 2694 523002 2746
rect 523002 2694 523014 2746
rect 523014 2694 523052 2746
rect 523076 2694 523078 2746
rect 523078 2694 523130 2746
rect 523130 2694 523132 2746
rect 523156 2694 523194 2746
rect 523194 2694 523206 2746
rect 523206 2694 523212 2746
rect 523236 2694 523258 2746
rect 523258 2694 523270 2746
rect 523270 2694 523292 2746
rect 523316 2694 523322 2746
rect 523322 2694 523334 2746
rect 523334 2694 523372 2746
rect 522836 2692 522892 2694
rect 522916 2692 522972 2694
rect 522996 2692 523052 2694
rect 523076 2692 523132 2694
rect 523156 2692 523212 2694
rect 523236 2692 523292 2694
rect 523316 2692 523372 2694
rect 540836 5466 540892 5468
rect 540916 5466 540972 5468
rect 540996 5466 541052 5468
rect 541076 5466 541132 5468
rect 541156 5466 541212 5468
rect 541236 5466 541292 5468
rect 541316 5466 541372 5468
rect 540836 5414 540874 5466
rect 540874 5414 540886 5466
rect 540886 5414 540892 5466
rect 540916 5414 540938 5466
rect 540938 5414 540950 5466
rect 540950 5414 540972 5466
rect 540996 5414 541002 5466
rect 541002 5414 541014 5466
rect 541014 5414 541052 5466
rect 541076 5414 541078 5466
rect 541078 5414 541130 5466
rect 541130 5414 541132 5466
rect 541156 5414 541194 5466
rect 541194 5414 541206 5466
rect 541206 5414 541212 5466
rect 541236 5414 541258 5466
rect 541258 5414 541270 5466
rect 541270 5414 541292 5466
rect 541316 5414 541322 5466
rect 541322 5414 541334 5466
rect 541334 5414 541372 5466
rect 540836 5412 540892 5414
rect 540916 5412 540972 5414
rect 540996 5412 541052 5414
rect 541076 5412 541132 5414
rect 541156 5412 541212 5414
rect 541236 5412 541292 5414
rect 541316 5412 541372 5414
rect 540836 4378 540892 4380
rect 540916 4378 540972 4380
rect 540996 4378 541052 4380
rect 541076 4378 541132 4380
rect 541156 4378 541212 4380
rect 541236 4378 541292 4380
rect 541316 4378 541372 4380
rect 540836 4326 540874 4378
rect 540874 4326 540886 4378
rect 540886 4326 540892 4378
rect 540916 4326 540938 4378
rect 540938 4326 540950 4378
rect 540950 4326 540972 4378
rect 540996 4326 541002 4378
rect 541002 4326 541014 4378
rect 541014 4326 541052 4378
rect 541076 4326 541078 4378
rect 541078 4326 541130 4378
rect 541130 4326 541132 4378
rect 541156 4326 541194 4378
rect 541194 4326 541206 4378
rect 541206 4326 541212 4378
rect 541236 4326 541258 4378
rect 541258 4326 541270 4378
rect 541270 4326 541292 4378
rect 541316 4326 541322 4378
rect 541322 4326 541334 4378
rect 541334 4326 541372 4378
rect 540836 4324 540892 4326
rect 540916 4324 540972 4326
rect 540996 4324 541052 4326
rect 541076 4324 541132 4326
rect 541156 4324 541212 4326
rect 541236 4324 541292 4326
rect 541316 4324 541372 4326
rect 540836 3290 540892 3292
rect 540916 3290 540972 3292
rect 540996 3290 541052 3292
rect 541076 3290 541132 3292
rect 541156 3290 541212 3292
rect 541236 3290 541292 3292
rect 541316 3290 541372 3292
rect 540836 3238 540874 3290
rect 540874 3238 540886 3290
rect 540886 3238 540892 3290
rect 540916 3238 540938 3290
rect 540938 3238 540950 3290
rect 540950 3238 540972 3290
rect 540996 3238 541002 3290
rect 541002 3238 541014 3290
rect 541014 3238 541052 3290
rect 541076 3238 541078 3290
rect 541078 3238 541130 3290
rect 541130 3238 541132 3290
rect 541156 3238 541194 3290
rect 541194 3238 541206 3290
rect 541206 3238 541212 3290
rect 541236 3238 541258 3290
rect 541258 3238 541270 3290
rect 541270 3238 541292 3290
rect 541316 3238 541322 3290
rect 541322 3238 541334 3290
rect 541334 3238 541372 3290
rect 540836 3236 540892 3238
rect 540916 3236 540972 3238
rect 540996 3236 541052 3238
rect 541076 3236 541132 3238
rect 541156 3236 541212 3238
rect 541236 3236 541292 3238
rect 541316 3236 541372 3238
rect 540836 2202 540892 2204
rect 540916 2202 540972 2204
rect 540996 2202 541052 2204
rect 541076 2202 541132 2204
rect 541156 2202 541212 2204
rect 541236 2202 541292 2204
rect 541316 2202 541372 2204
rect 540836 2150 540874 2202
rect 540874 2150 540886 2202
rect 540886 2150 540892 2202
rect 540916 2150 540938 2202
rect 540938 2150 540950 2202
rect 540950 2150 540972 2202
rect 540996 2150 541002 2202
rect 541002 2150 541014 2202
rect 541014 2150 541052 2202
rect 541076 2150 541078 2202
rect 541078 2150 541130 2202
rect 541130 2150 541132 2202
rect 541156 2150 541194 2202
rect 541194 2150 541206 2202
rect 541206 2150 541212 2202
rect 541236 2150 541258 2202
rect 541258 2150 541270 2202
rect 541270 2150 541292 2202
rect 541316 2150 541322 2202
rect 541322 2150 541334 2202
rect 541334 2150 541372 2202
rect 540836 2148 540892 2150
rect 540916 2148 540972 2150
rect 540996 2148 541052 2150
rect 541076 2148 541132 2150
rect 541156 2148 541212 2150
rect 541236 2148 541292 2150
rect 541316 2148 541372 2150
rect 558836 6010 558892 6012
rect 558916 6010 558972 6012
rect 558996 6010 559052 6012
rect 559076 6010 559132 6012
rect 559156 6010 559212 6012
rect 559236 6010 559292 6012
rect 559316 6010 559372 6012
rect 558836 5958 558874 6010
rect 558874 5958 558886 6010
rect 558886 5958 558892 6010
rect 558916 5958 558938 6010
rect 558938 5958 558950 6010
rect 558950 5958 558972 6010
rect 558996 5958 559002 6010
rect 559002 5958 559014 6010
rect 559014 5958 559052 6010
rect 559076 5958 559078 6010
rect 559078 5958 559130 6010
rect 559130 5958 559132 6010
rect 559156 5958 559194 6010
rect 559194 5958 559206 6010
rect 559206 5958 559212 6010
rect 559236 5958 559258 6010
rect 559258 5958 559270 6010
rect 559270 5958 559292 6010
rect 559316 5958 559322 6010
rect 559322 5958 559334 6010
rect 559334 5958 559372 6010
rect 558836 5956 558892 5958
rect 558916 5956 558972 5958
rect 558996 5956 559052 5958
rect 559076 5956 559132 5958
rect 559156 5956 559212 5958
rect 559236 5956 559292 5958
rect 559316 5956 559372 5958
rect 558836 4922 558892 4924
rect 558916 4922 558972 4924
rect 558996 4922 559052 4924
rect 559076 4922 559132 4924
rect 559156 4922 559212 4924
rect 559236 4922 559292 4924
rect 559316 4922 559372 4924
rect 558836 4870 558874 4922
rect 558874 4870 558886 4922
rect 558886 4870 558892 4922
rect 558916 4870 558938 4922
rect 558938 4870 558950 4922
rect 558950 4870 558972 4922
rect 558996 4870 559002 4922
rect 559002 4870 559014 4922
rect 559014 4870 559052 4922
rect 559076 4870 559078 4922
rect 559078 4870 559130 4922
rect 559130 4870 559132 4922
rect 559156 4870 559194 4922
rect 559194 4870 559206 4922
rect 559206 4870 559212 4922
rect 559236 4870 559258 4922
rect 559258 4870 559270 4922
rect 559270 4870 559292 4922
rect 559316 4870 559322 4922
rect 559322 4870 559334 4922
rect 559334 4870 559372 4922
rect 558836 4868 558892 4870
rect 558916 4868 558972 4870
rect 558996 4868 559052 4870
rect 559076 4868 559132 4870
rect 559156 4868 559212 4870
rect 559236 4868 559292 4870
rect 559316 4868 559372 4870
rect 558836 3834 558892 3836
rect 558916 3834 558972 3836
rect 558996 3834 559052 3836
rect 559076 3834 559132 3836
rect 559156 3834 559212 3836
rect 559236 3834 559292 3836
rect 559316 3834 559372 3836
rect 558836 3782 558874 3834
rect 558874 3782 558886 3834
rect 558886 3782 558892 3834
rect 558916 3782 558938 3834
rect 558938 3782 558950 3834
rect 558950 3782 558972 3834
rect 558996 3782 559002 3834
rect 559002 3782 559014 3834
rect 559014 3782 559052 3834
rect 559076 3782 559078 3834
rect 559078 3782 559130 3834
rect 559130 3782 559132 3834
rect 559156 3782 559194 3834
rect 559194 3782 559206 3834
rect 559206 3782 559212 3834
rect 559236 3782 559258 3834
rect 559258 3782 559270 3834
rect 559270 3782 559292 3834
rect 559316 3782 559322 3834
rect 559322 3782 559334 3834
rect 559334 3782 559372 3834
rect 558836 3780 558892 3782
rect 558916 3780 558972 3782
rect 558996 3780 559052 3782
rect 559076 3780 559132 3782
rect 559156 3780 559212 3782
rect 559236 3780 559292 3782
rect 559316 3780 559372 3782
rect 558836 2746 558892 2748
rect 558916 2746 558972 2748
rect 558996 2746 559052 2748
rect 559076 2746 559132 2748
rect 559156 2746 559212 2748
rect 559236 2746 559292 2748
rect 559316 2746 559372 2748
rect 558836 2694 558874 2746
rect 558874 2694 558886 2746
rect 558886 2694 558892 2746
rect 558916 2694 558938 2746
rect 558938 2694 558950 2746
rect 558950 2694 558972 2746
rect 558996 2694 559002 2746
rect 559002 2694 559014 2746
rect 559014 2694 559052 2746
rect 559076 2694 559078 2746
rect 559078 2694 559130 2746
rect 559130 2694 559132 2746
rect 559156 2694 559194 2746
rect 559194 2694 559206 2746
rect 559206 2694 559212 2746
rect 559236 2694 559258 2746
rect 559258 2694 559270 2746
rect 559270 2694 559292 2746
rect 559316 2694 559322 2746
rect 559322 2694 559334 2746
rect 559334 2694 559372 2746
rect 558836 2692 558892 2694
rect 558916 2692 558972 2694
rect 558996 2692 559052 2694
rect 559076 2692 559132 2694
rect 559156 2692 559212 2694
rect 559236 2692 559292 2694
rect 559316 2692 559372 2694
rect 561678 3460 561734 3496
rect 576836 5466 576892 5468
rect 576916 5466 576972 5468
rect 576996 5466 577052 5468
rect 577076 5466 577132 5468
rect 577156 5466 577212 5468
rect 577236 5466 577292 5468
rect 577316 5466 577372 5468
rect 576836 5414 576874 5466
rect 576874 5414 576886 5466
rect 576886 5414 576892 5466
rect 576916 5414 576938 5466
rect 576938 5414 576950 5466
rect 576950 5414 576972 5466
rect 576996 5414 577002 5466
rect 577002 5414 577014 5466
rect 577014 5414 577052 5466
rect 577076 5414 577078 5466
rect 577078 5414 577130 5466
rect 577130 5414 577132 5466
rect 577156 5414 577194 5466
rect 577194 5414 577206 5466
rect 577206 5414 577212 5466
rect 577236 5414 577258 5466
rect 577258 5414 577270 5466
rect 577270 5414 577292 5466
rect 577316 5414 577322 5466
rect 577322 5414 577334 5466
rect 577334 5414 577372 5466
rect 576836 5412 576892 5414
rect 576916 5412 576972 5414
rect 576996 5412 577052 5414
rect 577076 5412 577132 5414
rect 577156 5412 577212 5414
rect 577236 5412 577292 5414
rect 577316 5412 577372 5414
rect 576836 4378 576892 4380
rect 576916 4378 576972 4380
rect 576996 4378 577052 4380
rect 577076 4378 577132 4380
rect 577156 4378 577212 4380
rect 577236 4378 577292 4380
rect 577316 4378 577372 4380
rect 576836 4326 576874 4378
rect 576874 4326 576886 4378
rect 576886 4326 576892 4378
rect 576916 4326 576938 4378
rect 576938 4326 576950 4378
rect 576950 4326 576972 4378
rect 576996 4326 577002 4378
rect 577002 4326 577014 4378
rect 577014 4326 577052 4378
rect 577076 4326 577078 4378
rect 577078 4326 577130 4378
rect 577130 4326 577132 4378
rect 577156 4326 577194 4378
rect 577194 4326 577206 4378
rect 577206 4326 577212 4378
rect 577236 4326 577258 4378
rect 577258 4326 577270 4378
rect 577270 4326 577292 4378
rect 577316 4326 577322 4378
rect 577322 4326 577334 4378
rect 577334 4326 577372 4378
rect 576836 4324 576892 4326
rect 576916 4324 576972 4326
rect 576996 4324 577052 4326
rect 577076 4324 577132 4326
rect 577156 4324 577212 4326
rect 577236 4324 577292 4326
rect 577316 4324 577372 4326
rect 561678 3440 561680 3460
rect 561680 3440 561732 3460
rect 561732 3440 561734 3460
rect 564530 3440 564586 3496
rect 576836 3290 576892 3292
rect 576916 3290 576972 3292
rect 576996 3290 577052 3292
rect 577076 3290 577132 3292
rect 577156 3290 577212 3292
rect 577236 3290 577292 3292
rect 577316 3290 577372 3292
rect 576836 3238 576874 3290
rect 576874 3238 576886 3290
rect 576886 3238 576892 3290
rect 576916 3238 576938 3290
rect 576938 3238 576950 3290
rect 576950 3238 576972 3290
rect 576996 3238 577002 3290
rect 577002 3238 577014 3290
rect 577014 3238 577052 3290
rect 577076 3238 577078 3290
rect 577078 3238 577130 3290
rect 577130 3238 577132 3290
rect 577156 3238 577194 3290
rect 577194 3238 577206 3290
rect 577206 3238 577212 3290
rect 577236 3238 577258 3290
rect 577258 3238 577270 3290
rect 577270 3238 577292 3290
rect 577316 3238 577322 3290
rect 577322 3238 577334 3290
rect 577334 3238 577372 3290
rect 576836 3236 576892 3238
rect 576916 3236 576972 3238
rect 576996 3236 577052 3238
rect 577076 3236 577132 3238
rect 577156 3236 577212 3238
rect 577236 3236 577292 3238
rect 577316 3236 577372 3238
rect 576836 2202 576892 2204
rect 576916 2202 576972 2204
rect 576996 2202 577052 2204
rect 577076 2202 577132 2204
rect 577156 2202 577212 2204
rect 577236 2202 577292 2204
rect 577316 2202 577372 2204
rect 576836 2150 576874 2202
rect 576874 2150 576886 2202
rect 576886 2150 576892 2202
rect 576916 2150 576938 2202
rect 576938 2150 576950 2202
rect 576950 2150 576972 2202
rect 576996 2150 577002 2202
rect 577002 2150 577014 2202
rect 577014 2150 577052 2202
rect 577076 2150 577078 2202
rect 577078 2150 577130 2202
rect 577130 2150 577132 2202
rect 577156 2150 577194 2202
rect 577194 2150 577206 2202
rect 577206 2150 577212 2202
rect 577236 2150 577258 2202
rect 577258 2150 577270 2202
rect 577270 2150 577292 2202
rect 577316 2150 577322 2202
rect 577322 2150 577334 2202
rect 577334 2150 577372 2202
rect 576836 2148 576892 2150
rect 576916 2148 576972 2150
rect 576996 2148 577052 2150
rect 577076 2148 577132 2150
rect 577156 2148 577212 2150
rect 577236 2148 577292 2150
rect 577316 2148 577372 2150
<< metal3 >>
rect 36804 701792 37404 701793
rect 36804 701728 36832 701792
rect 36896 701728 36912 701792
rect 36976 701728 36992 701792
rect 37056 701728 37072 701792
rect 37136 701728 37152 701792
rect 37216 701728 37232 701792
rect 37296 701728 37312 701792
rect 37376 701728 37404 701792
rect 36804 701727 37404 701728
rect 72804 701792 73404 701793
rect 72804 701728 72832 701792
rect 72896 701728 72912 701792
rect 72976 701728 72992 701792
rect 73056 701728 73072 701792
rect 73136 701728 73152 701792
rect 73216 701728 73232 701792
rect 73296 701728 73312 701792
rect 73376 701728 73404 701792
rect 72804 701727 73404 701728
rect 108804 701792 109404 701793
rect 108804 701728 108832 701792
rect 108896 701728 108912 701792
rect 108976 701728 108992 701792
rect 109056 701728 109072 701792
rect 109136 701728 109152 701792
rect 109216 701728 109232 701792
rect 109296 701728 109312 701792
rect 109376 701728 109404 701792
rect 108804 701727 109404 701728
rect 144804 701792 145404 701793
rect 144804 701728 144832 701792
rect 144896 701728 144912 701792
rect 144976 701728 144992 701792
rect 145056 701728 145072 701792
rect 145136 701728 145152 701792
rect 145216 701728 145232 701792
rect 145296 701728 145312 701792
rect 145376 701728 145404 701792
rect 144804 701727 145404 701728
rect 180804 701792 181404 701793
rect 180804 701728 180832 701792
rect 180896 701728 180912 701792
rect 180976 701728 180992 701792
rect 181056 701728 181072 701792
rect 181136 701728 181152 701792
rect 181216 701728 181232 701792
rect 181296 701728 181312 701792
rect 181376 701728 181404 701792
rect 180804 701727 181404 701728
rect 216804 701792 217404 701793
rect 216804 701728 216832 701792
rect 216896 701728 216912 701792
rect 216976 701728 216992 701792
rect 217056 701728 217072 701792
rect 217136 701728 217152 701792
rect 217216 701728 217232 701792
rect 217296 701728 217312 701792
rect 217376 701728 217404 701792
rect 216804 701727 217404 701728
rect 252804 701792 253404 701793
rect 252804 701728 252832 701792
rect 252896 701728 252912 701792
rect 252976 701728 252992 701792
rect 253056 701728 253072 701792
rect 253136 701728 253152 701792
rect 253216 701728 253232 701792
rect 253296 701728 253312 701792
rect 253376 701728 253404 701792
rect 252804 701727 253404 701728
rect 288804 701792 289404 701793
rect 288804 701728 288832 701792
rect 288896 701728 288912 701792
rect 288976 701728 288992 701792
rect 289056 701728 289072 701792
rect 289136 701728 289152 701792
rect 289216 701728 289232 701792
rect 289296 701728 289312 701792
rect 289376 701728 289404 701792
rect 288804 701727 289404 701728
rect 324804 701792 325404 701793
rect 324804 701728 324832 701792
rect 324896 701728 324912 701792
rect 324976 701728 324992 701792
rect 325056 701728 325072 701792
rect 325136 701728 325152 701792
rect 325216 701728 325232 701792
rect 325296 701728 325312 701792
rect 325376 701728 325404 701792
rect 324804 701727 325404 701728
rect 360804 701792 361404 701793
rect 360804 701728 360832 701792
rect 360896 701728 360912 701792
rect 360976 701728 360992 701792
rect 361056 701728 361072 701792
rect 361136 701728 361152 701792
rect 361216 701728 361232 701792
rect 361296 701728 361312 701792
rect 361376 701728 361404 701792
rect 360804 701727 361404 701728
rect 396804 701792 397404 701793
rect 396804 701728 396832 701792
rect 396896 701728 396912 701792
rect 396976 701728 396992 701792
rect 397056 701728 397072 701792
rect 397136 701728 397152 701792
rect 397216 701728 397232 701792
rect 397296 701728 397312 701792
rect 397376 701728 397404 701792
rect 396804 701727 397404 701728
rect 432804 701792 433404 701793
rect 432804 701728 432832 701792
rect 432896 701728 432912 701792
rect 432976 701728 432992 701792
rect 433056 701728 433072 701792
rect 433136 701728 433152 701792
rect 433216 701728 433232 701792
rect 433296 701728 433312 701792
rect 433376 701728 433404 701792
rect 432804 701727 433404 701728
rect 468804 701792 469404 701793
rect 468804 701728 468832 701792
rect 468896 701728 468912 701792
rect 468976 701728 468992 701792
rect 469056 701728 469072 701792
rect 469136 701728 469152 701792
rect 469216 701728 469232 701792
rect 469296 701728 469312 701792
rect 469376 701728 469404 701792
rect 468804 701727 469404 701728
rect 504804 701792 505404 701793
rect 504804 701728 504832 701792
rect 504896 701728 504912 701792
rect 504976 701728 504992 701792
rect 505056 701728 505072 701792
rect 505136 701728 505152 701792
rect 505216 701728 505232 701792
rect 505296 701728 505312 701792
rect 505376 701728 505404 701792
rect 504804 701727 505404 701728
rect 540804 701792 541404 701793
rect 540804 701728 540832 701792
rect 540896 701728 540912 701792
rect 540976 701728 540992 701792
rect 541056 701728 541072 701792
rect 541136 701728 541152 701792
rect 541216 701728 541232 701792
rect 541296 701728 541312 701792
rect 541376 701728 541404 701792
rect 540804 701727 541404 701728
rect 576804 701792 577404 701793
rect 576804 701728 576832 701792
rect 576896 701728 576912 701792
rect 576976 701728 576992 701792
rect 577056 701728 577072 701792
rect 577136 701728 577152 701792
rect 577216 701728 577232 701792
rect 577296 701728 577312 701792
rect 577376 701728 577404 701792
rect 576804 701727 577404 701728
rect 18804 701248 19404 701249
rect 18804 701184 18832 701248
rect 18896 701184 18912 701248
rect 18976 701184 18992 701248
rect 19056 701184 19072 701248
rect 19136 701184 19152 701248
rect 19216 701184 19232 701248
rect 19296 701184 19312 701248
rect 19376 701184 19404 701248
rect 18804 701183 19404 701184
rect 54804 701248 55404 701249
rect 54804 701184 54832 701248
rect 54896 701184 54912 701248
rect 54976 701184 54992 701248
rect 55056 701184 55072 701248
rect 55136 701184 55152 701248
rect 55216 701184 55232 701248
rect 55296 701184 55312 701248
rect 55376 701184 55404 701248
rect 54804 701183 55404 701184
rect 90804 701248 91404 701249
rect 90804 701184 90832 701248
rect 90896 701184 90912 701248
rect 90976 701184 90992 701248
rect 91056 701184 91072 701248
rect 91136 701184 91152 701248
rect 91216 701184 91232 701248
rect 91296 701184 91312 701248
rect 91376 701184 91404 701248
rect 90804 701183 91404 701184
rect 126804 701248 127404 701249
rect 126804 701184 126832 701248
rect 126896 701184 126912 701248
rect 126976 701184 126992 701248
rect 127056 701184 127072 701248
rect 127136 701184 127152 701248
rect 127216 701184 127232 701248
rect 127296 701184 127312 701248
rect 127376 701184 127404 701248
rect 126804 701183 127404 701184
rect 162804 701248 163404 701249
rect 162804 701184 162832 701248
rect 162896 701184 162912 701248
rect 162976 701184 162992 701248
rect 163056 701184 163072 701248
rect 163136 701184 163152 701248
rect 163216 701184 163232 701248
rect 163296 701184 163312 701248
rect 163376 701184 163404 701248
rect 162804 701183 163404 701184
rect 198804 701248 199404 701249
rect 198804 701184 198832 701248
rect 198896 701184 198912 701248
rect 198976 701184 198992 701248
rect 199056 701184 199072 701248
rect 199136 701184 199152 701248
rect 199216 701184 199232 701248
rect 199296 701184 199312 701248
rect 199376 701184 199404 701248
rect 198804 701183 199404 701184
rect 234804 701248 235404 701249
rect 234804 701184 234832 701248
rect 234896 701184 234912 701248
rect 234976 701184 234992 701248
rect 235056 701184 235072 701248
rect 235136 701184 235152 701248
rect 235216 701184 235232 701248
rect 235296 701184 235312 701248
rect 235376 701184 235404 701248
rect 234804 701183 235404 701184
rect 270804 701248 271404 701249
rect 270804 701184 270832 701248
rect 270896 701184 270912 701248
rect 270976 701184 270992 701248
rect 271056 701184 271072 701248
rect 271136 701184 271152 701248
rect 271216 701184 271232 701248
rect 271296 701184 271312 701248
rect 271376 701184 271404 701248
rect 270804 701183 271404 701184
rect 306804 701248 307404 701249
rect 306804 701184 306832 701248
rect 306896 701184 306912 701248
rect 306976 701184 306992 701248
rect 307056 701184 307072 701248
rect 307136 701184 307152 701248
rect 307216 701184 307232 701248
rect 307296 701184 307312 701248
rect 307376 701184 307404 701248
rect 306804 701183 307404 701184
rect 342804 701248 343404 701249
rect 342804 701184 342832 701248
rect 342896 701184 342912 701248
rect 342976 701184 342992 701248
rect 343056 701184 343072 701248
rect 343136 701184 343152 701248
rect 343216 701184 343232 701248
rect 343296 701184 343312 701248
rect 343376 701184 343404 701248
rect 342804 701183 343404 701184
rect 378804 701248 379404 701249
rect 378804 701184 378832 701248
rect 378896 701184 378912 701248
rect 378976 701184 378992 701248
rect 379056 701184 379072 701248
rect 379136 701184 379152 701248
rect 379216 701184 379232 701248
rect 379296 701184 379312 701248
rect 379376 701184 379404 701248
rect 378804 701183 379404 701184
rect 414804 701248 415404 701249
rect 414804 701184 414832 701248
rect 414896 701184 414912 701248
rect 414976 701184 414992 701248
rect 415056 701184 415072 701248
rect 415136 701184 415152 701248
rect 415216 701184 415232 701248
rect 415296 701184 415312 701248
rect 415376 701184 415404 701248
rect 414804 701183 415404 701184
rect 450804 701248 451404 701249
rect 450804 701184 450832 701248
rect 450896 701184 450912 701248
rect 450976 701184 450992 701248
rect 451056 701184 451072 701248
rect 451136 701184 451152 701248
rect 451216 701184 451232 701248
rect 451296 701184 451312 701248
rect 451376 701184 451404 701248
rect 450804 701183 451404 701184
rect 486804 701248 487404 701249
rect 486804 701184 486832 701248
rect 486896 701184 486912 701248
rect 486976 701184 486992 701248
rect 487056 701184 487072 701248
rect 487136 701184 487152 701248
rect 487216 701184 487232 701248
rect 487296 701184 487312 701248
rect 487376 701184 487404 701248
rect 486804 701183 487404 701184
rect 522804 701248 523404 701249
rect 522804 701184 522832 701248
rect 522896 701184 522912 701248
rect 522976 701184 522992 701248
rect 523056 701184 523072 701248
rect 523136 701184 523152 701248
rect 523216 701184 523232 701248
rect 523296 701184 523312 701248
rect 523376 701184 523404 701248
rect 522804 701183 523404 701184
rect 558804 701248 559404 701249
rect 558804 701184 558832 701248
rect 558896 701184 558912 701248
rect 558976 701184 558992 701248
rect 559056 701184 559072 701248
rect 559136 701184 559152 701248
rect 559216 701184 559232 701248
rect 559296 701184 559312 701248
rect 559376 701184 559404 701248
rect 558804 701183 559404 701184
rect 40493 701042 40559 701045
rect 336917 701042 336983 701045
rect 40493 701040 336983 701042
rect 40493 700984 40498 701040
rect 40554 700984 336922 701040
rect 336978 700984 336983 701040
rect 40493 700982 336983 700984
rect 40493 700979 40559 700982
rect 336917 700979 336983 700982
rect 227989 700906 228055 700909
rect 527173 700906 527239 700909
rect 227989 700904 527239 700906
rect 227989 700848 227994 700904
rect 228050 700848 527178 700904
rect 527234 700848 527239 700904
rect 227989 700846 527239 700848
rect 227989 700843 228055 700846
rect 527173 700843 527239 700846
rect 36804 700704 37404 700705
rect 36804 700640 36832 700704
rect 36896 700640 36912 700704
rect 36976 700640 36992 700704
rect 37056 700640 37072 700704
rect 37136 700640 37152 700704
rect 37216 700640 37232 700704
rect 37296 700640 37312 700704
rect 37376 700640 37404 700704
rect 36804 700639 37404 700640
rect 72804 700704 73404 700705
rect 72804 700640 72832 700704
rect 72896 700640 72912 700704
rect 72976 700640 72992 700704
rect 73056 700640 73072 700704
rect 73136 700640 73152 700704
rect 73216 700640 73232 700704
rect 73296 700640 73312 700704
rect 73376 700640 73404 700704
rect 72804 700639 73404 700640
rect 108804 700704 109404 700705
rect 108804 700640 108832 700704
rect 108896 700640 108912 700704
rect 108976 700640 108992 700704
rect 109056 700640 109072 700704
rect 109136 700640 109152 700704
rect 109216 700640 109232 700704
rect 109296 700640 109312 700704
rect 109376 700640 109404 700704
rect 108804 700639 109404 700640
rect 144804 700704 145404 700705
rect 144804 700640 144832 700704
rect 144896 700640 144912 700704
rect 144976 700640 144992 700704
rect 145056 700640 145072 700704
rect 145136 700640 145152 700704
rect 145216 700640 145232 700704
rect 145296 700640 145312 700704
rect 145376 700640 145404 700704
rect 144804 700639 145404 700640
rect 180804 700704 181404 700705
rect 180804 700640 180832 700704
rect 180896 700640 180912 700704
rect 180976 700640 180992 700704
rect 181056 700640 181072 700704
rect 181136 700640 181152 700704
rect 181216 700640 181232 700704
rect 181296 700640 181312 700704
rect 181376 700640 181404 700704
rect 180804 700639 181404 700640
rect 216804 700704 217404 700705
rect 216804 700640 216832 700704
rect 216896 700640 216912 700704
rect 216976 700640 216992 700704
rect 217056 700640 217072 700704
rect 217136 700640 217152 700704
rect 217216 700640 217232 700704
rect 217296 700640 217312 700704
rect 217376 700640 217404 700704
rect 216804 700639 217404 700640
rect 252804 700704 253404 700705
rect 252804 700640 252832 700704
rect 252896 700640 252912 700704
rect 252976 700640 252992 700704
rect 253056 700640 253072 700704
rect 253136 700640 253152 700704
rect 253216 700640 253232 700704
rect 253296 700640 253312 700704
rect 253376 700640 253404 700704
rect 252804 700639 253404 700640
rect 288804 700704 289404 700705
rect 288804 700640 288832 700704
rect 288896 700640 288912 700704
rect 288976 700640 288992 700704
rect 289056 700640 289072 700704
rect 289136 700640 289152 700704
rect 289216 700640 289232 700704
rect 289296 700640 289312 700704
rect 289376 700640 289404 700704
rect 288804 700639 289404 700640
rect 324804 700704 325404 700705
rect 324804 700640 324832 700704
rect 324896 700640 324912 700704
rect 324976 700640 324992 700704
rect 325056 700640 325072 700704
rect 325136 700640 325152 700704
rect 325216 700640 325232 700704
rect 325296 700640 325312 700704
rect 325376 700640 325404 700704
rect 324804 700639 325404 700640
rect 360804 700704 361404 700705
rect 360804 700640 360832 700704
rect 360896 700640 360912 700704
rect 360976 700640 360992 700704
rect 361056 700640 361072 700704
rect 361136 700640 361152 700704
rect 361216 700640 361232 700704
rect 361296 700640 361312 700704
rect 361376 700640 361404 700704
rect 360804 700639 361404 700640
rect 396804 700704 397404 700705
rect 396804 700640 396832 700704
rect 396896 700640 396912 700704
rect 396976 700640 396992 700704
rect 397056 700640 397072 700704
rect 397136 700640 397152 700704
rect 397216 700640 397232 700704
rect 397296 700640 397312 700704
rect 397376 700640 397404 700704
rect 396804 700639 397404 700640
rect 432804 700704 433404 700705
rect 432804 700640 432832 700704
rect 432896 700640 432912 700704
rect 432976 700640 432992 700704
rect 433056 700640 433072 700704
rect 433136 700640 433152 700704
rect 433216 700640 433232 700704
rect 433296 700640 433312 700704
rect 433376 700640 433404 700704
rect 432804 700639 433404 700640
rect 468804 700704 469404 700705
rect 468804 700640 468832 700704
rect 468896 700640 468912 700704
rect 468976 700640 468992 700704
rect 469056 700640 469072 700704
rect 469136 700640 469152 700704
rect 469216 700640 469232 700704
rect 469296 700640 469312 700704
rect 469376 700640 469404 700704
rect 468804 700639 469404 700640
rect 504804 700704 505404 700705
rect 504804 700640 504832 700704
rect 504896 700640 504912 700704
rect 504976 700640 504992 700704
rect 505056 700640 505072 700704
rect 505136 700640 505152 700704
rect 505216 700640 505232 700704
rect 505296 700640 505312 700704
rect 505376 700640 505404 700704
rect 504804 700639 505404 700640
rect 540804 700704 541404 700705
rect 540804 700640 540832 700704
rect 540896 700640 540912 700704
rect 540976 700640 540992 700704
rect 541056 700640 541072 700704
rect 541136 700640 541152 700704
rect 541216 700640 541232 700704
rect 541296 700640 541312 700704
rect 541376 700640 541404 700704
rect 540804 700639 541404 700640
rect 576804 700704 577404 700705
rect 576804 700640 576832 700704
rect 576896 700640 576912 700704
rect 576976 700640 576992 700704
rect 577056 700640 577072 700704
rect 577136 700640 577152 700704
rect 577216 700640 577232 700704
rect 577296 700640 577312 700704
rect 577376 700640 577404 700704
rect 576804 700639 577404 700640
rect 24301 700498 24367 700501
rect 346301 700498 346367 700501
rect 24301 700496 346367 700498
rect 24301 700440 24306 700496
rect 24362 700440 346306 700496
rect 346362 700440 346367 700496
rect 24301 700438 346367 700440
rect 24301 700435 24367 700438
rect 346301 700435 346367 700438
rect 8109 700362 8175 700365
rect 341609 700362 341675 700365
rect 8109 700360 341675 700362
rect 8109 700304 8114 700360
rect 8170 700304 341614 700360
rect 341670 700304 341675 700360
rect 8109 700302 341675 700304
rect 8109 700299 8175 700302
rect 341609 700299 341675 700302
rect 296529 700226 296595 700229
rect 298645 700226 298711 700229
rect 296529 700224 298711 700226
rect 296529 700168 296534 700224
rect 296590 700168 298650 700224
rect 298706 700168 298711 700224
rect 296529 700166 298711 700168
rect 296529 700163 296595 700166
rect 298645 700163 298711 700166
rect 18804 700160 19404 700161
rect 18804 700096 18832 700160
rect 18896 700096 18912 700160
rect 18976 700096 18992 700160
rect 19056 700096 19072 700160
rect 19136 700096 19152 700160
rect 19216 700096 19232 700160
rect 19296 700096 19312 700160
rect 19376 700096 19404 700160
rect 18804 700095 19404 700096
rect 54804 700160 55404 700161
rect 54804 700096 54832 700160
rect 54896 700096 54912 700160
rect 54976 700096 54992 700160
rect 55056 700096 55072 700160
rect 55136 700096 55152 700160
rect 55216 700096 55232 700160
rect 55296 700096 55312 700160
rect 55376 700096 55404 700160
rect 54804 700095 55404 700096
rect 90804 700160 91404 700161
rect 90804 700096 90832 700160
rect 90896 700096 90912 700160
rect 90976 700096 90992 700160
rect 91056 700096 91072 700160
rect 91136 700096 91152 700160
rect 91216 700096 91232 700160
rect 91296 700096 91312 700160
rect 91376 700096 91404 700160
rect 90804 700095 91404 700096
rect 126804 700160 127404 700161
rect 126804 700096 126832 700160
rect 126896 700096 126912 700160
rect 126976 700096 126992 700160
rect 127056 700096 127072 700160
rect 127136 700096 127152 700160
rect 127216 700096 127232 700160
rect 127296 700096 127312 700160
rect 127376 700096 127404 700160
rect 126804 700095 127404 700096
rect 162804 700160 163404 700161
rect 162804 700096 162832 700160
rect 162896 700096 162912 700160
rect 162976 700096 162992 700160
rect 163056 700096 163072 700160
rect 163136 700096 163152 700160
rect 163216 700096 163232 700160
rect 163296 700096 163312 700160
rect 163376 700096 163404 700160
rect 162804 700095 163404 700096
rect 198804 700160 199404 700161
rect 198804 700096 198832 700160
rect 198896 700096 198912 700160
rect 198976 700096 198992 700160
rect 199056 700096 199072 700160
rect 199136 700096 199152 700160
rect 199216 700096 199232 700160
rect 199296 700096 199312 700160
rect 199376 700096 199404 700160
rect 198804 700095 199404 700096
rect 234804 700160 235404 700161
rect 234804 700096 234832 700160
rect 234896 700096 234912 700160
rect 234976 700096 234992 700160
rect 235056 700096 235072 700160
rect 235136 700096 235152 700160
rect 235216 700096 235232 700160
rect 235296 700096 235312 700160
rect 235376 700096 235404 700160
rect 234804 700095 235404 700096
rect 270804 700160 271404 700161
rect 270804 700096 270832 700160
rect 270896 700096 270912 700160
rect 270976 700096 270992 700160
rect 271056 700096 271072 700160
rect 271136 700096 271152 700160
rect 271216 700096 271232 700160
rect 271296 700096 271312 700160
rect 271376 700096 271404 700160
rect 270804 700095 271404 700096
rect 306804 700160 307404 700161
rect 306804 700096 306832 700160
rect 306896 700096 306912 700160
rect 306976 700096 306992 700160
rect 307056 700096 307072 700160
rect 307136 700096 307152 700160
rect 307216 700096 307232 700160
rect 307296 700096 307312 700160
rect 307376 700096 307404 700160
rect 306804 700095 307404 700096
rect 342804 700160 343404 700161
rect 342804 700096 342832 700160
rect 342896 700096 342912 700160
rect 342976 700096 342992 700160
rect 343056 700096 343072 700160
rect 343136 700096 343152 700160
rect 343216 700096 343232 700160
rect 343296 700096 343312 700160
rect 343376 700096 343404 700160
rect 342804 700095 343404 700096
rect 378804 700160 379404 700161
rect 378804 700096 378832 700160
rect 378896 700096 378912 700160
rect 378976 700096 378992 700160
rect 379056 700096 379072 700160
rect 379136 700096 379152 700160
rect 379216 700096 379232 700160
rect 379296 700096 379312 700160
rect 379376 700096 379404 700160
rect 378804 700095 379404 700096
rect 414804 700160 415404 700161
rect 414804 700096 414832 700160
rect 414896 700096 414912 700160
rect 414976 700096 414992 700160
rect 415056 700096 415072 700160
rect 415136 700096 415152 700160
rect 415216 700096 415232 700160
rect 415296 700096 415312 700160
rect 415376 700096 415404 700160
rect 414804 700095 415404 700096
rect 450804 700160 451404 700161
rect 450804 700096 450832 700160
rect 450896 700096 450912 700160
rect 450976 700096 450992 700160
rect 451056 700096 451072 700160
rect 451136 700096 451152 700160
rect 451216 700096 451232 700160
rect 451296 700096 451312 700160
rect 451376 700096 451404 700160
rect 450804 700095 451404 700096
rect 486804 700160 487404 700161
rect 486804 700096 486832 700160
rect 486896 700096 486912 700160
rect 486976 700096 486992 700160
rect 487056 700096 487072 700160
rect 487136 700096 487152 700160
rect 487216 700096 487232 700160
rect 487296 700096 487312 700160
rect 487376 700096 487404 700160
rect 486804 700095 487404 700096
rect 522804 700160 523404 700161
rect 522804 700096 522832 700160
rect 522896 700096 522912 700160
rect 522976 700096 522992 700160
rect 523056 700096 523072 700160
rect 523136 700096 523152 700160
rect 523216 700096 523232 700160
rect 523296 700096 523312 700160
rect 523376 700096 523404 700160
rect 522804 700095 523404 700096
rect 558804 700160 559404 700161
rect 558804 700096 558832 700160
rect 558896 700096 558912 700160
rect 558976 700096 558992 700160
rect 559056 700096 559072 700160
rect 559136 700096 559152 700160
rect 559216 700096 559232 700160
rect 559296 700096 559312 700160
rect 559376 700096 559404 700160
rect 558804 700095 559404 700096
rect 283097 700090 283163 700093
rect 296621 700090 296687 700093
rect 283097 700088 296687 700090
rect 283097 700032 283102 700088
rect 283158 700032 296626 700088
rect 296682 700032 296687 700088
rect 283097 700030 296687 700032
rect 283097 700027 283163 700030
rect 296621 700027 296687 700030
rect 298001 699954 298067 699957
rect 300117 699954 300183 699957
rect 298001 699952 300183 699954
rect 298001 699896 298006 699952
rect 298062 699896 300122 699952
rect 300178 699896 300183 699952
rect 298001 699894 300183 699896
rect 298001 699891 298067 699894
rect 300117 699891 300183 699894
rect 302325 699954 302391 699957
rect 308581 699954 308647 699957
rect 302325 699952 308647 699954
rect 302325 699896 302330 699952
rect 302386 699896 308586 699952
rect 308642 699896 308647 699952
rect 302325 699894 308647 699896
rect 302325 699891 302391 699894
rect 308581 699891 308647 699894
rect 269062 699756 269068 699820
rect 269132 699818 269138 699820
rect 273897 699818 273963 699821
rect 269132 699816 273963 699818
rect 269132 699760 273902 699816
rect 273958 699760 273963 699816
rect 269132 699758 273963 699760
rect 269132 699756 269138 699758
rect 273897 699755 273963 699758
rect 283741 699818 283807 699821
rect 288709 699818 288775 699821
rect 283741 699816 288775 699818
rect 283741 699760 283746 699816
rect 283802 699760 288714 699816
rect 288770 699760 288775 699816
rect 283741 699758 288775 699760
rect 283741 699755 283807 699758
rect 288709 699755 288775 699758
rect 296713 699818 296779 699821
rect 303613 699818 303679 699821
rect 296713 699816 303679 699818
rect 296713 699760 296718 699816
rect 296774 699760 303618 699816
rect 303674 699760 303679 699816
rect 296713 699758 303679 699760
rect 296713 699755 296779 699758
rect 303613 699755 303679 699758
rect 280061 699682 280127 699685
rect 283005 699682 283071 699685
rect 280061 699680 283071 699682
rect 280061 699624 280066 699680
rect 280122 699624 283010 699680
rect 283066 699624 283071 699680
rect 280061 699622 283071 699624
rect 280061 699619 280127 699622
rect 283005 699619 283071 699622
rect 36804 699616 37404 699617
rect 36804 699552 36832 699616
rect 36896 699552 36912 699616
rect 36976 699552 36992 699616
rect 37056 699552 37072 699616
rect 37136 699552 37152 699616
rect 37216 699552 37232 699616
rect 37296 699552 37312 699616
rect 37376 699552 37404 699616
rect 36804 699551 37404 699552
rect 72804 699616 73404 699617
rect 72804 699552 72832 699616
rect 72896 699552 72912 699616
rect 72976 699552 72992 699616
rect 73056 699552 73072 699616
rect 73136 699552 73152 699616
rect 73216 699552 73232 699616
rect 73296 699552 73312 699616
rect 73376 699552 73404 699616
rect 72804 699551 73404 699552
rect 108804 699616 109404 699617
rect 108804 699552 108832 699616
rect 108896 699552 108912 699616
rect 108976 699552 108992 699616
rect 109056 699552 109072 699616
rect 109136 699552 109152 699616
rect 109216 699552 109232 699616
rect 109296 699552 109312 699616
rect 109376 699552 109404 699616
rect 108804 699551 109404 699552
rect 144804 699616 145404 699617
rect 144804 699552 144832 699616
rect 144896 699552 144912 699616
rect 144976 699552 144992 699616
rect 145056 699552 145072 699616
rect 145136 699552 145152 699616
rect 145216 699552 145232 699616
rect 145296 699552 145312 699616
rect 145376 699552 145404 699616
rect 144804 699551 145404 699552
rect 180804 699616 181404 699617
rect 180804 699552 180832 699616
rect 180896 699552 180912 699616
rect 180976 699552 180992 699616
rect 181056 699552 181072 699616
rect 181136 699552 181152 699616
rect 181216 699552 181232 699616
rect 181296 699552 181312 699616
rect 181376 699552 181404 699616
rect 180804 699551 181404 699552
rect 216804 699616 217404 699617
rect 216804 699552 216832 699616
rect 216896 699552 216912 699616
rect 216976 699552 216992 699616
rect 217056 699552 217072 699616
rect 217136 699552 217152 699616
rect 217216 699552 217232 699616
rect 217296 699552 217312 699616
rect 217376 699552 217404 699616
rect 216804 699551 217404 699552
rect 252804 699616 253404 699617
rect 252804 699552 252832 699616
rect 252896 699552 252912 699616
rect 252976 699552 252992 699616
rect 253056 699552 253072 699616
rect 253136 699552 253152 699616
rect 253216 699552 253232 699616
rect 253296 699552 253312 699616
rect 253376 699552 253404 699616
rect 252804 699551 253404 699552
rect 288804 699616 289404 699617
rect 288804 699552 288832 699616
rect 288896 699552 288912 699616
rect 288976 699552 288992 699616
rect 289056 699552 289072 699616
rect 289136 699552 289152 699616
rect 289216 699552 289232 699616
rect 289296 699552 289312 699616
rect 289376 699552 289404 699616
rect 288804 699551 289404 699552
rect 324804 699616 325404 699617
rect 324804 699552 324832 699616
rect 324896 699552 324912 699616
rect 324976 699552 324992 699616
rect 325056 699552 325072 699616
rect 325136 699552 325152 699616
rect 325216 699552 325232 699616
rect 325296 699552 325312 699616
rect 325376 699552 325404 699616
rect 324804 699551 325404 699552
rect 360804 699616 361404 699617
rect 360804 699552 360832 699616
rect 360896 699552 360912 699616
rect 360976 699552 360992 699616
rect 361056 699552 361072 699616
rect 361136 699552 361152 699616
rect 361216 699552 361232 699616
rect 361296 699552 361312 699616
rect 361376 699552 361404 699616
rect 360804 699551 361404 699552
rect 396804 699616 397404 699617
rect 396804 699552 396832 699616
rect 396896 699552 396912 699616
rect 396976 699552 396992 699616
rect 397056 699552 397072 699616
rect 397136 699552 397152 699616
rect 397216 699552 397232 699616
rect 397296 699552 397312 699616
rect 397376 699552 397404 699616
rect 396804 699551 397404 699552
rect 432804 699616 433404 699617
rect 432804 699552 432832 699616
rect 432896 699552 432912 699616
rect 432976 699552 432992 699616
rect 433056 699552 433072 699616
rect 433136 699552 433152 699616
rect 433216 699552 433232 699616
rect 433296 699552 433312 699616
rect 433376 699552 433404 699616
rect 432804 699551 433404 699552
rect 468804 699616 469404 699617
rect 468804 699552 468832 699616
rect 468896 699552 468912 699616
rect 468976 699552 468992 699616
rect 469056 699552 469072 699616
rect 469136 699552 469152 699616
rect 469216 699552 469232 699616
rect 469296 699552 469312 699616
rect 469376 699552 469404 699616
rect 468804 699551 469404 699552
rect 504804 699616 505404 699617
rect 504804 699552 504832 699616
rect 504896 699552 504912 699616
rect 504976 699552 504992 699616
rect 505056 699552 505072 699616
rect 505136 699552 505152 699616
rect 505216 699552 505232 699616
rect 505296 699552 505312 699616
rect 505376 699552 505404 699616
rect 504804 699551 505404 699552
rect 540804 699616 541404 699617
rect 540804 699552 540832 699616
rect 540896 699552 540912 699616
rect 540976 699552 540992 699616
rect 541056 699552 541072 699616
rect 541136 699552 541152 699616
rect 541216 699552 541232 699616
rect 541296 699552 541312 699616
rect 541376 699552 541404 699616
rect 540804 699551 541404 699552
rect 576804 699616 577404 699617
rect 576804 699552 576832 699616
rect 576896 699552 576912 699616
rect 576976 699552 576992 699616
rect 577056 699552 577072 699616
rect 577136 699552 577152 699616
rect 577216 699552 577232 699616
rect 577296 699552 577312 699616
rect 577376 699552 577404 699616
rect 576804 699551 577404 699552
rect 259453 699546 259519 699549
rect 269062 699546 269068 699548
rect 259453 699544 269068 699546
rect 259453 699488 259458 699544
rect 259514 699488 269068 699544
rect 259453 699486 269068 699488
rect 259453 699483 259519 699486
rect 269062 699484 269068 699486
rect 269132 699484 269138 699548
rect 289721 699546 289787 699549
rect 296897 699546 296963 699549
rect 289721 699544 296963 699546
rect 289721 699488 289726 699544
rect 289782 699488 296902 699544
rect 296958 699488 296963 699544
rect 289721 699486 296963 699488
rect 289721 699483 289787 699486
rect 296897 699483 296963 699486
rect 273253 699410 273319 699413
rect 283005 699410 283071 699413
rect 273253 699408 283071 699410
rect 273253 699352 273258 699408
rect 273314 699352 283010 699408
rect 283066 699352 283071 699408
rect 273253 699350 283071 699352
rect 273253 699347 273319 699350
rect 283005 699347 283071 699350
rect 292389 699410 292455 699413
rect 294045 699410 294111 699413
rect 292389 699408 294111 699410
rect 292389 699352 292394 699408
rect 292450 699352 294050 699408
rect 294106 699352 294111 699408
rect 292389 699350 294111 699352
rect 292389 699347 292455 699350
rect 294045 699347 294111 699350
rect 186129 699274 186195 699277
rect 244089 699274 244155 699277
rect 186129 699272 244155 699274
rect 186129 699216 186134 699272
rect 186190 699216 244094 699272
rect 244150 699216 244155 699272
rect 186129 699214 244155 699216
rect 186129 699211 186195 699214
rect 244089 699211 244155 699214
rect 244273 699274 244339 699277
rect 267641 699274 267707 699277
rect 273345 699274 273411 699277
rect 244273 699272 267707 699274
rect 244273 699216 244278 699272
rect 244334 699216 267646 699272
rect 267702 699216 267707 699272
rect 244273 699214 267707 699216
rect 244273 699211 244339 699214
rect 267641 699211 267707 699214
rect 269070 699272 273411 699274
rect 269070 699216 273350 699272
rect 273406 699216 273411 699272
rect 269070 699214 273411 699216
rect 18804 699072 19404 699073
rect 18804 699008 18832 699072
rect 18896 699008 18912 699072
rect 18976 699008 18992 699072
rect 19056 699008 19072 699072
rect 19136 699008 19152 699072
rect 19216 699008 19232 699072
rect 19296 699008 19312 699072
rect 19376 699008 19404 699072
rect 18804 699007 19404 699008
rect 54804 699072 55404 699073
rect 54804 699008 54832 699072
rect 54896 699008 54912 699072
rect 54976 699008 54992 699072
rect 55056 699008 55072 699072
rect 55136 699008 55152 699072
rect 55216 699008 55232 699072
rect 55296 699008 55312 699072
rect 55376 699008 55404 699072
rect 54804 699007 55404 699008
rect 90804 699072 91404 699073
rect 90804 699008 90832 699072
rect 90896 699008 90912 699072
rect 90976 699008 90992 699072
rect 91056 699008 91072 699072
rect 91136 699008 91152 699072
rect 91216 699008 91232 699072
rect 91296 699008 91312 699072
rect 91376 699008 91404 699072
rect 90804 699007 91404 699008
rect 126804 699072 127404 699073
rect 126804 699008 126832 699072
rect 126896 699008 126912 699072
rect 126976 699008 126992 699072
rect 127056 699008 127072 699072
rect 127136 699008 127152 699072
rect 127216 699008 127232 699072
rect 127296 699008 127312 699072
rect 127376 699008 127404 699072
rect 126804 699007 127404 699008
rect 162804 699072 163404 699073
rect 162804 699008 162832 699072
rect 162896 699008 162912 699072
rect 162976 699008 162992 699072
rect 163056 699008 163072 699072
rect 163136 699008 163152 699072
rect 163216 699008 163232 699072
rect 163296 699008 163312 699072
rect 163376 699008 163404 699072
rect 162804 699007 163404 699008
rect 198804 699072 199404 699073
rect 198804 699008 198832 699072
rect 198896 699008 198912 699072
rect 198976 699008 198992 699072
rect 199056 699008 199072 699072
rect 199136 699008 199152 699072
rect 199216 699008 199232 699072
rect 199296 699008 199312 699072
rect 199376 699008 199404 699072
rect 198804 699007 199404 699008
rect 234804 699072 235404 699073
rect 234804 699008 234832 699072
rect 234896 699008 234912 699072
rect 234976 699008 234992 699072
rect 235056 699008 235072 699072
rect 235136 699008 235152 699072
rect 235216 699008 235232 699072
rect 235296 699008 235312 699072
rect 235376 699008 235404 699072
rect 234804 699007 235404 699008
rect 244089 699002 244155 699005
rect 244365 699002 244431 699005
rect 244089 699000 244431 699002
rect 244089 698944 244094 699000
rect 244150 698944 244370 699000
rect 244426 698944 244431 699000
rect 244089 698942 244431 698944
rect 244089 698939 244155 698942
rect 244365 698939 244431 698942
rect 253749 699002 253815 699005
rect 269070 699002 269130 699214
rect 273345 699211 273411 699214
rect 277393 699274 277459 699277
rect 292481 699274 292547 699277
rect 277393 699272 292547 699274
rect 277393 699216 277398 699272
rect 277454 699216 292486 699272
rect 292542 699216 292547 699272
rect 277393 699214 292547 699216
rect 277393 699211 277459 699214
rect 292481 699211 292547 699214
rect 296529 699274 296595 699277
rect 302325 699274 302391 699277
rect 296529 699272 302391 699274
rect 296529 699216 296534 699272
rect 296590 699216 302330 699272
rect 302386 699216 302391 699272
rect 296529 699214 302391 699216
rect 296529 699211 296595 699214
rect 302325 699211 302391 699214
rect 311985 699274 312051 699277
rect 321645 699274 321711 699277
rect 311985 699272 321711 699274
rect 311985 699216 311990 699272
rect 312046 699216 321650 699272
rect 321706 699216 321711 699272
rect 311985 699214 321711 699216
rect 311985 699211 312051 699214
rect 321645 699211 321711 699214
rect 331029 699274 331095 699277
rect 331305 699274 331371 699277
rect 331029 699272 331371 699274
rect 331029 699216 331034 699272
rect 331090 699216 331310 699272
rect 331366 699216 331371 699272
rect 331029 699214 331371 699216
rect 331029 699211 331095 699214
rect 331305 699211 331371 699214
rect 340689 699274 340755 699277
rect 344921 699274 344987 699277
rect 340689 699272 344987 699274
rect 340689 699216 340694 699272
rect 340750 699216 344926 699272
rect 344982 699216 344987 699272
rect 340689 699214 344987 699216
rect 340689 699211 340755 699214
rect 344921 699211 344987 699214
rect 364333 699274 364399 699277
rect 373901 699274 373967 699277
rect 364333 699272 373967 699274
rect 364333 699216 364338 699272
rect 364394 699216 373906 699272
rect 373962 699216 373967 699272
rect 364333 699214 373967 699216
rect 364333 699211 364399 699214
rect 373901 699211 373967 699214
rect 374085 699274 374151 699277
rect 383561 699274 383627 699277
rect 374085 699272 383627 699274
rect 374085 699216 374090 699272
rect 374146 699216 383566 699272
rect 383622 699216 383627 699272
rect 374085 699214 383627 699216
rect 374085 699211 374151 699214
rect 383561 699211 383627 699214
rect 503478 699212 503484 699276
rect 503548 699274 503554 699276
rect 526253 699274 526319 699277
rect 503548 699272 526319 699274
rect 503548 699216 526258 699272
rect 526314 699216 526319 699272
rect 503548 699214 526319 699216
rect 503548 699212 503554 699214
rect 526253 699211 526319 699214
rect 282913 699138 282979 699141
rect 296621 699138 296687 699141
rect 282913 699136 296687 699138
rect 282913 699080 282918 699136
rect 282974 699080 296626 699136
rect 296682 699080 296687 699136
rect 282913 699078 296687 699080
rect 282913 699075 282979 699078
rect 296621 699075 296687 699078
rect 321553 699138 321619 699141
rect 331121 699138 331187 699141
rect 321553 699136 331187 699138
rect 321553 699080 321558 699136
rect 321614 699080 331126 699136
rect 331182 699080 331187 699136
rect 321553 699078 331187 699080
rect 321553 699075 321619 699078
rect 331121 699075 331187 699078
rect 270804 699072 271404 699073
rect 270804 699008 270832 699072
rect 270896 699008 270912 699072
rect 270976 699008 270992 699072
rect 271056 699008 271072 699072
rect 271136 699008 271152 699072
rect 271216 699008 271232 699072
rect 271296 699008 271312 699072
rect 271376 699008 271404 699072
rect 270804 699007 271404 699008
rect 306804 699072 307404 699073
rect 306804 699008 306832 699072
rect 306896 699008 306912 699072
rect 306976 699008 306992 699072
rect 307056 699008 307072 699072
rect 307136 699008 307152 699072
rect 307216 699008 307232 699072
rect 307296 699008 307312 699072
rect 307376 699008 307404 699072
rect 306804 699007 307404 699008
rect 342804 699072 343404 699073
rect 342804 699008 342832 699072
rect 342896 699008 342912 699072
rect 342976 699008 342992 699072
rect 343056 699008 343072 699072
rect 343136 699008 343152 699072
rect 343216 699008 343232 699072
rect 343296 699008 343312 699072
rect 343376 699008 343404 699072
rect 342804 699007 343404 699008
rect 378804 699072 379404 699073
rect 378804 699008 378832 699072
rect 378896 699008 378912 699072
rect 378976 699008 378992 699072
rect 379056 699008 379072 699072
rect 379136 699008 379152 699072
rect 379216 699008 379232 699072
rect 379296 699008 379312 699072
rect 379376 699008 379404 699072
rect 378804 699007 379404 699008
rect 414804 699072 415404 699073
rect 414804 699008 414832 699072
rect 414896 699008 414912 699072
rect 414976 699008 414992 699072
rect 415056 699008 415072 699072
rect 415136 699008 415152 699072
rect 415216 699008 415232 699072
rect 415296 699008 415312 699072
rect 415376 699008 415404 699072
rect 414804 699007 415404 699008
rect 450804 699072 451404 699073
rect 450804 699008 450832 699072
rect 450896 699008 450912 699072
rect 450976 699008 450992 699072
rect 451056 699008 451072 699072
rect 451136 699008 451152 699072
rect 451216 699008 451232 699072
rect 451296 699008 451312 699072
rect 451376 699008 451404 699072
rect 450804 699007 451404 699008
rect 486804 699072 487404 699073
rect 486804 699008 486832 699072
rect 486896 699008 486912 699072
rect 486976 699008 486992 699072
rect 487056 699008 487072 699072
rect 487136 699008 487152 699072
rect 487216 699008 487232 699072
rect 487296 699008 487312 699072
rect 487376 699008 487404 699072
rect 486804 699007 487404 699008
rect 522804 699072 523404 699073
rect 522804 699008 522832 699072
rect 522896 699008 522912 699072
rect 522976 699008 522992 699072
rect 523056 699008 523072 699072
rect 523136 699008 523152 699072
rect 523216 699008 523232 699072
rect 523296 699008 523312 699072
rect 523376 699008 523404 699072
rect 522804 699007 523404 699008
rect 558804 699072 559404 699073
rect 558804 699008 558832 699072
rect 558896 699008 558912 699072
rect 558976 699008 558992 699072
rect 559056 699008 559072 699072
rect 559136 699008 559152 699072
rect 559216 699008 559232 699072
rect 559296 699008 559312 699072
rect 559376 699008 559404 699072
rect 558804 699007 559404 699008
rect 253749 699000 269130 699002
rect 253749 698944 253754 699000
rect 253810 698944 269130 699000
rect 253749 698942 269130 698944
rect 311985 699002 312051 699005
rect 321645 699002 321711 699005
rect 311985 699000 321711 699002
rect 311985 698944 311990 699000
rect 312046 698944 321650 699000
rect 321706 698944 321711 699000
rect 311985 698942 321711 698944
rect 253749 698939 253815 698942
rect 311985 698939 312051 698942
rect 321645 698939 321711 698942
rect 4797 698866 4863 698869
rect 545113 698866 545179 698869
rect 4797 698864 545179 698866
rect 4797 698808 4802 698864
rect 4858 698808 545118 698864
rect 545174 698808 545179 698864
rect 4797 698806 545179 698808
rect 4797 698803 4863 698806
rect 545113 698803 545179 698806
rect 4981 698730 5047 698733
rect 516777 698730 516843 698733
rect 4981 698728 516843 698730
rect 4981 698672 4986 698728
rect 5042 698672 516782 698728
rect 516838 698672 516843 698728
rect 4981 698670 516843 698672
rect 4981 698667 5047 698670
rect 516777 698667 516843 698670
rect 36804 698528 37404 698529
rect 36804 698464 36832 698528
rect 36896 698464 36912 698528
rect 36976 698464 36992 698528
rect 37056 698464 37072 698528
rect 37136 698464 37152 698528
rect 37216 698464 37232 698528
rect 37296 698464 37312 698528
rect 37376 698464 37404 698528
rect 36804 698463 37404 698464
rect 72804 698528 73404 698529
rect 72804 698464 72832 698528
rect 72896 698464 72912 698528
rect 72976 698464 72992 698528
rect 73056 698464 73072 698528
rect 73136 698464 73152 698528
rect 73216 698464 73232 698528
rect 73296 698464 73312 698528
rect 73376 698464 73404 698528
rect 72804 698463 73404 698464
rect 108804 698528 109404 698529
rect 108804 698464 108832 698528
rect 108896 698464 108912 698528
rect 108976 698464 108992 698528
rect 109056 698464 109072 698528
rect 109136 698464 109152 698528
rect 109216 698464 109232 698528
rect 109296 698464 109312 698528
rect 109376 698464 109404 698528
rect 108804 698463 109404 698464
rect 144804 698528 145404 698529
rect 144804 698464 144832 698528
rect 144896 698464 144912 698528
rect 144976 698464 144992 698528
rect 145056 698464 145072 698528
rect 145136 698464 145152 698528
rect 145216 698464 145232 698528
rect 145296 698464 145312 698528
rect 145376 698464 145404 698528
rect 144804 698463 145404 698464
rect 180804 698528 181404 698529
rect 180804 698464 180832 698528
rect 180896 698464 180912 698528
rect 180976 698464 180992 698528
rect 181056 698464 181072 698528
rect 181136 698464 181152 698528
rect 181216 698464 181232 698528
rect 181296 698464 181312 698528
rect 181376 698464 181404 698528
rect 180804 698463 181404 698464
rect 216804 698528 217404 698529
rect 216804 698464 216832 698528
rect 216896 698464 216912 698528
rect 216976 698464 216992 698528
rect 217056 698464 217072 698528
rect 217136 698464 217152 698528
rect 217216 698464 217232 698528
rect 217296 698464 217312 698528
rect 217376 698464 217404 698528
rect 216804 698463 217404 698464
rect 252804 698528 253404 698529
rect 252804 698464 252832 698528
rect 252896 698464 252912 698528
rect 252976 698464 252992 698528
rect 253056 698464 253072 698528
rect 253136 698464 253152 698528
rect 253216 698464 253232 698528
rect 253296 698464 253312 698528
rect 253376 698464 253404 698528
rect 252804 698463 253404 698464
rect 288804 698528 289404 698529
rect 288804 698464 288832 698528
rect 288896 698464 288912 698528
rect 288976 698464 288992 698528
rect 289056 698464 289072 698528
rect 289136 698464 289152 698528
rect 289216 698464 289232 698528
rect 289296 698464 289312 698528
rect 289376 698464 289404 698528
rect 288804 698463 289404 698464
rect 324804 698528 325404 698529
rect 324804 698464 324832 698528
rect 324896 698464 324912 698528
rect 324976 698464 324992 698528
rect 325056 698464 325072 698528
rect 325136 698464 325152 698528
rect 325216 698464 325232 698528
rect 325296 698464 325312 698528
rect 325376 698464 325404 698528
rect 324804 698463 325404 698464
rect 360804 698528 361404 698529
rect 360804 698464 360832 698528
rect 360896 698464 360912 698528
rect 360976 698464 360992 698528
rect 361056 698464 361072 698528
rect 361136 698464 361152 698528
rect 361216 698464 361232 698528
rect 361296 698464 361312 698528
rect 361376 698464 361404 698528
rect 360804 698463 361404 698464
rect 396804 698528 397404 698529
rect 396804 698464 396832 698528
rect 396896 698464 396912 698528
rect 396976 698464 396992 698528
rect 397056 698464 397072 698528
rect 397136 698464 397152 698528
rect 397216 698464 397232 698528
rect 397296 698464 397312 698528
rect 397376 698464 397404 698528
rect 396804 698463 397404 698464
rect 432804 698528 433404 698529
rect 432804 698464 432832 698528
rect 432896 698464 432912 698528
rect 432976 698464 432992 698528
rect 433056 698464 433072 698528
rect 433136 698464 433152 698528
rect 433216 698464 433232 698528
rect 433296 698464 433312 698528
rect 433376 698464 433404 698528
rect 432804 698463 433404 698464
rect 468804 698528 469404 698529
rect 468804 698464 468832 698528
rect 468896 698464 468912 698528
rect 468976 698464 468992 698528
rect 469056 698464 469072 698528
rect 469136 698464 469152 698528
rect 469216 698464 469232 698528
rect 469296 698464 469312 698528
rect 469376 698464 469404 698528
rect 468804 698463 469404 698464
rect 504804 698528 505404 698529
rect 504804 698464 504832 698528
rect 504896 698464 504912 698528
rect 504976 698464 504992 698528
rect 505056 698464 505072 698528
rect 505136 698464 505152 698528
rect 505216 698464 505232 698528
rect 505296 698464 505312 698528
rect 505376 698464 505404 698528
rect 504804 698463 505404 698464
rect 540804 698528 541404 698529
rect 540804 698464 540832 698528
rect 540896 698464 540912 698528
rect 540976 698464 540992 698528
rect 541056 698464 541072 698528
rect 541136 698464 541152 698528
rect 541216 698464 541232 698528
rect 541296 698464 541312 698528
rect 541376 698464 541404 698528
rect 540804 698463 541404 698464
rect 576804 698528 577404 698529
rect 576804 698464 576832 698528
rect 576896 698464 576912 698528
rect 576976 698464 576992 698528
rect 577056 698464 577072 698528
rect 577136 698464 577152 698528
rect 577216 698464 577232 698528
rect 577296 698464 577312 698528
rect 577376 698464 577404 698528
rect 576804 698463 577404 698464
rect 218053 698458 218119 698461
rect 218421 698458 218487 698461
rect 218053 698456 218487 698458
rect 218053 698400 218058 698456
rect 218114 698400 218426 698456
rect 218482 698400 218487 698456
rect 218053 698398 218487 698400
rect 218053 698395 218119 698398
rect 218421 698395 218487 698398
rect 218053 698322 218119 698325
rect 218421 698322 218487 698325
rect 218053 698320 218487 698322
rect 218053 698264 218058 698320
rect 218114 698264 218426 698320
rect 218482 698264 218487 698320
rect 218053 698262 218487 698264
rect 218053 698259 218119 698262
rect 218421 698259 218487 698262
rect 226333 698322 226399 698325
rect 235901 698322 235967 698325
rect 226333 698320 235967 698322
rect 226333 698264 226338 698320
rect 226394 698264 235906 698320
rect 235962 698264 235967 698320
rect 226333 698262 235967 698264
rect 226333 698259 226399 698262
rect 235901 698259 235967 698262
rect 248321 698322 248387 698325
rect 253841 698322 253907 698325
rect 248321 698320 253907 698322
rect 248321 698264 248326 698320
rect 248382 698264 253846 698320
rect 253902 698264 253907 698320
rect 248321 698262 253907 698264
rect 248321 698259 248387 698262
rect 253841 698259 253907 698262
rect 208945 698186 209011 698189
rect 215109 698186 215175 698189
rect 208945 698184 215175 698186
rect 208945 698128 208950 698184
rect 209006 698128 215114 698184
rect 215170 698128 215175 698184
rect 208945 698126 215175 698128
rect 208945 698123 209011 698126
rect 215109 698123 215175 698126
rect 237373 698186 237439 698189
rect 237557 698186 237623 698189
rect 237373 698184 237623 698186
rect 237373 698128 237378 698184
rect 237434 698128 237562 698184
rect 237618 698128 237623 698184
rect 237373 698126 237623 698128
rect 237373 698123 237439 698126
rect 237557 698123 237623 698126
rect 253841 698186 253907 698189
rect 254025 698186 254091 698189
rect 253841 698184 254091 698186
rect 253841 698128 253846 698184
rect 253902 698128 254030 698184
rect 254086 698128 254091 698184
rect 253841 698126 254091 698128
rect 253841 698123 253907 698126
rect 254025 698123 254091 698126
rect 275737 698186 275803 698189
rect 277393 698186 277459 698189
rect 275737 698184 277459 698186
rect 275737 698128 275742 698184
rect 275798 698128 277398 698184
rect 277454 698128 277459 698184
rect 275737 698126 277459 698128
rect 275737 698123 275803 698126
rect 277393 698123 277459 698126
rect 350441 698186 350507 698189
rect 350717 698186 350783 698189
rect 350441 698184 350783 698186
rect 350441 698128 350446 698184
rect 350502 698128 350722 698184
rect 350778 698128 350783 698184
rect 350441 698126 350783 698128
rect 350441 698123 350507 698126
rect 350717 698123 350783 698126
rect 193305 698050 193371 698053
rect 202781 698050 202847 698053
rect 193305 698048 202847 698050
rect 193305 697992 193310 698048
rect 193366 697992 202786 698048
rect 202842 697992 202847 698048
rect 193305 697990 202847 697992
rect 193305 697987 193371 697990
rect 202781 697987 202847 697990
rect 579613 698050 579679 698053
rect 583520 698050 584960 698140
rect 579613 698048 584960 698050
rect 579613 697992 579618 698048
rect 579674 697992 584960 698048
rect 579613 697990 584960 697992
rect 579613 697987 579679 697990
rect 583520 697900 584960 697990
rect 6177 697098 6243 697101
rect 540421 697098 540487 697101
rect 6177 697096 540487 697098
rect 6177 697040 6182 697096
rect 6238 697040 540426 697096
rect 540482 697040 540487 697096
rect 6177 697038 540487 697040
rect 6177 697035 6243 697038
rect 540421 697035 540487 697038
rect 10317 696962 10383 696965
rect 574737 696962 574803 696965
rect 10317 696960 574803 696962
rect 10317 696904 10322 696960
rect 10378 696904 574742 696960
rect 574798 696904 574803 696960
rect 10317 696902 574803 696904
rect 10317 696899 10383 696902
rect 574737 696899 574803 696902
rect 232957 696826 233023 696829
rect 234521 696826 234587 696829
rect 232957 696824 234587 696826
rect -960 696540 480 696780
rect 232957 696768 232962 696824
rect 233018 696768 234526 696824
rect 234582 696768 234587 696824
rect 232957 696766 234587 696768
rect 232957 696763 233023 696766
rect 234521 696763 234587 696766
rect 244273 696826 244339 696829
rect 248413 696826 248479 696829
rect 244273 696824 248479 696826
rect 244273 696768 244278 696824
rect 244334 696768 248418 696824
rect 248474 696768 248479 696824
rect 244273 696766 248479 696768
rect 244273 696763 244339 696766
rect 248413 696763 248479 696766
rect 309133 696826 309199 696829
rect 318609 696826 318675 696829
rect 309133 696824 318675 696826
rect 309133 696768 309138 696824
rect 309194 696768 318614 696824
rect 318670 696768 318675 696824
rect 309133 696766 318675 696768
rect 309133 696763 309199 696766
rect 318609 696763 318675 696766
rect 338113 696826 338179 696829
rect 342621 696826 342687 696829
rect 338113 696824 342687 696826
rect 338113 696768 338118 696824
rect 338174 696768 342626 696824
rect 342682 696768 342687 696824
rect 338113 696766 342687 696768
rect 338113 696763 338179 696766
rect 342621 696763 342687 696766
rect 299473 696690 299539 696693
rect 309041 696690 309107 696693
rect 299473 696688 309107 696690
rect 299473 696632 299478 696688
rect 299534 696632 309046 696688
rect 309102 696632 309107 696688
rect 299473 696630 309107 696632
rect 299473 696627 299539 696630
rect 309041 696627 309107 696630
rect 318793 696690 318859 696693
rect 321553 696690 321619 696693
rect 318793 696688 321619 696690
rect 318793 696632 318798 696688
rect 318854 696632 321558 696688
rect 321614 696632 321619 696688
rect 318793 696630 321619 696632
rect 318793 696627 318859 696630
rect 321553 696627 321619 696630
rect 328453 696690 328519 696693
rect 338021 696690 338087 696693
rect 328453 696688 338087 696690
rect 328453 696632 328458 696688
rect 328514 696632 338026 696688
rect 338082 696632 338087 696688
rect 328453 696630 338087 696632
rect 328453 696627 328519 696630
rect 338021 696627 338087 696630
rect 224953 696418 225019 696421
rect 234521 696418 234587 696421
rect 224953 696416 234587 696418
rect 224953 696360 224958 696416
rect 225014 696360 234526 696416
rect 234582 696360 234587 696416
rect 224953 696358 234587 696360
rect 224953 696355 225019 696358
rect 234521 696355 234587 696358
rect 244273 696418 244339 696421
rect 253841 696418 253907 696421
rect 244273 696416 253907 696418
rect 244273 696360 244278 696416
rect 244334 696360 253846 696416
rect 253902 696360 253907 696416
rect 244273 696358 253907 696360
rect 244273 696355 244339 696358
rect 253841 696355 253907 696358
rect 263593 696418 263659 696421
rect 273161 696418 273227 696421
rect 263593 696416 273227 696418
rect 263593 696360 263598 696416
rect 263654 696360 273166 696416
rect 273222 696360 273227 696416
rect 263593 696358 273227 696360
rect 263593 696355 263659 696358
rect 273161 696355 273227 696358
rect 282913 696418 282979 696421
rect 292481 696418 292547 696421
rect 282913 696416 292547 696418
rect 282913 696360 282918 696416
rect 282974 696360 292486 696416
rect 292542 696360 292547 696416
rect 282913 696358 292547 696360
rect 282913 696355 282979 696358
rect 292481 696355 292547 696358
rect 89713 696146 89779 696149
rect 580257 696146 580323 696149
rect 89713 696144 580323 696146
rect 89713 696088 89718 696144
rect 89774 696088 580262 696144
rect 580318 696088 580323 696144
rect 89713 696086 580323 696088
rect 89713 696083 89779 696086
rect 580257 696083 580323 696086
rect 19977 696010 20043 696013
rect 205541 696010 205607 696013
rect 213729 696010 213795 696013
rect 19977 696008 29010 696010
rect 19977 695952 19982 696008
rect 20038 695952 29010 696008
rect 19977 695950 29010 695952
rect 19977 695947 20043 695950
rect 28950 695874 29010 695950
rect 205541 696008 213795 696010
rect 205541 695952 205546 696008
rect 205602 695952 213734 696008
rect 213790 695952 213795 696008
rect 205541 695950 213795 695952
rect 205541 695947 205607 695950
rect 213729 695947 213795 695950
rect 229001 696010 229067 696013
rect 230381 696010 230447 696013
rect 229001 696008 230447 696010
rect 229001 695952 229006 696008
rect 229062 695952 230386 696008
rect 230442 695952 230447 696008
rect 229001 695950 230447 695952
rect 229001 695947 229067 695950
rect 230381 695947 230447 695950
rect 241462 695948 241468 696012
rect 241532 696010 241538 696012
rect 251081 696010 251147 696013
rect 241532 696008 251147 696010
rect 241532 695952 251086 696008
rect 251142 695952 251147 696008
rect 241532 695950 251147 695952
rect 241532 695948 241538 695950
rect 251081 695947 251147 695950
rect 260782 695948 260788 696012
rect 260852 696010 260858 696012
rect 265617 696010 265683 696013
rect 260852 696008 265683 696010
rect 260852 695952 265622 696008
rect 265678 695952 265683 696008
rect 260852 695950 265683 695952
rect 260852 695948 260858 695950
rect 265617 695947 265683 695950
rect 318742 695948 318748 696012
rect 318812 696010 318818 696012
rect 328361 696010 328427 696013
rect 371877 696010 371943 696013
rect 468477 696010 468543 696013
rect 318812 696008 328427 696010
rect 318812 695952 328366 696008
rect 328422 695952 328427 696008
rect 318812 695950 328427 695952
rect 318812 695948 318818 695950
rect 328361 695947 328427 695950
rect 367142 696008 371943 696010
rect 367142 695952 371882 696008
rect 371938 695952 371943 696008
rect 367142 695950 371943 695952
rect 28950 695814 29194 695874
rect 29134 695738 29194 695814
rect 144862 695812 144868 695876
rect 144932 695874 144938 695876
rect 292665 695874 292731 695877
rect 299381 695874 299447 695877
rect 367142 695876 367202 695950
rect 371877 695947 371943 695950
rect 463742 696008 468543 696010
rect 463742 695952 468482 696008
rect 468538 695952 468543 696008
rect 463742 695950 468543 695952
rect 347630 695874 347636 695876
rect 144932 695814 181546 695874
rect 144932 695812 144938 695814
rect 119981 695738 120047 695741
rect 29134 695736 120047 695738
rect 29134 695680 119986 695736
rect 120042 695680 120047 695736
rect 29134 695678 120047 695680
rect 119981 695675 120047 695678
rect 120165 695602 120231 695605
rect 144862 695602 144868 695604
rect 120165 695600 144868 695602
rect 120165 695544 120170 695600
rect 120226 695544 144868 695600
rect 120165 695542 144868 695544
rect 120165 695539 120231 695542
rect 144862 695540 144868 695542
rect 144932 695540 144938 695604
rect 176193 695602 176259 695605
rect 176510 695602 176516 695604
rect 176193 695600 176516 695602
rect 176193 695544 176198 695600
rect 176254 695544 176516 695600
rect 176193 695542 176516 695544
rect 176193 695539 176259 695542
rect 176510 695540 176516 695542
rect 176580 695540 176586 695604
rect 181486 695602 181546 695814
rect 270542 695814 280124 695874
rect 234613 695738 234679 695741
rect 241462 695738 241468 695740
rect 234613 695736 241468 695738
rect 234613 695680 234618 695736
rect 234674 695680 241468 695736
rect 234613 695678 241468 695680
rect 234613 695675 234679 695678
rect 241462 695676 241468 695678
rect 241532 695676 241538 695740
rect 253933 695738 253999 695741
rect 260782 695738 260788 695740
rect 253933 695736 260788 695738
rect 253933 695680 253938 695736
rect 253994 695680 260788 695736
rect 253933 695678 260788 695680
rect 253933 695675 253999 695678
rect 260782 695676 260788 695678
rect 260852 695676 260858 695740
rect 265617 695738 265683 695741
rect 270542 695738 270602 695814
rect 265617 695736 270602 695738
rect 265617 695680 265622 695736
rect 265678 695680 270602 695736
rect 265617 695678 270602 695680
rect 280064 695738 280124 695814
rect 292665 695872 299447 695874
rect 292665 695816 292670 695872
rect 292726 695816 299386 695872
rect 299442 695816 299447 695872
rect 292665 695814 299447 695816
rect 292665 695811 292731 695814
rect 299381 695811 299447 695814
rect 340692 695814 347636 695874
rect 292481 695738 292547 695741
rect 280064 695736 292547 695738
rect 280064 695680 292486 695736
rect 292542 695680 292547 695736
rect 280064 695678 292547 695680
rect 265617 695675 265683 695678
rect 292481 695675 292547 695678
rect 309225 695738 309291 695741
rect 318742 695738 318748 695740
rect 309225 695736 318748 695738
rect 309225 695680 309230 695736
rect 309286 695680 318748 695736
rect 309225 695678 318748 695680
rect 309225 695675 309291 695678
rect 318742 695676 318748 695678
rect 318812 695676 318818 695740
rect 331213 695738 331279 695741
rect 340692 695738 340752 695814
rect 347630 695812 347636 695814
rect 347700 695812 347706 695876
rect 367134 695812 367140 695876
rect 367204 695812 367210 695876
rect 422201 695874 422267 695877
rect 425053 695874 425119 695877
rect 422201 695872 425119 695874
rect 422201 695816 422206 695872
rect 422262 695816 425058 695872
rect 425114 695816 425119 695872
rect 422201 695814 425119 695816
rect 422201 695811 422267 695814
rect 425053 695811 425119 695814
rect 434662 695812 434668 695876
rect 434732 695874 434738 695876
rect 437289 695874 437355 695877
rect 434732 695872 437355 695874
rect 434732 695816 437294 695872
rect 437350 695816 437355 695872
rect 434732 695814 437355 695816
rect 434732 695812 434738 695814
rect 437289 695811 437355 695814
rect 437473 695874 437539 695877
rect 463742 695876 463802 695950
rect 468477 695947 468543 695950
rect 473302 695948 473308 696012
rect 473372 696010 473378 696012
rect 482921 696010 482987 696013
rect 473372 696008 482987 696010
rect 473372 695952 482926 696008
rect 482982 695952 482987 696008
rect 473372 695950 482987 695952
rect 473372 695948 473378 695950
rect 482921 695947 482987 695950
rect 442942 695874 442948 695876
rect 437473 695872 442948 695874
rect 437473 695816 437478 695872
rect 437534 695816 442948 695872
rect 437473 695814 442948 695816
rect 437473 695811 437539 695814
rect 442942 695812 442948 695814
rect 443012 695812 443018 695876
rect 463734 695812 463740 695876
rect 463804 695812 463810 695876
rect 495390 695814 505202 695874
rect 331213 695736 340752 695738
rect 331213 695680 331218 695736
rect 331274 695680 340752 695736
rect 331213 695678 340752 695680
rect 360285 695738 360351 695741
rect 367134 695738 367140 695740
rect 360285 695736 367140 695738
rect 360285 695680 360290 695736
rect 360346 695680 367140 695736
rect 360285 695678 367140 695680
rect 331213 695675 331279 695678
rect 360285 695675 360351 695678
rect 367134 695676 367140 695678
rect 367204 695676 367210 695740
rect 384941 695738 385007 695741
rect 386597 695738 386663 695741
rect 398741 695738 398807 695741
rect 384941 695736 386522 695738
rect 384941 695680 384946 695736
rect 385002 695680 386522 695736
rect 384941 695678 386522 695680
rect 384941 695675 385007 695678
rect 386462 695605 386522 695678
rect 386597 695736 398807 695738
rect 386597 695680 386602 695736
rect 386658 695680 398746 695736
rect 398802 695680 398807 695736
rect 386597 695678 398807 695680
rect 386597 695675 386663 695678
rect 398741 695675 398807 695678
rect 403065 695738 403131 695741
rect 412582 695738 412588 695740
rect 403065 695736 412588 695738
rect 403065 695680 403070 695736
rect 403126 695680 412588 695736
rect 403065 695678 412588 695680
rect 403065 695675 403131 695678
rect 412582 695676 412588 695678
rect 412652 695676 412658 695740
rect 452561 695738 452627 695741
rect 463734 695738 463740 695740
rect 452561 695736 463740 695738
rect 452561 695680 452566 695736
rect 452622 695680 463740 695736
rect 452561 695678 463740 695680
rect 452561 695675 452627 695678
rect 463734 695676 463740 695678
rect 463804 695676 463810 695740
rect 482921 695738 482987 695741
rect 485773 695738 485839 695741
rect 482921 695736 485839 695738
rect 482921 695680 482926 695736
rect 482982 695680 485778 695736
rect 485834 695680 485839 695736
rect 482921 695678 485839 695680
rect 482921 695675 482987 695678
rect 485773 695675 485839 695678
rect 205541 695602 205607 695605
rect 181486 695600 205607 695602
rect 181486 695544 205546 695600
rect 205602 695544 205607 695600
rect 181486 695542 205607 695544
rect 205541 695539 205607 695542
rect 213729 695602 213795 695605
rect 215201 695602 215267 695605
rect 213729 695600 215267 695602
rect 213729 695544 213734 695600
rect 213790 695544 215206 695600
rect 215262 695544 215267 695600
rect 213729 695542 215267 695544
rect 213729 695539 213795 695542
rect 215201 695539 215267 695542
rect 230381 695602 230447 695605
rect 234521 695602 234587 695605
rect 230381 695600 234587 695602
rect 230381 695544 230386 695600
rect 230442 695544 234526 695600
rect 234582 695544 234587 695600
rect 230381 695542 234587 695544
rect 230381 695539 230447 695542
rect 234521 695539 234587 695542
rect 251081 695602 251147 695605
rect 253841 695602 253907 695605
rect 251081 695600 253907 695602
rect 251081 695544 251086 695600
rect 251142 695544 253846 695600
rect 253902 695544 253907 695600
rect 251081 695542 253907 695544
rect 251081 695539 251147 695542
rect 253841 695539 253907 695542
rect 299381 695602 299447 695605
rect 309133 695602 309199 695605
rect 299381 695600 309199 695602
rect 299381 695544 299386 695600
rect 299442 695544 309138 695600
rect 309194 695544 309199 695600
rect 299381 695542 309199 695544
rect 299381 695539 299447 695542
rect 309133 695539 309199 695542
rect 328361 695602 328427 695605
rect 331121 695602 331187 695605
rect 328361 695600 331187 695602
rect 328361 695544 328366 695600
rect 328422 695544 331126 695600
rect 331182 695544 331187 695600
rect 328361 695542 331187 695544
rect 328361 695539 328427 695542
rect 331121 695539 331187 695542
rect 347630 695540 347636 695604
rect 347700 695602 347706 695604
rect 357433 695602 357499 695605
rect 347700 695600 357499 695602
rect 347700 695544 357438 695600
rect 357494 695544 357499 695600
rect 347700 695542 357499 695544
rect 347700 695540 347706 695542
rect 357433 695539 357499 695542
rect 357617 695602 357683 695605
rect 360101 695602 360167 695605
rect 357617 695600 360167 695602
rect 357617 695544 357622 695600
rect 357678 695544 360106 695600
rect 360162 695544 360167 695600
rect 357617 695542 360167 695544
rect 357617 695539 357683 695542
rect 360101 695539 360167 695542
rect 371877 695602 371943 695605
rect 375373 695602 375439 695605
rect 371877 695600 375439 695602
rect 371877 695544 371882 695600
rect 371938 695544 375378 695600
rect 375434 695544 375439 695600
rect 371877 695542 375439 695544
rect 386462 695600 386571 695605
rect 386462 695544 386510 695600
rect 386566 695544 386571 695600
rect 386462 695542 386571 695544
rect 371877 695539 371943 695542
rect 375373 695539 375439 695542
rect 386505 695539 386571 695542
rect 398925 695602 398991 695605
rect 402973 695602 403039 695605
rect 398925 695600 403039 695602
rect 398925 695544 398930 695600
rect 398986 695544 402978 695600
rect 403034 695544 403039 695600
rect 398925 695542 403039 695544
rect 398925 695539 398991 695542
rect 402973 695539 403039 695542
rect 426382 695540 426388 695604
rect 426452 695602 426458 695604
rect 426525 695602 426591 695605
rect 426452 695600 426591 695602
rect 426452 695544 426530 695600
rect 426586 695544 426591 695600
rect 426452 695542 426591 695544
rect 426452 695540 426458 695542
rect 426525 695539 426591 695542
rect 426893 695602 426959 695605
rect 434662 695602 434668 695604
rect 426893 695600 434668 695602
rect 426893 695544 426898 695600
rect 426954 695544 434668 695600
rect 426893 695542 434668 695544
rect 426893 695539 426959 695542
rect 434662 695540 434668 695542
rect 434732 695540 434738 695604
rect 468477 695602 468543 695605
rect 473302 695602 473308 695604
rect 468477 695600 473308 695602
rect 468477 695544 468482 695600
rect 468538 695544 473308 695600
rect 468477 695542 473308 695544
rect 468477 695539 468543 695542
rect 473302 695540 473308 695542
rect 473372 695540 473378 695604
rect 492581 695602 492647 695605
rect 495390 695602 495450 695814
rect 505142 695738 505202 695814
rect 543825 695738 543891 695741
rect 553209 695738 553275 695741
rect 505142 695678 524522 695738
rect 492581 695600 495450 695602
rect 492581 695544 492586 695600
rect 492642 695544 495450 695600
rect 492581 695542 495450 695544
rect 524462 695602 524522 695678
rect 543825 695736 553275 695738
rect 543825 695680 543830 695736
rect 543886 695680 553214 695736
rect 553270 695680 553275 695736
rect 543825 695678 553275 695680
rect 543825 695675 543891 695678
rect 553209 695675 553275 695678
rect 553393 695738 553459 695741
rect 562317 695738 562383 695741
rect 553393 695736 562383 695738
rect 553393 695680 553398 695736
rect 553454 695680 562322 695736
rect 562378 695680 562383 695736
rect 553393 695678 562383 695680
rect 553393 695675 553459 695678
rect 562317 695675 562383 695678
rect 567101 695738 567167 695741
rect 569309 695738 569375 695741
rect 567101 695736 569375 695738
rect 567101 695680 567106 695736
rect 567162 695680 569314 695736
rect 569370 695680 569375 695736
rect 567101 695678 569375 695680
rect 567101 695675 567167 695678
rect 569309 695675 569375 695678
rect 540973 695602 541039 695605
rect 524462 695600 541039 695602
rect 524462 695544 540978 695600
rect 541034 695544 541039 695600
rect 524462 695542 541039 695544
rect 492581 695539 492647 695542
rect 540973 695539 541039 695542
rect 215293 695466 215359 695469
rect 229001 695466 229067 695469
rect 215293 695464 229067 695466
rect 215293 695408 215298 695464
rect 215354 695408 229006 695464
rect 229062 695408 229067 695464
rect 215293 695406 229067 695408
rect 215293 695403 215359 695406
rect 229001 695403 229067 695406
rect 442942 695404 442948 695468
rect 443012 695466 443018 695468
rect 452561 695466 452627 695469
rect 443012 695464 452627 695466
rect 443012 695408 452566 695464
rect 452622 695408 452627 695464
rect 443012 695406 452627 695408
rect 443012 695404 443018 695406
rect 452561 695403 452627 695406
rect 15377 695330 15443 695333
rect 157057 695332 157123 695333
rect 17166 695330 17172 695332
rect 15377 695328 17172 695330
rect 15377 695272 15382 695328
rect 15438 695272 17172 695328
rect 15377 695270 17172 695272
rect 15377 695267 15443 695270
rect 17166 695268 17172 695270
rect 17236 695268 17242 695332
rect 157006 695330 157012 695332
rect 156966 695270 157012 695330
rect 157076 695328 157123 695332
rect 157118 695272 157123 695328
rect 157006 695268 157012 695270
rect 157076 695268 157123 695272
rect 412582 695268 412588 695332
rect 412652 695330 412658 695332
rect 422201 695330 422267 695333
rect 521377 695332 521443 695333
rect 521326 695330 521332 695332
rect 412652 695328 422267 695330
rect 412652 695272 422206 695328
rect 422262 695272 422267 695328
rect 412652 695270 422267 695272
rect 521286 695270 521332 695330
rect 521396 695328 521443 695332
rect 521438 695272 521443 695328
rect 412652 695268 412658 695270
rect 157057 695267 157123 695268
rect 422201 695267 422267 695270
rect 521326 695268 521332 695270
rect 521396 695268 521443 695272
rect 521377 695267 521443 695268
rect 176510 694860 176516 694924
rect 176580 694922 176586 694924
rect 178902 694922 178908 694924
rect 176580 694862 178908 694922
rect 176580 694860 176586 694862
rect 178902 694860 178908 694862
rect 178972 694860 178978 694924
rect 311566 694860 311572 694924
rect 311636 694922 311642 694924
rect 311636 694862 318626 694922
rect 311636 694860 311642 694862
rect 124254 694724 124260 694788
rect 124324 694786 124330 694788
rect 133638 694786 133644 694788
rect 124324 694726 133644 694786
rect 124324 694724 124330 694726
rect 133638 694724 133644 694726
rect 133708 694724 133714 694788
rect 153326 694724 153332 694788
rect 153396 694786 153402 694788
rect 153396 694726 165538 694786
rect 153396 694724 153402 694726
rect 111006 694452 111012 694516
rect 111076 694514 111082 694516
rect 115606 694514 115612 694516
rect 111076 694454 115612 694514
rect 111076 694452 111082 694454
rect 115606 694452 115612 694454
rect 115676 694452 115682 694516
rect 165478 694514 165538 694726
rect 273294 694724 273300 694788
rect 273364 694786 273370 694788
rect 279918 694786 279924 694788
rect 273364 694726 279924 694786
rect 273364 694724 273370 694726
rect 279918 694724 279924 694726
rect 279988 694724 279994 694788
rect 299790 694724 299796 694788
rect 299860 694786 299866 694788
rect 311198 694786 311204 694788
rect 299860 694726 311204 694786
rect 299860 694724 299866 694726
rect 311198 694724 311204 694726
rect 311268 694724 311274 694788
rect 318566 694786 318626 694862
rect 321502 694860 321508 694924
rect 321572 694922 321578 694924
rect 323710 694922 323716 694924
rect 321572 694862 323716 694922
rect 321572 694860 321578 694862
rect 323710 694860 323716 694862
rect 323780 694860 323786 694924
rect 489678 694860 489684 694924
rect 489748 694922 489754 694924
rect 489748 694862 491218 694922
rect 489748 694860 489754 694862
rect 318742 694786 318748 694788
rect 318566 694726 318748 694786
rect 318742 694724 318748 694726
rect 318812 694724 318818 694788
rect 331070 694786 331076 694788
rect 328502 694726 331076 694786
rect 186262 694588 186268 694652
rect 186332 694650 186338 694652
rect 255998 694650 256004 694652
rect 186332 694590 256004 694650
rect 186332 694588 186338 694590
rect 255998 694588 256004 694590
rect 256068 694588 256074 694652
rect 275318 694588 275324 694652
rect 275388 694650 275394 694652
rect 284886 694650 284892 694652
rect 275388 694590 284892 694650
rect 275388 694588 275394 694590
rect 284886 694588 284892 694590
rect 284956 694588 284962 694652
rect 311750 694650 311756 694652
rect 299476 694590 311756 694650
rect 165478 694454 186882 694514
rect 96662 694318 106106 694378
rect 17166 694180 17172 694244
rect 17236 694242 17242 694244
rect 96662 694242 96722 694318
rect 17236 694182 96722 694242
rect 106046 694242 106106 694318
rect 133638 694316 133644 694380
rect 133708 694378 133714 694380
rect 153142 694378 153148 694380
rect 133708 694318 153148 694378
rect 133708 694316 133714 694318
rect 153142 694316 153148 694318
rect 153212 694316 153218 694380
rect 160870 694316 160876 694380
rect 160940 694378 160946 694380
rect 164182 694378 164188 694380
rect 160940 694318 164188 694378
rect 160940 694316 160946 694318
rect 164182 694316 164188 694318
rect 164252 694316 164258 694380
rect 185894 694316 185900 694380
rect 185964 694378 185970 694380
rect 186822 694378 186882 694454
rect 196014 694452 196020 694516
rect 196084 694514 196090 694516
rect 196084 694454 206202 694514
rect 196084 694452 196090 694454
rect 195830 694378 195836 694380
rect 185964 694318 186514 694378
rect 186822 694318 195836 694378
rect 185964 694316 185970 694318
rect 124254 694242 124260 694244
rect 106046 694182 124260 694242
rect 17236 694180 17242 694182
rect 124254 694180 124260 694182
rect 124324 694180 124330 694244
rect 178902 694180 178908 694244
rect 178972 694242 178978 694244
rect 178972 694182 186146 694242
rect 178972 694180 178978 694182
rect 6637 694106 6703 694109
rect 9622 694106 9628 694108
rect 6637 694104 9628 694106
rect 6637 694048 6642 694104
rect 6698 694048 9628 694104
rect 6637 694046 9628 694048
rect 6637 694043 6703 694046
rect 9622 694044 9628 694046
rect 9692 694044 9698 694108
rect 31518 694106 31524 694108
rect 19198 694046 31524 694106
rect 9806 693908 9812 693972
rect 9876 693970 9882 693972
rect 19198 693970 19258 694046
rect 31518 694044 31524 694046
rect 31588 694044 31594 694108
rect 89846 694044 89852 694108
rect 89916 694106 89922 694108
rect 96654 694106 96660 694108
rect 89916 694046 96660 694106
rect 89916 694044 89922 694046
rect 96654 694044 96660 694046
rect 96724 694044 96730 694108
rect 140814 694044 140820 694108
rect 140884 694106 140890 694108
rect 143574 694106 143580 694108
rect 140884 694046 143580 694106
rect 140884 694044 140890 694046
rect 143574 694044 143580 694046
rect 143644 694044 143650 694108
rect 152958 694044 152964 694108
rect 153028 694106 153034 694108
rect 160870 694106 160876 694108
rect 153028 694046 160876 694106
rect 153028 694044 153034 694046
rect 160870 694044 160876 694046
rect 160940 694044 160946 694108
rect 164182 694044 164188 694108
rect 164252 694106 164258 694108
rect 185894 694106 185900 694108
rect 164252 694046 185900 694106
rect 164252 694044 164258 694046
rect 185894 694044 185900 694046
rect 185964 694044 185970 694108
rect 186086 694106 186146 694182
rect 186262 694106 186268 694108
rect 186086 694046 186268 694106
rect 186262 694044 186268 694046
rect 186332 694044 186338 694108
rect 186454 694106 186514 694318
rect 195830 694316 195836 694318
rect 195900 694316 195906 694380
rect 206142 694378 206202 694454
rect 215334 694452 215340 694516
rect 215404 694514 215410 694516
rect 215404 694454 225522 694514
rect 215404 694452 215410 694454
rect 215150 694378 215156 694380
rect 206142 694318 215156 694378
rect 215150 694316 215156 694318
rect 215220 694316 215226 694380
rect 225462 694378 225522 694454
rect 234616 694454 244842 694514
rect 234616 694378 234676 694454
rect 225462 694318 234676 694378
rect 244782 694378 244842 694454
rect 263542 694452 263548 694516
rect 263612 694514 263618 694516
rect 273662 694514 273668 694516
rect 263612 694454 273668 694514
rect 263612 694452 263618 694454
rect 273662 694452 273668 694454
rect 273732 694452 273738 694516
rect 283046 694452 283052 694516
rect 283116 694514 283122 694516
rect 299476 694514 299536 694590
rect 311750 694588 311756 694590
rect 311820 694588 311826 694652
rect 318926 694588 318932 694652
rect 318996 694650 319002 694652
rect 328502 694650 328562 694726
rect 331070 694724 331076 694726
rect 331140 694724 331146 694788
rect 424910 694786 424916 694788
rect 410382 694726 424916 694786
rect 318996 694590 328562 694650
rect 318996 694588 319002 694590
rect 331254 694588 331260 694652
rect 331324 694650 331330 694652
rect 331324 694590 333530 694650
rect 331324 694588 331330 694590
rect 323526 694514 323532 694516
rect 283116 694454 293234 694514
rect 283116 694452 283122 694454
rect 253790 694378 253796 694380
rect 244782 694318 253796 694378
rect 253790 694316 253796 694318
rect 253860 694316 253866 694380
rect 254342 694316 254348 694380
rect 254412 694378 254418 694380
rect 254412 694318 268394 694378
rect 254412 694316 254418 694318
rect 255998 694180 256004 694244
rect 256068 694242 256074 694244
rect 268334 694242 268394 694318
rect 280056 694316 280062 694380
rect 280126 694378 280132 694380
rect 282678 694378 282684 694380
rect 280126 694318 282684 694378
rect 280126 694316 280132 694318
rect 282678 694316 282684 694318
rect 282748 694316 282754 694380
rect 283230 694316 283236 694380
rect 283300 694378 283306 694380
rect 293174 694378 293234 694454
rect 299430 694454 299536 694514
rect 318566 694454 323532 694514
rect 299430 694378 299490 694454
rect 311566 694378 311572 694380
rect 283300 694318 292130 694378
rect 293174 694318 299490 694378
rect 302926 694318 311572 694378
rect 283300 694316 283306 694318
rect 273294 694242 273300 694244
rect 256068 694182 263794 694242
rect 268334 694182 273300 694242
rect 256068 694180 256074 694182
rect 195830 694106 195836 694108
rect 186454 694046 195836 694106
rect 195830 694044 195836 694046
rect 195900 694044 195906 694108
rect 196014 694044 196020 694108
rect 196084 694106 196090 694108
rect 205398 694106 205404 694108
rect 196084 694046 205404 694106
rect 196084 694044 196090 694046
rect 205398 694044 205404 694046
rect 205468 694044 205474 694108
rect 205950 694044 205956 694108
rect 206020 694106 206026 694108
rect 215150 694106 215156 694108
rect 206020 694046 215156 694106
rect 206020 694044 206026 694046
rect 215150 694044 215156 694046
rect 215220 694044 215226 694108
rect 215334 694044 215340 694108
rect 215404 694106 215410 694108
rect 224718 694106 224724 694108
rect 215404 694046 224724 694106
rect 215404 694044 215410 694046
rect 224718 694044 224724 694046
rect 224788 694044 224794 694108
rect 225270 694044 225276 694108
rect 225340 694106 225346 694108
rect 244038 694106 244044 694108
rect 225340 694046 244044 694106
rect 225340 694044 225346 694046
rect 244038 694044 244044 694046
rect 244108 694044 244114 694108
rect 244590 694044 244596 694108
rect 244660 694106 244666 694108
rect 263542 694106 263548 694108
rect 244660 694046 263548 694106
rect 244660 694044 244666 694046
rect 263542 694044 263548 694046
rect 263612 694044 263618 694108
rect 263734 694106 263794 694182
rect 273294 694180 273300 694182
rect 273364 694180 273370 694244
rect 275318 694242 275324 694244
rect 273486 694182 275324 694242
rect 273486 694106 273546 694182
rect 275318 694180 275324 694182
rect 275388 694180 275394 694244
rect 292070 694242 292130 694318
rect 302926 694242 302986 694318
rect 311566 694316 311572 694318
rect 311636 694316 311642 694380
rect 311750 694316 311756 694380
rect 311820 694378 311826 694380
rect 318566 694378 318626 694454
rect 323526 694452 323532 694454
rect 323596 694452 323602 694516
rect 323710 694452 323716 694516
rect 323780 694514 323786 694516
rect 323780 694454 328424 694514
rect 323780 694452 323786 694454
rect 311820 694318 318626 694378
rect 311820 694316 311826 694318
rect 292070 694182 302986 694242
rect 328364 694242 328424 694454
rect 330702 694452 330708 694516
rect 330772 694514 330778 694516
rect 333470 694514 333530 694590
rect 340822 694588 340828 694652
rect 340892 694650 340898 694652
rect 371918 694650 371924 694652
rect 340892 694590 371924 694650
rect 340892 694588 340898 694590
rect 371918 694588 371924 694590
rect 371988 694588 371994 694652
rect 379094 694588 379100 694652
rect 379164 694650 379170 694652
rect 391238 694650 391244 694652
rect 379164 694590 391244 694650
rect 379164 694588 379170 694590
rect 391238 694588 391244 694590
rect 391308 694588 391314 694652
rect 398414 694588 398420 694652
rect 398484 694650 398490 694652
rect 410382 694650 410442 694726
rect 424910 694724 424916 694726
rect 424980 694724 424986 694788
rect 425094 694724 425100 694788
rect 425164 694786 425170 694788
rect 434294 694786 434300 694788
rect 425164 694726 434300 694786
rect 425164 694724 425170 694726
rect 434294 694724 434300 694726
rect 434364 694724 434370 694788
rect 461158 694724 461164 694788
rect 461228 694786 461234 694788
rect 470358 694786 470364 694788
rect 461228 694726 470364 694786
rect 461228 694724 461234 694726
rect 470358 694724 470364 694726
rect 470428 694724 470434 694788
rect 398484 694590 410442 694650
rect 398484 694588 398490 694590
rect 470542 694588 470548 694652
rect 470612 694650 470618 694652
rect 470612 694590 480178 694650
rect 470612 694588 470618 694590
rect 359958 694514 359964 694516
rect 330772 694454 333346 694514
rect 333470 694454 341442 694514
rect 330772 694452 330778 694454
rect 333286 694378 333346 694454
rect 341382 694378 341442 694454
rect 352606 694454 359964 694514
rect 352606 694378 352666 694454
rect 359958 694452 359964 694454
rect 360028 694452 360034 694516
rect 369894 694452 369900 694516
rect 369964 694514 369970 694516
rect 369964 694454 380082 694514
rect 369964 694452 369970 694454
rect 333286 694318 341074 694378
rect 341382 694318 352666 694378
rect 328364 694182 330954 694242
rect 263734 694046 273546 694106
rect 273662 694044 273668 694108
rect 273732 694106 273738 694108
rect 282862 694106 282868 694108
rect 273732 694046 282868 694106
rect 273732 694044 273738 694046
rect 282862 694044 282868 694046
rect 282932 694044 282938 694108
rect 284886 694044 284892 694108
rect 284956 694106 284962 694108
rect 299238 694106 299244 694108
rect 284956 694046 299244 694106
rect 284956 694044 284962 694046
rect 299238 694044 299244 694046
rect 299308 694044 299314 694108
rect 311198 694044 311204 694108
rect 311268 694106 311274 694108
rect 321502 694106 321508 694108
rect 311268 694046 321508 694106
rect 311268 694044 311274 694046
rect 321502 694044 321508 694046
rect 321572 694044 321578 694108
rect 323526 694044 323532 694108
rect 323596 694106 323602 694108
rect 330702 694106 330708 694108
rect 323596 694046 330708 694106
rect 323596 694044 323602 694046
rect 330702 694044 330708 694046
rect 330772 694044 330778 694108
rect 330894 694106 330954 694182
rect 340822 694106 340828 694108
rect 330894 694046 340828 694106
rect 340822 694044 340828 694046
rect 340892 694044 340898 694108
rect 341014 694106 341074 694318
rect 360326 694316 360332 694380
rect 360396 694378 360402 694380
rect 369710 694378 369716 694380
rect 360396 694318 369716 694378
rect 360396 694316 360402 694318
rect 369710 694316 369716 694318
rect 369780 694316 369786 694380
rect 380022 694378 380082 694454
rect 390134 694452 390140 694516
rect 390204 694514 390210 694516
rect 390204 694454 399402 694514
rect 390204 694452 390210 694454
rect 389214 694378 389220 694380
rect 380022 694318 389220 694378
rect 389214 694316 389220 694318
rect 389284 694316 389290 694380
rect 399342 694378 399402 694454
rect 410566 694454 420010 694514
rect 410566 694378 410626 694454
rect 399342 694318 410626 694378
rect 419950 694378 420010 694454
rect 420126 694452 420132 694516
rect 420196 694514 420202 694516
rect 426382 694514 426388 694516
rect 420196 694454 426388 694514
rect 420196 694452 420202 694454
rect 426382 694452 426388 694454
rect 426452 694452 426458 694516
rect 433382 694454 434730 694514
rect 433382 694378 433442 694454
rect 419950 694318 433442 694378
rect 434670 694378 434730 694454
rect 434670 694318 447058 694378
rect 371918 694180 371924 694244
rect 371988 694242 371994 694244
rect 379094 694242 379100 694244
rect 371988 694182 379100 694242
rect 371988 694180 371994 694182
rect 379094 694180 379100 694182
rect 379164 694180 379170 694244
rect 391238 694180 391244 694244
rect 391308 694242 391314 694244
rect 398414 694242 398420 694244
rect 391308 694182 398420 694242
rect 391308 694180 391314 694182
rect 398414 694180 398420 694182
rect 398484 694180 398490 694244
rect 420310 694180 420316 694244
rect 420380 694242 420386 694244
rect 424726 694242 424732 694244
rect 420380 694182 424732 694242
rect 420380 694180 420386 694182
rect 424726 694180 424732 694182
rect 424796 694180 424802 694244
rect 424910 694180 424916 694244
rect 424980 694180 424986 694244
rect 446998 694242 447058 694318
rect 470358 694316 470364 694380
rect 470428 694378 470434 694380
rect 470542 694378 470548 694380
rect 470428 694318 470548 694378
rect 470428 694316 470434 694318
rect 470542 694316 470548 694318
rect 470612 694316 470618 694380
rect 480118 694378 480178 694590
rect 491158 694514 491218 694862
rect 531262 694724 531268 694788
rect 531332 694786 531338 694788
rect 531332 694726 539610 694786
rect 531332 694724 531338 694726
rect 511942 694588 511948 694652
rect 512012 694650 512018 694652
rect 521510 694650 521516 694652
rect 512012 694590 521516 694650
rect 512012 694588 512018 694590
rect 521510 694588 521516 694590
rect 521580 694588 521586 694652
rect 539550 694650 539610 694726
rect 539550 694590 539794 694650
rect 491158 694454 495634 694514
rect 489494 694378 489500 694380
rect 480118 694318 489500 694378
rect 489494 694316 489500 694318
rect 489564 694316 489570 694380
rect 460974 694242 460980 694244
rect 446998 694182 460980 694242
rect 460974 694180 460980 694182
rect 461044 694180 461050 694244
rect 495574 694242 495634 694454
rect 500902 694452 500908 694516
rect 500972 694514 500978 694516
rect 500972 694454 521578 694514
rect 500972 694452 500978 694454
rect 500902 694242 500908 694244
rect 495574 694182 500908 694242
rect 500902 694180 500908 694182
rect 500972 694180 500978 694244
rect 521518 694242 521578 694454
rect 521694 694452 521700 694516
rect 521764 694514 521770 694516
rect 531262 694514 531268 694516
rect 521764 694454 531268 694514
rect 521764 694452 521770 694454
rect 531262 694452 531268 694454
rect 531332 694452 531338 694516
rect 539734 694514 539794 694590
rect 550582 694514 550588 694516
rect 539734 694454 550588 694514
rect 550582 694452 550588 694454
rect 550652 694452 550658 694516
rect 576117 694378 576183 694381
rect 563102 694376 576183 694378
rect 563102 694320 576122 694376
rect 576178 694320 576183 694376
rect 563102 694318 576183 694320
rect 521694 694242 521700 694244
rect 521518 694182 521700 694242
rect 521694 694180 521700 694182
rect 521764 694180 521770 694244
rect 550582 694180 550588 694244
rect 550652 694242 550658 694244
rect 563102 694242 563162 694318
rect 576117 694315 576183 694318
rect 550652 694182 563162 694242
rect 550652 694180 550658 694182
rect 359958 694106 359964 694108
rect 341014 694046 359964 694106
rect 359958 694044 359964 694046
rect 360028 694044 360034 694108
rect 360326 694044 360332 694108
rect 360396 694106 360402 694108
rect 369710 694106 369716 694108
rect 360396 694046 369716 694106
rect 360396 694044 360402 694046
rect 369710 694044 369716 694046
rect 369780 694044 369786 694108
rect 369894 694044 369900 694108
rect 369964 694106 369970 694108
rect 420126 694106 420132 694108
rect 369964 694046 420132 694106
rect 369964 694044 369970 694046
rect 420126 694044 420132 694046
rect 420196 694044 420202 694108
rect 424918 694106 424978 694180
rect 425094 694106 425100 694108
rect 424918 694046 425100 694106
rect 425094 694044 425100 694046
rect 425164 694044 425170 694108
rect 434478 694044 434484 694108
rect 434548 694106 434554 694108
rect 434662 694106 434668 694108
rect 434548 694046 434668 694106
rect 434548 694044 434554 694046
rect 434662 694044 434668 694046
rect 434732 694044 434738 694108
rect 435030 694044 435036 694108
rect 435100 694106 435106 694108
rect 511942 694106 511948 694108
rect 435100 694046 511948 694106
rect 435100 694044 435106 694046
rect 511942 694044 511948 694046
rect 512012 694044 512018 694108
rect 521510 694044 521516 694108
rect 521580 694106 521586 694108
rect 521694 694106 521700 694108
rect 521580 694046 521700 694106
rect 521580 694044 521586 694046
rect 521694 694044 521700 694046
rect 521764 694044 521770 694108
rect 524454 694044 524460 694108
rect 524524 694106 524530 694108
rect 539542 694106 539548 694108
rect 524524 694046 539548 694106
rect 524524 694044 524530 694046
rect 539542 694044 539548 694046
rect 539612 694044 539618 694108
rect 9876 693910 19258 693970
rect 9876 693908 9882 693910
rect 31886 693908 31892 693972
rect 31956 693970 31962 693972
rect 37222 693970 37228 693972
rect 31956 693910 37228 693970
rect 31956 693908 31962 693910
rect 37222 693908 37228 693910
rect 37292 693908 37298 693972
rect 46790 693908 46796 693972
rect 46860 693970 46866 693972
rect 56542 693970 56548 693972
rect 46860 693910 56548 693970
rect 46860 693908 46866 693910
rect 56542 693908 56548 693910
rect 56612 693908 56618 693972
rect 66110 693908 66116 693972
rect 66180 693970 66186 693972
rect 75862 693970 75868 693972
rect 66180 693910 75868 693970
rect 66180 693908 66186 693910
rect 75862 693908 75868 693910
rect 75932 693908 75938 693972
rect 85430 693908 85436 693972
rect 85500 693970 85506 693972
rect 89478 693970 89484 693972
rect 85500 693910 89484 693970
rect 85500 693908 85506 693910
rect 89478 693908 89484 693910
rect 89548 693908 89554 693972
rect 96838 693908 96844 693972
rect 96908 693970 96914 693972
rect 111006 693970 111012 693972
rect 96908 693910 111012 693970
rect 96908 693908 96914 693910
rect 111006 693908 111012 693910
rect 111076 693908 111082 693972
rect 115606 693908 115612 693972
rect 115676 693970 115682 693972
rect 124254 693970 124260 693972
rect 115676 693910 124260 693970
rect 115676 693908 115682 693910
rect 124254 693908 124260 693910
rect 124324 693908 124330 693972
rect 133638 693908 133644 693972
rect 133708 693970 133714 693972
rect 140630 693970 140636 693972
rect 133708 693910 140636 693970
rect 133708 693908 133714 693910
rect 140630 693908 140636 693910
rect 140700 693908 140706 693972
rect 157006 693908 157012 693972
rect 157076 693970 157082 693972
rect 173934 693970 173940 693972
rect 157076 693910 173940 693970
rect 157076 693908 157082 693910
rect 173934 693908 173940 693910
rect 174004 693908 174010 693972
rect 174118 693908 174124 693972
rect 174188 693970 174194 693972
rect 420310 693970 420316 693972
rect 174188 693910 420316 693970
rect 174188 693908 174194 693910
rect 420310 693908 420316 693910
rect 420380 693908 420386 693972
rect 424910 693908 424916 693972
rect 424980 693970 424986 693972
rect 434662 693970 434668 693972
rect 424980 693910 434668 693970
rect 424980 693908 424986 693910
rect 434662 693908 434668 693910
rect 434732 693908 434738 693972
rect 435030 693908 435036 693972
rect 435100 693970 435106 693972
rect 543590 693970 543596 693972
rect 435100 693910 543596 693970
rect 435100 693908 435106 693910
rect 543590 693908 543596 693910
rect 543660 693908 543666 693972
rect 543774 693908 543780 693972
rect 543844 693970 543850 693972
rect 562910 693970 562916 693972
rect 543844 693910 562916 693970
rect 543844 693908 543850 693910
rect 562910 693908 562916 693910
rect 562980 693908 562986 693972
rect 563094 693908 563100 693972
rect 563164 693970 563170 693972
rect 577957 693970 578023 693973
rect 563164 693968 578023 693970
rect 563164 693912 577962 693968
rect 578018 693912 578023 693968
rect 563164 693910 578023 693912
rect 563164 693908 563170 693910
rect 577957 693907 578023 693910
rect 3417 693834 3483 693837
rect 55622 693834 55628 693836
rect 3417 693832 55628 693834
rect 3417 693776 3422 693832
rect 3478 693776 55628 693832
rect 3417 693774 55628 693776
rect 3417 693771 3483 693774
rect 55622 693772 55628 693774
rect 55692 693772 55698 693836
rect 56358 693772 56364 693836
rect 56428 693834 56434 693836
rect 74942 693834 74948 693836
rect 56428 693774 74948 693834
rect 56428 693772 56434 693774
rect 74942 693772 74948 693774
rect 75012 693772 75018 693836
rect 75678 693772 75684 693836
rect 75748 693834 75754 693836
rect 108798 693834 108804 693836
rect 75748 693774 108804 693834
rect 75748 693772 75754 693774
rect 108798 693772 108804 693774
rect 108868 693772 108874 693836
rect 114134 693772 114140 693836
rect 114204 693834 114210 693836
rect 162894 693834 162900 693836
rect 114204 693774 162900 693834
rect 114204 693772 114210 693774
rect 162894 693772 162900 693774
rect 162964 693772 162970 693836
rect 163814 693772 163820 693836
rect 163884 693834 163890 693836
rect 424174 693834 424180 693836
rect 163884 693774 424180 693834
rect 163884 693772 163890 693774
rect 424174 693772 424180 693774
rect 424244 693772 424250 693836
rect 424910 693772 424916 693836
rect 424980 693834 424986 693836
rect 434110 693834 434116 693836
rect 424980 693774 434116 693834
rect 424980 693772 424986 693774
rect 434110 693772 434116 693774
rect 434180 693772 434186 693836
rect 434478 693772 434484 693836
rect 434548 693834 434554 693836
rect 434662 693834 434668 693836
rect 434548 693774 434668 693834
rect 434548 693772 434554 693774
rect 434662 693772 434668 693774
rect 434732 693772 434738 693836
rect 435214 693772 435220 693836
rect 435284 693834 435290 693836
rect 503478 693834 503484 693836
rect 435284 693774 503484 693834
rect 435284 693772 435290 693774
rect 503478 693772 503484 693774
rect 503548 693772 503554 693836
rect 521694 693772 521700 693836
rect 521764 693834 521770 693836
rect 524454 693834 524460 693836
rect 521764 693774 524460 693834
rect 521764 693772 521770 693774
rect 524454 693772 524460 693774
rect 524524 693772 524530 693836
rect 549110 693772 549116 693836
rect 549180 693834 549186 693836
rect 568481 693834 568547 693837
rect 549180 693774 550650 693834
rect 549180 693772 549186 693774
rect 7649 693698 7715 693701
rect 550590 693700 550650 693774
rect 568481 693832 569970 693834
rect 568481 693776 568486 693832
rect 568542 693776 569970 693832
rect 568481 693774 569970 693776
rect 568481 693771 568547 693774
rect 123702 693698 123708 693700
rect 7649 693696 123708 693698
rect 7649 693640 7654 693696
rect 7710 693640 123708 693696
rect 7649 693638 123708 693640
rect 7649 693635 7715 693638
rect 123702 693636 123708 693638
rect 123772 693636 123778 693700
rect 124070 693636 124076 693700
rect 124140 693698 124146 693700
rect 163078 693698 163084 693700
rect 124140 693638 163084 693698
rect 124140 693636 124146 693638
rect 163078 693636 163084 693638
rect 163148 693636 163154 693700
rect 163630 693636 163636 693700
rect 163700 693698 163706 693700
rect 423990 693698 423996 693700
rect 163700 693638 423996 693698
rect 163700 693636 163706 693638
rect 423990 693636 423996 693638
rect 424060 693636 424066 693700
rect 424726 693636 424732 693700
rect 424796 693698 424802 693700
rect 433926 693698 433932 693700
rect 424796 693638 433932 693698
rect 424796 693636 424802 693638
rect 433926 693636 433932 693638
rect 433996 693636 434002 693700
rect 434478 693636 434484 693700
rect 434548 693698 434554 693700
rect 473486 693698 473492 693700
rect 434548 693638 473492 693698
rect 434548 693636 434554 693638
rect 473486 693636 473492 693638
rect 473556 693636 473562 693700
rect 474038 693636 474044 693700
rect 474108 693698 474114 693700
rect 521326 693698 521332 693700
rect 474108 693638 521332 693698
rect 474108 693636 474114 693638
rect 521326 693636 521332 693638
rect 521396 693636 521402 693700
rect 550582 693636 550588 693700
rect 550652 693636 550658 693700
rect 550766 693636 550772 693700
rect 550836 693698 550842 693700
rect 558862 693698 558868 693700
rect 550836 693638 558868 693698
rect 550836 693636 550842 693638
rect 558862 693636 558868 693638
rect 558932 693636 558938 693700
rect 569910 693562 569970 693774
rect 579429 693562 579495 693565
rect 569910 693560 579495 693562
rect 569910 693504 579434 693560
rect 579490 693504 579495 693560
rect 569910 693502 579495 693504
rect 579429 693499 579495 693502
rect 565670 693364 565676 693428
rect 565740 693426 565746 693428
rect 568481 693426 568547 693429
rect 565740 693424 568547 693426
rect 565740 693368 568486 693424
rect 568542 693368 568547 693424
rect 565740 693366 568547 693368
rect 565740 693364 565746 693366
rect 568481 693363 568547 693366
rect 580901 686354 580967 686357
rect 583520 686354 584960 686444
rect 580901 686352 584960 686354
rect 580901 686296 580906 686352
rect 580962 686296 584960 686352
rect 580901 686294 584960 686296
rect 580901 686291 580967 686294
rect 583520 686204 584960 686294
rect -960 682274 480 682364
rect 2957 682274 3023 682277
rect -960 682272 3023 682274
rect -960 682216 2962 682272
rect 3018 682216 3023 682272
rect -960 682214 3023 682216
rect -960 682124 480 682214
rect 2957 682211 3023 682214
rect 579797 674658 579863 674661
rect 583520 674658 584960 674748
rect 579797 674656 584960 674658
rect 579797 674600 579802 674656
rect 579858 674600 584960 674656
rect 579797 674598 584960 674600
rect 579797 674595 579863 674598
rect 583520 674508 584960 674598
rect -960 667994 480 668084
rect 2773 667994 2839 667997
rect -960 667992 2839 667994
rect -960 667936 2778 667992
rect 2834 667936 2839 667992
rect -960 667934 2839 667936
rect -960 667844 480 667934
rect 2773 667931 2839 667934
rect 583520 662676 584960 662916
rect -960 653578 480 653668
rect 3049 653578 3115 653581
rect -960 653576 3115 653578
rect -960 653520 3054 653576
rect 3110 653520 3115 653576
rect -960 653518 3115 653520
rect -960 653428 480 653518
rect 3049 653515 3115 653518
rect 579613 651130 579679 651133
rect 583520 651130 584960 651220
rect 579613 651128 584960 651130
rect 579613 651072 579618 651128
rect 579674 651072 584960 651128
rect 579613 651070 584960 651072
rect 579613 651067 579679 651070
rect 583520 650980 584960 651070
rect 580901 639434 580967 639437
rect 583520 639434 584960 639524
rect 580901 639432 584960 639434
rect 580901 639376 580906 639432
rect 580962 639376 584960 639432
rect 580901 639374 584960 639376
rect 580901 639371 580967 639374
rect 583520 639284 584960 639374
rect -960 639012 480 639252
rect 574645 628010 574711 628013
rect 575473 628010 575539 628013
rect 574645 628008 575539 628010
rect 574645 627952 574650 628008
rect 574706 627952 575478 628008
rect 575534 627952 575539 628008
rect 574645 627950 575539 627952
rect 574645 627947 574711 627950
rect 575473 627947 575539 627950
rect 579797 627738 579863 627741
rect 583520 627738 584960 627828
rect 579797 627736 584960 627738
rect 579797 627680 579802 627736
rect 579858 627680 584960 627736
rect 579797 627678 584960 627680
rect 579797 627675 579863 627678
rect 583520 627588 584960 627678
rect -960 624882 480 624972
rect 2957 624882 3023 624885
rect -960 624880 3023 624882
rect -960 624824 2962 624880
rect 3018 624824 3023 624880
rect -960 624822 3023 624824
rect -960 624732 480 624822
rect 2957 624819 3023 624822
rect 583520 615756 584960 615996
rect -960 610466 480 610556
rect 3141 610466 3207 610469
rect -960 610464 3207 610466
rect -960 610408 3146 610464
rect 3202 610408 3207 610464
rect -960 610406 3207 610408
rect -960 610316 480 610406
rect 3141 610403 3207 610406
rect 579613 604210 579679 604213
rect 583520 604210 584960 604300
rect 579613 604208 584960 604210
rect 579613 604152 579618 604208
rect 579674 604152 584960 604208
rect 579613 604150 584960 604152
rect 579613 604147 579679 604150
rect 583520 604060 584960 604150
rect -960 596050 480 596140
rect 3141 596050 3207 596053
rect -960 596048 3207 596050
rect -960 595992 3146 596048
rect 3202 595992 3207 596048
rect -960 595990 3207 595992
rect -960 595900 480 595990
rect 3141 595987 3207 595990
rect 579521 592514 579587 592517
rect 583520 592514 584960 592604
rect 579521 592512 584960 592514
rect 579521 592456 579526 592512
rect 579582 592456 584960 592512
rect 579521 592454 584960 592456
rect 579521 592451 579587 592454
rect 583520 592364 584960 592454
rect -960 581620 480 581860
rect 580165 580818 580231 580821
rect 583520 580818 584960 580908
rect 580165 580816 584960 580818
rect 580165 580760 580170 580816
rect 580226 580760 584960 580816
rect 580165 580758 584960 580760
rect 580165 580755 580231 580758
rect 583520 580668 584960 580758
rect 583520 568836 584960 569076
rect -960 567354 480 567444
rect 3049 567354 3115 567357
rect -960 567352 3115 567354
rect -960 567296 3054 567352
rect 3110 567296 3115 567352
rect -960 567294 3115 567296
rect -960 567204 480 567294
rect 3049 567291 3115 567294
rect 579613 557290 579679 557293
rect 583520 557290 584960 557380
rect 579613 557288 584960 557290
rect 579613 557232 579618 557288
rect 579674 557232 584960 557288
rect 579613 557230 584960 557232
rect 579613 557227 579679 557230
rect 583520 557140 584960 557230
rect -960 553074 480 553164
rect 3877 553074 3943 553077
rect -960 553072 3943 553074
rect -960 553016 3882 553072
rect 3938 553016 3943 553072
rect -960 553014 3943 553016
rect -960 552924 480 553014
rect 3877 553011 3943 553014
rect 579429 545594 579495 545597
rect 583520 545594 584960 545684
rect 579429 545592 584960 545594
rect 579429 545536 579434 545592
rect 579490 545536 584960 545592
rect 579429 545534 584960 545536
rect 579429 545531 579495 545534
rect 583520 545444 584960 545534
rect -960 538658 480 538748
rect 3233 538658 3299 538661
rect -960 538656 3299 538658
rect -960 538600 3238 538656
rect 3294 538600 3299 538656
rect -960 538598 3299 538600
rect -960 538508 480 538598
rect 3233 538595 3299 538598
rect 579797 533898 579863 533901
rect 583520 533898 584960 533988
rect 579797 533896 584960 533898
rect 579797 533840 579802 533896
rect 579858 533840 584960 533896
rect 579797 533838 584960 533840
rect 579797 533835 579863 533838
rect 583520 533748 584960 533838
rect -960 524092 480 524332
rect 583520 521916 584960 522156
rect 580073 510370 580139 510373
rect 583520 510370 584960 510460
rect 580073 510368 584960 510370
rect 580073 510312 580078 510368
rect 580134 510312 584960 510368
rect 580073 510310 584960 510312
rect 580073 510307 580139 510310
rect 583520 510220 584960 510310
rect -960 509962 480 510052
rect 3049 509962 3115 509965
rect -960 509960 3115 509962
rect -960 509904 3054 509960
rect 3110 509904 3115 509960
rect -960 509902 3115 509904
rect -960 509812 480 509902
rect 3049 509899 3115 509902
rect 579337 498674 579403 498677
rect 583520 498674 584960 498764
rect 579337 498672 584960 498674
rect 579337 498616 579342 498672
rect 579398 498616 584960 498672
rect 579337 498614 584960 498616
rect 579337 498611 579403 498614
rect 583520 498524 584960 498614
rect -960 495546 480 495636
rect 3325 495546 3391 495549
rect -960 495544 3391 495546
rect -960 495488 3330 495544
rect 3386 495488 3391 495544
rect -960 495486 3391 495488
rect -960 495396 480 495486
rect 3325 495483 3391 495486
rect 580165 486842 580231 486845
rect 583520 486842 584960 486932
rect 580165 486840 584960 486842
rect 580165 486784 580170 486840
rect 580226 486784 584960 486840
rect 580165 486782 584960 486784
rect 580165 486779 580231 486782
rect 583520 486692 584960 486782
rect -960 481130 480 481220
rect 3325 481130 3391 481133
rect -960 481128 3391 481130
rect -960 481072 3330 481128
rect 3386 481072 3391 481128
rect -960 481070 3391 481072
rect -960 480980 480 481070
rect 3325 481067 3391 481070
rect 583520 474996 584960 475236
rect -960 466700 480 466940
rect 580809 463450 580875 463453
rect 583520 463450 584960 463540
rect 580809 463448 584960 463450
rect 580809 463392 580814 463448
rect 580870 463392 584960 463448
rect 580809 463390 584960 463392
rect 580809 463387 580875 463390
rect 583520 463300 584960 463390
rect -960 452434 480 452524
rect 3325 452434 3391 452437
rect -960 452432 3391 452434
rect -960 452376 3330 452432
rect 3386 452376 3391 452432
rect -960 452374 3391 452376
rect -960 452284 480 452374
rect 3325 452371 3391 452374
rect 579245 451754 579311 451757
rect 583520 451754 584960 451844
rect 579245 451752 584960 451754
rect 579245 451696 579250 451752
rect 579306 451696 584960 451752
rect 579245 451694 584960 451696
rect 579245 451691 579311 451694
rect 583520 451604 584960 451694
rect 579981 439922 580047 439925
rect 583520 439922 584960 440012
rect 579981 439920 584960 439922
rect 579981 439864 579986 439920
rect 580042 439864 584960 439920
rect 579981 439862 584960 439864
rect 579981 439859 580047 439862
rect 583520 439772 584960 439862
rect -960 438018 480 438108
rect 4061 438018 4127 438021
rect -960 438016 4127 438018
rect -960 437960 4066 438016
rect 4122 437960 4127 438016
rect -960 437958 4127 437960
rect -960 437868 480 437958
rect 4061 437955 4127 437958
rect 583520 428076 584960 428316
rect -960 423738 480 423828
rect 2865 423738 2931 423741
rect -960 423736 2931 423738
rect -960 423680 2870 423736
rect 2926 423680 2931 423736
rect -960 423678 2931 423680
rect -960 423588 480 423678
rect 2865 423675 2931 423678
rect 579613 416530 579679 416533
rect 583520 416530 584960 416620
rect 579613 416528 584960 416530
rect 579613 416472 579618 416528
rect 579674 416472 584960 416528
rect 579613 416470 584960 416472
rect 579613 416467 579679 416470
rect 583520 416380 584960 416470
rect -960 409172 480 409412
rect 580717 404834 580783 404837
rect 583520 404834 584960 404924
rect 580717 404832 584960 404834
rect 580717 404776 580722 404832
rect 580778 404776 584960 404832
rect 580717 404774 584960 404776
rect 580717 404771 580783 404774
rect 583520 404684 584960 404774
rect -960 395042 480 395132
rect 3233 395042 3299 395045
rect -960 395040 3299 395042
rect -960 394984 3238 395040
rect 3294 394984 3299 395040
rect -960 394982 3299 394984
rect -960 394892 480 394982
rect 3233 394979 3299 394982
rect 579613 393002 579679 393005
rect 583520 393002 584960 393092
rect 579613 393000 584960 393002
rect 579613 392944 579618 393000
rect 579674 392944 584960 393000
rect 579613 392942 584960 392944
rect 579613 392939 579679 392942
rect 583520 392852 584960 392942
rect 583520 381156 584960 381396
rect -960 380626 480 380716
rect 2773 380626 2839 380629
rect -960 380624 2839 380626
rect -960 380568 2778 380624
rect 2834 380568 2839 380624
rect -960 380566 2839 380568
rect -960 380476 480 380566
rect 2773 380563 2839 380566
rect 580717 369610 580783 369613
rect 583520 369610 584960 369700
rect 580717 369608 584960 369610
rect 580717 369552 580722 369608
rect 580778 369552 584960 369608
rect 580717 369550 584960 369552
rect 580717 369547 580783 369550
rect 583520 369460 584960 369550
rect -960 366210 480 366300
rect 3233 366210 3299 366213
rect -960 366208 3299 366210
rect -960 366152 3238 366208
rect 3294 366152 3299 366208
rect -960 366150 3299 366152
rect -960 366060 480 366150
rect 3233 366147 3299 366150
rect 579153 357914 579219 357917
rect 583520 357914 584960 358004
rect 579153 357912 584960 357914
rect 579153 357856 579158 357912
rect 579214 357856 584960 357912
rect 579153 357854 584960 357856
rect 579153 357851 579219 357854
rect 583520 357764 584960 357854
rect -960 351780 480 352020
rect 580165 346082 580231 346085
rect 583520 346082 584960 346172
rect 580165 346080 584960 346082
rect 580165 346024 580170 346080
rect 580226 346024 584960 346080
rect 580165 346022 584960 346024
rect 580165 346019 580231 346022
rect 583520 345932 584960 346022
rect -960 337514 480 337604
rect 3233 337514 3299 337517
rect -960 337512 3299 337514
rect -960 337456 3238 337512
rect 3294 337456 3299 337512
rect -960 337454 3299 337456
rect -960 337364 480 337454
rect 3233 337451 3299 337454
rect 583520 334236 584960 334476
rect -960 323098 480 323188
rect 3969 323098 4035 323101
rect -960 323096 4035 323098
rect -960 323040 3974 323096
rect 4030 323040 4035 323096
rect -960 323038 4035 323040
rect -960 322948 480 323038
rect 3969 323035 4035 323038
rect 580625 322690 580691 322693
rect 583520 322690 584960 322780
rect 580625 322688 584960 322690
rect 580625 322632 580630 322688
rect 580686 322632 584960 322688
rect 580625 322630 584960 322632
rect 580625 322627 580691 322630
rect 583520 322540 584960 322630
rect 579061 310858 579127 310861
rect 583520 310858 584960 310948
rect 579061 310856 584960 310858
rect 579061 310800 579066 310856
rect 579122 310800 584960 310856
rect 579061 310798 584960 310800
rect 579061 310795 579127 310798
rect 583520 310708 584960 310798
rect -960 308818 480 308908
rect 3233 308818 3299 308821
rect -960 308816 3299 308818
rect -960 308760 3238 308816
rect 3294 308760 3299 308816
rect -960 308758 3299 308760
rect -960 308668 480 308758
rect 3233 308755 3299 308758
rect 580165 299162 580231 299165
rect 583520 299162 584960 299252
rect 580165 299160 584960 299162
rect 580165 299104 580170 299160
rect 580226 299104 584960 299160
rect 580165 299102 584960 299104
rect 580165 299099 580231 299102
rect 583520 299012 584960 299102
rect -960 294402 480 294492
rect 3233 294402 3299 294405
rect -960 294400 3299 294402
rect -960 294344 3238 294400
rect 3294 294344 3299 294400
rect -960 294342 3299 294344
rect -960 294252 480 294342
rect 3233 294339 3299 294342
rect 583520 287316 584960 287556
rect -960 280122 480 280212
rect 2773 280122 2839 280125
rect -960 280120 2839 280122
rect -960 280064 2778 280120
rect 2834 280064 2839 280120
rect -960 280062 2839 280064
rect -960 279972 480 280062
rect 2773 280059 2839 280062
rect 579613 275770 579679 275773
rect 583520 275770 584960 275860
rect 579613 275768 584960 275770
rect 579613 275712 579618 275768
rect 579674 275712 584960 275768
rect 579613 275710 584960 275712
rect 579613 275707 579679 275710
rect 583520 275620 584960 275710
rect -960 265706 480 265796
rect 2957 265706 3023 265709
rect -960 265704 3023 265706
rect -960 265648 2962 265704
rect 3018 265648 3023 265704
rect -960 265646 3023 265648
rect -960 265556 480 265646
rect 2957 265643 3023 265646
rect 578969 263938 579035 263941
rect 583520 263938 584960 264028
rect 578969 263936 584960 263938
rect 578969 263880 578974 263936
rect 579030 263880 584960 263936
rect 578969 263878 584960 263880
rect 578969 263875 579035 263878
rect 583520 263788 584960 263878
rect 580165 252242 580231 252245
rect 583520 252242 584960 252332
rect 580165 252240 584960 252242
rect 580165 252184 580170 252240
rect 580226 252184 584960 252240
rect 580165 252182 584960 252184
rect 580165 252179 580231 252182
rect 583520 252092 584960 252182
rect -960 251290 480 251380
rect 3233 251290 3299 251293
rect -960 251288 3299 251290
rect -960 251232 3238 251288
rect 3294 251232 3299 251288
rect -960 251230 3299 251232
rect -960 251140 480 251230
rect 3233 251227 3299 251230
rect 583520 240396 584960 240636
rect -960 237010 480 237100
rect 3325 237010 3391 237013
rect -960 237008 3391 237010
rect -960 236952 3330 237008
rect 3386 236952 3391 237008
rect -960 236950 3391 236952
rect -960 236860 480 236950
rect 3325 236947 3391 236950
rect 580533 228850 580599 228853
rect 583520 228850 584960 228940
rect 580533 228848 584960 228850
rect 580533 228792 580538 228848
rect 580594 228792 584960 228848
rect 580533 228790 584960 228792
rect 580533 228787 580599 228790
rect 583520 228700 584960 228790
rect -960 222594 480 222684
rect 3785 222594 3851 222597
rect -960 222592 3851 222594
rect -960 222536 3790 222592
rect 3846 222536 3851 222592
rect -960 222534 3851 222536
rect -960 222444 480 222534
rect 3785 222531 3851 222534
rect 578877 217018 578943 217021
rect 583520 217018 584960 217108
rect 578877 217016 584960 217018
rect 578877 216960 578882 217016
rect 578938 216960 584960 217016
rect 578877 216958 584960 216960
rect 578877 216955 578943 216958
rect 583520 216868 584960 216958
rect -960 208178 480 208268
rect 3325 208178 3391 208181
rect -960 208176 3391 208178
rect -960 208120 3330 208176
rect 3386 208120 3391 208176
rect -960 208118 3391 208120
rect -960 208028 480 208118
rect 3325 208115 3391 208118
rect 580165 205322 580231 205325
rect 583520 205322 584960 205412
rect 580165 205320 584960 205322
rect 580165 205264 580170 205320
rect 580226 205264 584960 205320
rect 580165 205262 584960 205264
rect 580165 205259 580231 205262
rect 583520 205172 584960 205262
rect -960 193898 480 193988
rect 2773 193898 2839 193901
rect -960 193896 2839 193898
rect -960 193840 2778 193896
rect 2834 193840 2839 193896
rect -960 193838 2839 193840
rect -960 193748 480 193838
rect 2773 193835 2839 193838
rect 583520 193476 584960 193716
rect 580441 181930 580507 181933
rect 583520 181930 584960 182020
rect 580441 181928 584960 181930
rect 580441 181872 580446 181928
rect 580502 181872 584960 181928
rect 580441 181870 584960 181872
rect 580441 181867 580507 181870
rect 583520 181780 584960 181870
rect -960 179482 480 179572
rect 3693 179482 3759 179485
rect -960 179480 3759 179482
rect -960 179424 3698 179480
rect 3754 179424 3759 179480
rect -960 179422 3759 179424
rect -960 179332 480 179422
rect 3693 179419 3759 179422
rect 580625 170098 580691 170101
rect 583520 170098 584960 170188
rect 580625 170096 584960 170098
rect 580625 170040 580630 170096
rect 580686 170040 584960 170096
rect 580625 170038 584960 170040
rect 580625 170035 580691 170038
rect 583520 169948 584960 170038
rect -960 165066 480 165156
rect 3325 165066 3391 165069
rect -960 165064 3391 165066
rect -960 165008 3330 165064
rect 3386 165008 3391 165064
rect -960 165006 3391 165008
rect -960 164916 480 165006
rect 3325 165003 3391 165006
rect 579613 158402 579679 158405
rect 583520 158402 584960 158492
rect 579613 158400 584960 158402
rect 579613 158344 579618 158400
rect 579674 158344 584960 158400
rect 579613 158342 584960 158344
rect 579613 158339 579679 158342
rect 583520 158252 584960 158342
rect -960 150786 480 150876
rect 3877 150786 3943 150789
rect -960 150784 3943 150786
rect -960 150728 3882 150784
rect 3938 150728 3943 150784
rect -960 150726 3943 150728
rect -960 150636 480 150726
rect 3877 150723 3943 150726
rect 583520 146556 584960 146796
rect -960 136370 480 136460
rect 3325 136370 3391 136373
rect -960 136368 3391 136370
rect -960 136312 3330 136368
rect 3386 136312 3391 136368
rect -960 136310 3391 136312
rect -960 136220 480 136310
rect 3325 136307 3391 136310
rect 580165 134874 580231 134877
rect 583520 134874 584960 134964
rect 580165 134872 584960 134874
rect 580165 134816 580170 134872
rect 580226 134816 584960 134872
rect 580165 134814 584960 134816
rect 580165 134811 580231 134814
rect 583520 134724 584960 134814
rect 580349 123178 580415 123181
rect 583520 123178 584960 123268
rect 580349 123176 584960 123178
rect 580349 123120 580354 123176
rect 580410 123120 584960 123176
rect 580349 123118 584960 123120
rect 580349 123115 580415 123118
rect 583520 123028 584960 123118
rect -960 122090 480 122180
rect 3325 122090 3391 122093
rect -960 122088 3391 122090
rect -960 122032 3330 122088
rect 3386 122032 3391 122088
rect -960 122030 3391 122032
rect -960 121940 480 122030
rect 3325 122027 3391 122030
rect 580165 111482 580231 111485
rect 583520 111482 584960 111572
rect 580165 111480 584960 111482
rect 580165 111424 580170 111480
rect 580226 111424 584960 111480
rect 580165 111422 584960 111424
rect 580165 111419 580231 111422
rect 583520 111332 584960 111422
rect -960 107674 480 107764
rect 2773 107674 2839 107677
rect -960 107672 2839 107674
rect -960 107616 2778 107672
rect 2834 107616 2839 107672
rect -960 107614 2839 107616
rect -960 107524 480 107614
rect 2773 107611 2839 107614
rect 583520 99636 584960 99876
rect -960 93258 480 93348
rect 3601 93258 3667 93261
rect -960 93256 3667 93258
rect -960 93200 3606 93256
rect 3662 93200 3667 93256
rect -960 93198 3667 93200
rect -960 93108 480 93198
rect 3601 93195 3667 93198
rect 579889 87954 579955 87957
rect 583520 87954 584960 88044
rect 579889 87952 584960 87954
rect 579889 87896 579894 87952
rect 579950 87896 584960 87952
rect 579889 87894 584960 87896
rect 579889 87891 579955 87894
rect 583520 87804 584960 87894
rect -960 78978 480 79068
rect 3049 78978 3115 78981
rect -960 78976 3115 78978
rect -960 78920 3054 78976
rect 3110 78920 3115 78976
rect -960 78918 3115 78920
rect -960 78828 480 78918
rect 3049 78915 3115 78918
rect 580257 76258 580323 76261
rect 583520 76258 584960 76348
rect 580257 76256 584960 76258
rect 580257 76200 580262 76256
rect 580318 76200 584960 76256
rect 580257 76198 584960 76200
rect 580257 76195 580323 76198
rect 583520 76108 584960 76198
rect -960 64562 480 64652
rect 3509 64562 3575 64565
rect -960 64560 3575 64562
rect -960 64504 3514 64560
rect 3570 64504 3575 64560
rect -960 64502 3575 64504
rect -960 64412 480 64502
rect 3509 64499 3575 64502
rect 579797 64562 579863 64565
rect 583520 64562 584960 64652
rect 579797 64560 584960 64562
rect 579797 64504 579802 64560
rect 579858 64504 584960 64560
rect 579797 64502 584960 64504
rect 579797 64499 579863 64502
rect 583520 64412 584960 64502
rect 583520 52716 584960 52956
rect -960 50146 480 50236
rect 3417 50146 3483 50149
rect -960 50144 3483 50146
rect -960 50088 3422 50144
rect 3478 50088 3483 50144
rect -960 50086 3483 50088
rect -960 49996 480 50086
rect 3417 50083 3483 50086
rect 580165 41034 580231 41037
rect 583520 41034 584960 41124
rect 580165 41032 584960 41034
rect 580165 40976 580170 41032
rect 580226 40976 584960 41032
rect 580165 40974 584960 40976
rect 580165 40971 580231 40974
rect 583520 40884 584960 40974
rect -960 35866 480 35956
rect 3417 35866 3483 35869
rect -960 35864 3483 35866
rect -960 35808 3422 35864
rect 3478 35808 3483 35864
rect -960 35806 3483 35808
rect -960 35716 480 35806
rect 3417 35803 3483 35806
rect 579613 29338 579679 29341
rect 583520 29338 584960 29428
rect 579613 29336 584960 29338
rect 579613 29280 579618 29336
rect 579674 29280 584960 29336
rect 579613 29278 584960 29280
rect 579613 29275 579679 29278
rect 583520 29188 584960 29278
rect -960 21450 480 21540
rect 2773 21450 2839 21453
rect -960 21448 2839 21450
rect -960 21392 2778 21448
rect 2834 21392 2839 21448
rect -960 21390 2839 21392
rect -960 21300 480 21390
rect 2773 21387 2839 21390
rect 580165 17642 580231 17645
rect 583520 17642 584960 17732
rect 580165 17640 584960 17642
rect 580165 17584 580170 17640
rect 580226 17584 584960 17640
rect 580165 17582 584960 17584
rect 580165 17579 580231 17582
rect 583520 17492 584960 17582
rect -960 7170 480 7260
rect 3141 7170 3207 7173
rect -960 7168 3207 7170
rect -960 7112 3146 7168
rect 3202 7112 3207 7168
rect -960 7110 3207 7112
rect -960 7020 480 7110
rect 3141 7107 3207 7110
rect 18804 6016 19404 6017
rect 18804 5952 18832 6016
rect 18896 5952 18912 6016
rect 18976 5952 18992 6016
rect 19056 5952 19072 6016
rect 19136 5952 19152 6016
rect 19216 5952 19232 6016
rect 19296 5952 19312 6016
rect 19376 5952 19404 6016
rect 18804 5951 19404 5952
rect 54804 6016 55404 6017
rect 54804 5952 54832 6016
rect 54896 5952 54912 6016
rect 54976 5952 54992 6016
rect 55056 5952 55072 6016
rect 55136 5952 55152 6016
rect 55216 5952 55232 6016
rect 55296 5952 55312 6016
rect 55376 5952 55404 6016
rect 54804 5951 55404 5952
rect 90804 6016 91404 6017
rect 90804 5952 90832 6016
rect 90896 5952 90912 6016
rect 90976 5952 90992 6016
rect 91056 5952 91072 6016
rect 91136 5952 91152 6016
rect 91216 5952 91232 6016
rect 91296 5952 91312 6016
rect 91376 5952 91404 6016
rect 90804 5951 91404 5952
rect 126804 6016 127404 6017
rect 126804 5952 126832 6016
rect 126896 5952 126912 6016
rect 126976 5952 126992 6016
rect 127056 5952 127072 6016
rect 127136 5952 127152 6016
rect 127216 5952 127232 6016
rect 127296 5952 127312 6016
rect 127376 5952 127404 6016
rect 126804 5951 127404 5952
rect 162804 6016 163404 6017
rect 162804 5952 162832 6016
rect 162896 5952 162912 6016
rect 162976 5952 162992 6016
rect 163056 5952 163072 6016
rect 163136 5952 163152 6016
rect 163216 5952 163232 6016
rect 163296 5952 163312 6016
rect 163376 5952 163404 6016
rect 162804 5951 163404 5952
rect 198804 6016 199404 6017
rect 198804 5952 198832 6016
rect 198896 5952 198912 6016
rect 198976 5952 198992 6016
rect 199056 5952 199072 6016
rect 199136 5952 199152 6016
rect 199216 5952 199232 6016
rect 199296 5952 199312 6016
rect 199376 5952 199404 6016
rect 198804 5951 199404 5952
rect 234804 6016 235404 6017
rect 234804 5952 234832 6016
rect 234896 5952 234912 6016
rect 234976 5952 234992 6016
rect 235056 5952 235072 6016
rect 235136 5952 235152 6016
rect 235216 5952 235232 6016
rect 235296 5952 235312 6016
rect 235376 5952 235404 6016
rect 234804 5951 235404 5952
rect 270804 6016 271404 6017
rect 270804 5952 270832 6016
rect 270896 5952 270912 6016
rect 270976 5952 270992 6016
rect 271056 5952 271072 6016
rect 271136 5952 271152 6016
rect 271216 5952 271232 6016
rect 271296 5952 271312 6016
rect 271376 5952 271404 6016
rect 270804 5951 271404 5952
rect 306804 6016 307404 6017
rect 306804 5952 306832 6016
rect 306896 5952 306912 6016
rect 306976 5952 306992 6016
rect 307056 5952 307072 6016
rect 307136 5952 307152 6016
rect 307216 5952 307232 6016
rect 307296 5952 307312 6016
rect 307376 5952 307404 6016
rect 306804 5951 307404 5952
rect 342804 6016 343404 6017
rect 342804 5952 342832 6016
rect 342896 5952 342912 6016
rect 342976 5952 342992 6016
rect 343056 5952 343072 6016
rect 343136 5952 343152 6016
rect 343216 5952 343232 6016
rect 343296 5952 343312 6016
rect 343376 5952 343404 6016
rect 342804 5951 343404 5952
rect 378804 6016 379404 6017
rect 378804 5952 378832 6016
rect 378896 5952 378912 6016
rect 378976 5952 378992 6016
rect 379056 5952 379072 6016
rect 379136 5952 379152 6016
rect 379216 5952 379232 6016
rect 379296 5952 379312 6016
rect 379376 5952 379404 6016
rect 378804 5951 379404 5952
rect 414804 6016 415404 6017
rect 414804 5952 414832 6016
rect 414896 5952 414912 6016
rect 414976 5952 414992 6016
rect 415056 5952 415072 6016
rect 415136 5952 415152 6016
rect 415216 5952 415232 6016
rect 415296 5952 415312 6016
rect 415376 5952 415404 6016
rect 414804 5951 415404 5952
rect 450804 6016 451404 6017
rect 450804 5952 450832 6016
rect 450896 5952 450912 6016
rect 450976 5952 450992 6016
rect 451056 5952 451072 6016
rect 451136 5952 451152 6016
rect 451216 5952 451232 6016
rect 451296 5952 451312 6016
rect 451376 5952 451404 6016
rect 450804 5951 451404 5952
rect 486804 6016 487404 6017
rect 486804 5952 486832 6016
rect 486896 5952 486912 6016
rect 486976 5952 486992 6016
rect 487056 5952 487072 6016
rect 487136 5952 487152 6016
rect 487216 5952 487232 6016
rect 487296 5952 487312 6016
rect 487376 5952 487404 6016
rect 486804 5951 487404 5952
rect 522804 6016 523404 6017
rect 522804 5952 522832 6016
rect 522896 5952 522912 6016
rect 522976 5952 522992 6016
rect 523056 5952 523072 6016
rect 523136 5952 523152 6016
rect 523216 5952 523232 6016
rect 523296 5952 523312 6016
rect 523376 5952 523404 6016
rect 522804 5951 523404 5952
rect 558804 6016 559404 6017
rect 558804 5952 558832 6016
rect 558896 5952 558912 6016
rect 558976 5952 558992 6016
rect 559056 5952 559072 6016
rect 559136 5952 559152 6016
rect 559216 5952 559232 6016
rect 559296 5952 559312 6016
rect 559376 5952 559404 6016
rect 558804 5951 559404 5952
rect 583520 5796 584960 6036
rect 36804 5472 37404 5473
rect 36804 5408 36832 5472
rect 36896 5408 36912 5472
rect 36976 5408 36992 5472
rect 37056 5408 37072 5472
rect 37136 5408 37152 5472
rect 37216 5408 37232 5472
rect 37296 5408 37312 5472
rect 37376 5408 37404 5472
rect 36804 5407 37404 5408
rect 72804 5472 73404 5473
rect 72804 5408 72832 5472
rect 72896 5408 72912 5472
rect 72976 5408 72992 5472
rect 73056 5408 73072 5472
rect 73136 5408 73152 5472
rect 73216 5408 73232 5472
rect 73296 5408 73312 5472
rect 73376 5408 73404 5472
rect 72804 5407 73404 5408
rect 108804 5472 109404 5473
rect 108804 5408 108832 5472
rect 108896 5408 108912 5472
rect 108976 5408 108992 5472
rect 109056 5408 109072 5472
rect 109136 5408 109152 5472
rect 109216 5408 109232 5472
rect 109296 5408 109312 5472
rect 109376 5408 109404 5472
rect 108804 5407 109404 5408
rect 144804 5472 145404 5473
rect 144804 5408 144832 5472
rect 144896 5408 144912 5472
rect 144976 5408 144992 5472
rect 145056 5408 145072 5472
rect 145136 5408 145152 5472
rect 145216 5408 145232 5472
rect 145296 5408 145312 5472
rect 145376 5408 145404 5472
rect 144804 5407 145404 5408
rect 180804 5472 181404 5473
rect 180804 5408 180832 5472
rect 180896 5408 180912 5472
rect 180976 5408 180992 5472
rect 181056 5408 181072 5472
rect 181136 5408 181152 5472
rect 181216 5408 181232 5472
rect 181296 5408 181312 5472
rect 181376 5408 181404 5472
rect 180804 5407 181404 5408
rect 216804 5472 217404 5473
rect 216804 5408 216832 5472
rect 216896 5408 216912 5472
rect 216976 5408 216992 5472
rect 217056 5408 217072 5472
rect 217136 5408 217152 5472
rect 217216 5408 217232 5472
rect 217296 5408 217312 5472
rect 217376 5408 217404 5472
rect 216804 5407 217404 5408
rect 252804 5472 253404 5473
rect 252804 5408 252832 5472
rect 252896 5408 252912 5472
rect 252976 5408 252992 5472
rect 253056 5408 253072 5472
rect 253136 5408 253152 5472
rect 253216 5408 253232 5472
rect 253296 5408 253312 5472
rect 253376 5408 253404 5472
rect 252804 5407 253404 5408
rect 288804 5472 289404 5473
rect 288804 5408 288832 5472
rect 288896 5408 288912 5472
rect 288976 5408 288992 5472
rect 289056 5408 289072 5472
rect 289136 5408 289152 5472
rect 289216 5408 289232 5472
rect 289296 5408 289312 5472
rect 289376 5408 289404 5472
rect 288804 5407 289404 5408
rect 324804 5472 325404 5473
rect 324804 5408 324832 5472
rect 324896 5408 324912 5472
rect 324976 5408 324992 5472
rect 325056 5408 325072 5472
rect 325136 5408 325152 5472
rect 325216 5408 325232 5472
rect 325296 5408 325312 5472
rect 325376 5408 325404 5472
rect 324804 5407 325404 5408
rect 360804 5472 361404 5473
rect 360804 5408 360832 5472
rect 360896 5408 360912 5472
rect 360976 5408 360992 5472
rect 361056 5408 361072 5472
rect 361136 5408 361152 5472
rect 361216 5408 361232 5472
rect 361296 5408 361312 5472
rect 361376 5408 361404 5472
rect 360804 5407 361404 5408
rect 396804 5472 397404 5473
rect 396804 5408 396832 5472
rect 396896 5408 396912 5472
rect 396976 5408 396992 5472
rect 397056 5408 397072 5472
rect 397136 5408 397152 5472
rect 397216 5408 397232 5472
rect 397296 5408 397312 5472
rect 397376 5408 397404 5472
rect 396804 5407 397404 5408
rect 432804 5472 433404 5473
rect 432804 5408 432832 5472
rect 432896 5408 432912 5472
rect 432976 5408 432992 5472
rect 433056 5408 433072 5472
rect 433136 5408 433152 5472
rect 433216 5408 433232 5472
rect 433296 5408 433312 5472
rect 433376 5408 433404 5472
rect 432804 5407 433404 5408
rect 468804 5472 469404 5473
rect 468804 5408 468832 5472
rect 468896 5408 468912 5472
rect 468976 5408 468992 5472
rect 469056 5408 469072 5472
rect 469136 5408 469152 5472
rect 469216 5408 469232 5472
rect 469296 5408 469312 5472
rect 469376 5408 469404 5472
rect 468804 5407 469404 5408
rect 504804 5472 505404 5473
rect 504804 5408 504832 5472
rect 504896 5408 504912 5472
rect 504976 5408 504992 5472
rect 505056 5408 505072 5472
rect 505136 5408 505152 5472
rect 505216 5408 505232 5472
rect 505296 5408 505312 5472
rect 505376 5408 505404 5472
rect 504804 5407 505404 5408
rect 540804 5472 541404 5473
rect 540804 5408 540832 5472
rect 540896 5408 540912 5472
rect 540976 5408 540992 5472
rect 541056 5408 541072 5472
rect 541136 5408 541152 5472
rect 541216 5408 541232 5472
rect 541296 5408 541312 5472
rect 541376 5408 541404 5472
rect 540804 5407 541404 5408
rect 576804 5472 577404 5473
rect 576804 5408 576832 5472
rect 576896 5408 576912 5472
rect 576976 5408 576992 5472
rect 577056 5408 577072 5472
rect 577136 5408 577152 5472
rect 577216 5408 577232 5472
rect 577296 5408 577312 5472
rect 577376 5408 577404 5472
rect 576804 5407 577404 5408
rect 18804 4928 19404 4929
rect 18804 4864 18832 4928
rect 18896 4864 18912 4928
rect 18976 4864 18992 4928
rect 19056 4864 19072 4928
rect 19136 4864 19152 4928
rect 19216 4864 19232 4928
rect 19296 4864 19312 4928
rect 19376 4864 19404 4928
rect 18804 4863 19404 4864
rect 54804 4928 55404 4929
rect 54804 4864 54832 4928
rect 54896 4864 54912 4928
rect 54976 4864 54992 4928
rect 55056 4864 55072 4928
rect 55136 4864 55152 4928
rect 55216 4864 55232 4928
rect 55296 4864 55312 4928
rect 55376 4864 55404 4928
rect 54804 4863 55404 4864
rect 90804 4928 91404 4929
rect 90804 4864 90832 4928
rect 90896 4864 90912 4928
rect 90976 4864 90992 4928
rect 91056 4864 91072 4928
rect 91136 4864 91152 4928
rect 91216 4864 91232 4928
rect 91296 4864 91312 4928
rect 91376 4864 91404 4928
rect 90804 4863 91404 4864
rect 126804 4928 127404 4929
rect 126804 4864 126832 4928
rect 126896 4864 126912 4928
rect 126976 4864 126992 4928
rect 127056 4864 127072 4928
rect 127136 4864 127152 4928
rect 127216 4864 127232 4928
rect 127296 4864 127312 4928
rect 127376 4864 127404 4928
rect 126804 4863 127404 4864
rect 162804 4928 163404 4929
rect 162804 4864 162832 4928
rect 162896 4864 162912 4928
rect 162976 4864 162992 4928
rect 163056 4864 163072 4928
rect 163136 4864 163152 4928
rect 163216 4864 163232 4928
rect 163296 4864 163312 4928
rect 163376 4864 163404 4928
rect 162804 4863 163404 4864
rect 198804 4928 199404 4929
rect 198804 4864 198832 4928
rect 198896 4864 198912 4928
rect 198976 4864 198992 4928
rect 199056 4864 199072 4928
rect 199136 4864 199152 4928
rect 199216 4864 199232 4928
rect 199296 4864 199312 4928
rect 199376 4864 199404 4928
rect 198804 4863 199404 4864
rect 234804 4928 235404 4929
rect 234804 4864 234832 4928
rect 234896 4864 234912 4928
rect 234976 4864 234992 4928
rect 235056 4864 235072 4928
rect 235136 4864 235152 4928
rect 235216 4864 235232 4928
rect 235296 4864 235312 4928
rect 235376 4864 235404 4928
rect 234804 4863 235404 4864
rect 270804 4928 271404 4929
rect 270804 4864 270832 4928
rect 270896 4864 270912 4928
rect 270976 4864 270992 4928
rect 271056 4864 271072 4928
rect 271136 4864 271152 4928
rect 271216 4864 271232 4928
rect 271296 4864 271312 4928
rect 271376 4864 271404 4928
rect 270804 4863 271404 4864
rect 306804 4928 307404 4929
rect 306804 4864 306832 4928
rect 306896 4864 306912 4928
rect 306976 4864 306992 4928
rect 307056 4864 307072 4928
rect 307136 4864 307152 4928
rect 307216 4864 307232 4928
rect 307296 4864 307312 4928
rect 307376 4864 307404 4928
rect 306804 4863 307404 4864
rect 342804 4928 343404 4929
rect 342804 4864 342832 4928
rect 342896 4864 342912 4928
rect 342976 4864 342992 4928
rect 343056 4864 343072 4928
rect 343136 4864 343152 4928
rect 343216 4864 343232 4928
rect 343296 4864 343312 4928
rect 343376 4864 343404 4928
rect 342804 4863 343404 4864
rect 378804 4928 379404 4929
rect 378804 4864 378832 4928
rect 378896 4864 378912 4928
rect 378976 4864 378992 4928
rect 379056 4864 379072 4928
rect 379136 4864 379152 4928
rect 379216 4864 379232 4928
rect 379296 4864 379312 4928
rect 379376 4864 379404 4928
rect 378804 4863 379404 4864
rect 414804 4928 415404 4929
rect 414804 4864 414832 4928
rect 414896 4864 414912 4928
rect 414976 4864 414992 4928
rect 415056 4864 415072 4928
rect 415136 4864 415152 4928
rect 415216 4864 415232 4928
rect 415296 4864 415312 4928
rect 415376 4864 415404 4928
rect 414804 4863 415404 4864
rect 450804 4928 451404 4929
rect 450804 4864 450832 4928
rect 450896 4864 450912 4928
rect 450976 4864 450992 4928
rect 451056 4864 451072 4928
rect 451136 4864 451152 4928
rect 451216 4864 451232 4928
rect 451296 4864 451312 4928
rect 451376 4864 451404 4928
rect 450804 4863 451404 4864
rect 486804 4928 487404 4929
rect 486804 4864 486832 4928
rect 486896 4864 486912 4928
rect 486976 4864 486992 4928
rect 487056 4864 487072 4928
rect 487136 4864 487152 4928
rect 487216 4864 487232 4928
rect 487296 4864 487312 4928
rect 487376 4864 487404 4928
rect 486804 4863 487404 4864
rect 522804 4928 523404 4929
rect 522804 4864 522832 4928
rect 522896 4864 522912 4928
rect 522976 4864 522992 4928
rect 523056 4864 523072 4928
rect 523136 4864 523152 4928
rect 523216 4864 523232 4928
rect 523296 4864 523312 4928
rect 523376 4864 523404 4928
rect 522804 4863 523404 4864
rect 558804 4928 559404 4929
rect 558804 4864 558832 4928
rect 558896 4864 558912 4928
rect 558976 4864 558992 4928
rect 559056 4864 559072 4928
rect 559136 4864 559152 4928
rect 559216 4864 559232 4928
rect 559296 4864 559312 4928
rect 559376 4864 559404 4928
rect 558804 4863 559404 4864
rect 36804 4384 37404 4385
rect 36804 4320 36832 4384
rect 36896 4320 36912 4384
rect 36976 4320 36992 4384
rect 37056 4320 37072 4384
rect 37136 4320 37152 4384
rect 37216 4320 37232 4384
rect 37296 4320 37312 4384
rect 37376 4320 37404 4384
rect 36804 4319 37404 4320
rect 72804 4384 73404 4385
rect 72804 4320 72832 4384
rect 72896 4320 72912 4384
rect 72976 4320 72992 4384
rect 73056 4320 73072 4384
rect 73136 4320 73152 4384
rect 73216 4320 73232 4384
rect 73296 4320 73312 4384
rect 73376 4320 73404 4384
rect 72804 4319 73404 4320
rect 108804 4384 109404 4385
rect 108804 4320 108832 4384
rect 108896 4320 108912 4384
rect 108976 4320 108992 4384
rect 109056 4320 109072 4384
rect 109136 4320 109152 4384
rect 109216 4320 109232 4384
rect 109296 4320 109312 4384
rect 109376 4320 109404 4384
rect 108804 4319 109404 4320
rect 144804 4384 145404 4385
rect 144804 4320 144832 4384
rect 144896 4320 144912 4384
rect 144976 4320 144992 4384
rect 145056 4320 145072 4384
rect 145136 4320 145152 4384
rect 145216 4320 145232 4384
rect 145296 4320 145312 4384
rect 145376 4320 145404 4384
rect 144804 4319 145404 4320
rect 180804 4384 181404 4385
rect 180804 4320 180832 4384
rect 180896 4320 180912 4384
rect 180976 4320 180992 4384
rect 181056 4320 181072 4384
rect 181136 4320 181152 4384
rect 181216 4320 181232 4384
rect 181296 4320 181312 4384
rect 181376 4320 181404 4384
rect 180804 4319 181404 4320
rect 216804 4384 217404 4385
rect 216804 4320 216832 4384
rect 216896 4320 216912 4384
rect 216976 4320 216992 4384
rect 217056 4320 217072 4384
rect 217136 4320 217152 4384
rect 217216 4320 217232 4384
rect 217296 4320 217312 4384
rect 217376 4320 217404 4384
rect 216804 4319 217404 4320
rect 252804 4384 253404 4385
rect 252804 4320 252832 4384
rect 252896 4320 252912 4384
rect 252976 4320 252992 4384
rect 253056 4320 253072 4384
rect 253136 4320 253152 4384
rect 253216 4320 253232 4384
rect 253296 4320 253312 4384
rect 253376 4320 253404 4384
rect 252804 4319 253404 4320
rect 288804 4384 289404 4385
rect 288804 4320 288832 4384
rect 288896 4320 288912 4384
rect 288976 4320 288992 4384
rect 289056 4320 289072 4384
rect 289136 4320 289152 4384
rect 289216 4320 289232 4384
rect 289296 4320 289312 4384
rect 289376 4320 289404 4384
rect 288804 4319 289404 4320
rect 324804 4384 325404 4385
rect 324804 4320 324832 4384
rect 324896 4320 324912 4384
rect 324976 4320 324992 4384
rect 325056 4320 325072 4384
rect 325136 4320 325152 4384
rect 325216 4320 325232 4384
rect 325296 4320 325312 4384
rect 325376 4320 325404 4384
rect 324804 4319 325404 4320
rect 360804 4384 361404 4385
rect 360804 4320 360832 4384
rect 360896 4320 360912 4384
rect 360976 4320 360992 4384
rect 361056 4320 361072 4384
rect 361136 4320 361152 4384
rect 361216 4320 361232 4384
rect 361296 4320 361312 4384
rect 361376 4320 361404 4384
rect 360804 4319 361404 4320
rect 396804 4384 397404 4385
rect 396804 4320 396832 4384
rect 396896 4320 396912 4384
rect 396976 4320 396992 4384
rect 397056 4320 397072 4384
rect 397136 4320 397152 4384
rect 397216 4320 397232 4384
rect 397296 4320 397312 4384
rect 397376 4320 397404 4384
rect 396804 4319 397404 4320
rect 432804 4384 433404 4385
rect 432804 4320 432832 4384
rect 432896 4320 432912 4384
rect 432976 4320 432992 4384
rect 433056 4320 433072 4384
rect 433136 4320 433152 4384
rect 433216 4320 433232 4384
rect 433296 4320 433312 4384
rect 433376 4320 433404 4384
rect 432804 4319 433404 4320
rect 468804 4384 469404 4385
rect 468804 4320 468832 4384
rect 468896 4320 468912 4384
rect 468976 4320 468992 4384
rect 469056 4320 469072 4384
rect 469136 4320 469152 4384
rect 469216 4320 469232 4384
rect 469296 4320 469312 4384
rect 469376 4320 469404 4384
rect 468804 4319 469404 4320
rect 504804 4384 505404 4385
rect 504804 4320 504832 4384
rect 504896 4320 504912 4384
rect 504976 4320 504992 4384
rect 505056 4320 505072 4384
rect 505136 4320 505152 4384
rect 505216 4320 505232 4384
rect 505296 4320 505312 4384
rect 505376 4320 505404 4384
rect 504804 4319 505404 4320
rect 540804 4384 541404 4385
rect 540804 4320 540832 4384
rect 540896 4320 540912 4384
rect 540976 4320 540992 4384
rect 541056 4320 541072 4384
rect 541136 4320 541152 4384
rect 541216 4320 541232 4384
rect 541296 4320 541312 4384
rect 541376 4320 541404 4384
rect 540804 4319 541404 4320
rect 576804 4384 577404 4385
rect 576804 4320 576832 4384
rect 576896 4320 576912 4384
rect 576976 4320 576992 4384
rect 577056 4320 577072 4384
rect 577136 4320 577152 4384
rect 577216 4320 577232 4384
rect 577296 4320 577312 4384
rect 577376 4320 577404 4384
rect 576804 4319 577404 4320
rect 18804 3840 19404 3841
rect 18804 3776 18832 3840
rect 18896 3776 18912 3840
rect 18976 3776 18992 3840
rect 19056 3776 19072 3840
rect 19136 3776 19152 3840
rect 19216 3776 19232 3840
rect 19296 3776 19312 3840
rect 19376 3776 19404 3840
rect 18804 3775 19404 3776
rect 54804 3840 55404 3841
rect 54804 3776 54832 3840
rect 54896 3776 54912 3840
rect 54976 3776 54992 3840
rect 55056 3776 55072 3840
rect 55136 3776 55152 3840
rect 55216 3776 55232 3840
rect 55296 3776 55312 3840
rect 55376 3776 55404 3840
rect 54804 3775 55404 3776
rect 90804 3840 91404 3841
rect 90804 3776 90832 3840
rect 90896 3776 90912 3840
rect 90976 3776 90992 3840
rect 91056 3776 91072 3840
rect 91136 3776 91152 3840
rect 91216 3776 91232 3840
rect 91296 3776 91312 3840
rect 91376 3776 91404 3840
rect 90804 3775 91404 3776
rect 126804 3840 127404 3841
rect 126804 3776 126832 3840
rect 126896 3776 126912 3840
rect 126976 3776 126992 3840
rect 127056 3776 127072 3840
rect 127136 3776 127152 3840
rect 127216 3776 127232 3840
rect 127296 3776 127312 3840
rect 127376 3776 127404 3840
rect 126804 3775 127404 3776
rect 162804 3840 163404 3841
rect 162804 3776 162832 3840
rect 162896 3776 162912 3840
rect 162976 3776 162992 3840
rect 163056 3776 163072 3840
rect 163136 3776 163152 3840
rect 163216 3776 163232 3840
rect 163296 3776 163312 3840
rect 163376 3776 163404 3840
rect 162804 3775 163404 3776
rect 198804 3840 199404 3841
rect 198804 3776 198832 3840
rect 198896 3776 198912 3840
rect 198976 3776 198992 3840
rect 199056 3776 199072 3840
rect 199136 3776 199152 3840
rect 199216 3776 199232 3840
rect 199296 3776 199312 3840
rect 199376 3776 199404 3840
rect 198804 3775 199404 3776
rect 234804 3840 235404 3841
rect 234804 3776 234832 3840
rect 234896 3776 234912 3840
rect 234976 3776 234992 3840
rect 235056 3776 235072 3840
rect 235136 3776 235152 3840
rect 235216 3776 235232 3840
rect 235296 3776 235312 3840
rect 235376 3776 235404 3840
rect 234804 3775 235404 3776
rect 270804 3840 271404 3841
rect 270804 3776 270832 3840
rect 270896 3776 270912 3840
rect 270976 3776 270992 3840
rect 271056 3776 271072 3840
rect 271136 3776 271152 3840
rect 271216 3776 271232 3840
rect 271296 3776 271312 3840
rect 271376 3776 271404 3840
rect 270804 3775 271404 3776
rect 306804 3840 307404 3841
rect 306804 3776 306832 3840
rect 306896 3776 306912 3840
rect 306976 3776 306992 3840
rect 307056 3776 307072 3840
rect 307136 3776 307152 3840
rect 307216 3776 307232 3840
rect 307296 3776 307312 3840
rect 307376 3776 307404 3840
rect 306804 3775 307404 3776
rect 342804 3840 343404 3841
rect 342804 3776 342832 3840
rect 342896 3776 342912 3840
rect 342976 3776 342992 3840
rect 343056 3776 343072 3840
rect 343136 3776 343152 3840
rect 343216 3776 343232 3840
rect 343296 3776 343312 3840
rect 343376 3776 343404 3840
rect 342804 3775 343404 3776
rect 378804 3840 379404 3841
rect 378804 3776 378832 3840
rect 378896 3776 378912 3840
rect 378976 3776 378992 3840
rect 379056 3776 379072 3840
rect 379136 3776 379152 3840
rect 379216 3776 379232 3840
rect 379296 3776 379312 3840
rect 379376 3776 379404 3840
rect 378804 3775 379404 3776
rect 414804 3840 415404 3841
rect 414804 3776 414832 3840
rect 414896 3776 414912 3840
rect 414976 3776 414992 3840
rect 415056 3776 415072 3840
rect 415136 3776 415152 3840
rect 415216 3776 415232 3840
rect 415296 3776 415312 3840
rect 415376 3776 415404 3840
rect 414804 3775 415404 3776
rect 450804 3840 451404 3841
rect 450804 3776 450832 3840
rect 450896 3776 450912 3840
rect 450976 3776 450992 3840
rect 451056 3776 451072 3840
rect 451136 3776 451152 3840
rect 451216 3776 451232 3840
rect 451296 3776 451312 3840
rect 451376 3776 451404 3840
rect 450804 3775 451404 3776
rect 486804 3840 487404 3841
rect 486804 3776 486832 3840
rect 486896 3776 486912 3840
rect 486976 3776 486992 3840
rect 487056 3776 487072 3840
rect 487136 3776 487152 3840
rect 487216 3776 487232 3840
rect 487296 3776 487312 3840
rect 487376 3776 487404 3840
rect 486804 3775 487404 3776
rect 522804 3840 523404 3841
rect 522804 3776 522832 3840
rect 522896 3776 522912 3840
rect 522976 3776 522992 3840
rect 523056 3776 523072 3840
rect 523136 3776 523152 3840
rect 523216 3776 523232 3840
rect 523296 3776 523312 3840
rect 523376 3776 523404 3840
rect 522804 3775 523404 3776
rect 558804 3840 559404 3841
rect 558804 3776 558832 3840
rect 558896 3776 558912 3840
rect 558976 3776 558992 3840
rect 559056 3776 559072 3840
rect 559136 3776 559152 3840
rect 559216 3776 559232 3840
rect 559296 3776 559312 3840
rect 559376 3776 559404 3840
rect 558804 3775 559404 3776
rect 561673 3498 561739 3501
rect 564525 3498 564591 3501
rect 561673 3496 564591 3498
rect 561673 3440 561678 3496
rect 561734 3440 564530 3496
rect 564586 3440 564591 3496
rect 561673 3438 564591 3440
rect 561673 3435 561739 3438
rect 564525 3435 564591 3438
rect 36804 3296 37404 3297
rect 36804 3232 36832 3296
rect 36896 3232 36912 3296
rect 36976 3232 36992 3296
rect 37056 3232 37072 3296
rect 37136 3232 37152 3296
rect 37216 3232 37232 3296
rect 37296 3232 37312 3296
rect 37376 3232 37404 3296
rect 36804 3231 37404 3232
rect 72804 3296 73404 3297
rect 72804 3232 72832 3296
rect 72896 3232 72912 3296
rect 72976 3232 72992 3296
rect 73056 3232 73072 3296
rect 73136 3232 73152 3296
rect 73216 3232 73232 3296
rect 73296 3232 73312 3296
rect 73376 3232 73404 3296
rect 72804 3231 73404 3232
rect 108804 3296 109404 3297
rect 108804 3232 108832 3296
rect 108896 3232 108912 3296
rect 108976 3232 108992 3296
rect 109056 3232 109072 3296
rect 109136 3232 109152 3296
rect 109216 3232 109232 3296
rect 109296 3232 109312 3296
rect 109376 3232 109404 3296
rect 108804 3231 109404 3232
rect 144804 3296 145404 3297
rect 144804 3232 144832 3296
rect 144896 3232 144912 3296
rect 144976 3232 144992 3296
rect 145056 3232 145072 3296
rect 145136 3232 145152 3296
rect 145216 3232 145232 3296
rect 145296 3232 145312 3296
rect 145376 3232 145404 3296
rect 144804 3231 145404 3232
rect 180804 3296 181404 3297
rect 180804 3232 180832 3296
rect 180896 3232 180912 3296
rect 180976 3232 180992 3296
rect 181056 3232 181072 3296
rect 181136 3232 181152 3296
rect 181216 3232 181232 3296
rect 181296 3232 181312 3296
rect 181376 3232 181404 3296
rect 180804 3231 181404 3232
rect 216804 3296 217404 3297
rect 216804 3232 216832 3296
rect 216896 3232 216912 3296
rect 216976 3232 216992 3296
rect 217056 3232 217072 3296
rect 217136 3232 217152 3296
rect 217216 3232 217232 3296
rect 217296 3232 217312 3296
rect 217376 3232 217404 3296
rect 216804 3231 217404 3232
rect 252804 3296 253404 3297
rect 252804 3232 252832 3296
rect 252896 3232 252912 3296
rect 252976 3232 252992 3296
rect 253056 3232 253072 3296
rect 253136 3232 253152 3296
rect 253216 3232 253232 3296
rect 253296 3232 253312 3296
rect 253376 3232 253404 3296
rect 252804 3231 253404 3232
rect 288804 3296 289404 3297
rect 288804 3232 288832 3296
rect 288896 3232 288912 3296
rect 288976 3232 288992 3296
rect 289056 3232 289072 3296
rect 289136 3232 289152 3296
rect 289216 3232 289232 3296
rect 289296 3232 289312 3296
rect 289376 3232 289404 3296
rect 288804 3231 289404 3232
rect 324804 3296 325404 3297
rect 324804 3232 324832 3296
rect 324896 3232 324912 3296
rect 324976 3232 324992 3296
rect 325056 3232 325072 3296
rect 325136 3232 325152 3296
rect 325216 3232 325232 3296
rect 325296 3232 325312 3296
rect 325376 3232 325404 3296
rect 324804 3231 325404 3232
rect 360804 3296 361404 3297
rect 360804 3232 360832 3296
rect 360896 3232 360912 3296
rect 360976 3232 360992 3296
rect 361056 3232 361072 3296
rect 361136 3232 361152 3296
rect 361216 3232 361232 3296
rect 361296 3232 361312 3296
rect 361376 3232 361404 3296
rect 360804 3231 361404 3232
rect 396804 3296 397404 3297
rect 396804 3232 396832 3296
rect 396896 3232 396912 3296
rect 396976 3232 396992 3296
rect 397056 3232 397072 3296
rect 397136 3232 397152 3296
rect 397216 3232 397232 3296
rect 397296 3232 397312 3296
rect 397376 3232 397404 3296
rect 396804 3231 397404 3232
rect 432804 3296 433404 3297
rect 432804 3232 432832 3296
rect 432896 3232 432912 3296
rect 432976 3232 432992 3296
rect 433056 3232 433072 3296
rect 433136 3232 433152 3296
rect 433216 3232 433232 3296
rect 433296 3232 433312 3296
rect 433376 3232 433404 3296
rect 432804 3231 433404 3232
rect 468804 3296 469404 3297
rect 468804 3232 468832 3296
rect 468896 3232 468912 3296
rect 468976 3232 468992 3296
rect 469056 3232 469072 3296
rect 469136 3232 469152 3296
rect 469216 3232 469232 3296
rect 469296 3232 469312 3296
rect 469376 3232 469404 3296
rect 468804 3231 469404 3232
rect 504804 3296 505404 3297
rect 504804 3232 504832 3296
rect 504896 3232 504912 3296
rect 504976 3232 504992 3296
rect 505056 3232 505072 3296
rect 505136 3232 505152 3296
rect 505216 3232 505232 3296
rect 505296 3232 505312 3296
rect 505376 3232 505404 3296
rect 504804 3231 505404 3232
rect 540804 3296 541404 3297
rect 540804 3232 540832 3296
rect 540896 3232 540912 3296
rect 540976 3232 540992 3296
rect 541056 3232 541072 3296
rect 541136 3232 541152 3296
rect 541216 3232 541232 3296
rect 541296 3232 541312 3296
rect 541376 3232 541404 3296
rect 540804 3231 541404 3232
rect 576804 3296 577404 3297
rect 576804 3232 576832 3296
rect 576896 3232 576912 3296
rect 576976 3232 576992 3296
rect 577056 3232 577072 3296
rect 577136 3232 577152 3296
rect 577216 3232 577232 3296
rect 577296 3232 577312 3296
rect 577376 3232 577404 3296
rect 576804 3231 577404 3232
rect 18804 2752 19404 2753
rect 18804 2688 18832 2752
rect 18896 2688 18912 2752
rect 18976 2688 18992 2752
rect 19056 2688 19072 2752
rect 19136 2688 19152 2752
rect 19216 2688 19232 2752
rect 19296 2688 19312 2752
rect 19376 2688 19404 2752
rect 18804 2687 19404 2688
rect 54804 2752 55404 2753
rect 54804 2688 54832 2752
rect 54896 2688 54912 2752
rect 54976 2688 54992 2752
rect 55056 2688 55072 2752
rect 55136 2688 55152 2752
rect 55216 2688 55232 2752
rect 55296 2688 55312 2752
rect 55376 2688 55404 2752
rect 54804 2687 55404 2688
rect 90804 2752 91404 2753
rect 90804 2688 90832 2752
rect 90896 2688 90912 2752
rect 90976 2688 90992 2752
rect 91056 2688 91072 2752
rect 91136 2688 91152 2752
rect 91216 2688 91232 2752
rect 91296 2688 91312 2752
rect 91376 2688 91404 2752
rect 90804 2687 91404 2688
rect 126804 2752 127404 2753
rect 126804 2688 126832 2752
rect 126896 2688 126912 2752
rect 126976 2688 126992 2752
rect 127056 2688 127072 2752
rect 127136 2688 127152 2752
rect 127216 2688 127232 2752
rect 127296 2688 127312 2752
rect 127376 2688 127404 2752
rect 126804 2687 127404 2688
rect 162804 2752 163404 2753
rect 162804 2688 162832 2752
rect 162896 2688 162912 2752
rect 162976 2688 162992 2752
rect 163056 2688 163072 2752
rect 163136 2688 163152 2752
rect 163216 2688 163232 2752
rect 163296 2688 163312 2752
rect 163376 2688 163404 2752
rect 162804 2687 163404 2688
rect 198804 2752 199404 2753
rect 198804 2688 198832 2752
rect 198896 2688 198912 2752
rect 198976 2688 198992 2752
rect 199056 2688 199072 2752
rect 199136 2688 199152 2752
rect 199216 2688 199232 2752
rect 199296 2688 199312 2752
rect 199376 2688 199404 2752
rect 198804 2687 199404 2688
rect 234804 2752 235404 2753
rect 234804 2688 234832 2752
rect 234896 2688 234912 2752
rect 234976 2688 234992 2752
rect 235056 2688 235072 2752
rect 235136 2688 235152 2752
rect 235216 2688 235232 2752
rect 235296 2688 235312 2752
rect 235376 2688 235404 2752
rect 234804 2687 235404 2688
rect 270804 2752 271404 2753
rect 270804 2688 270832 2752
rect 270896 2688 270912 2752
rect 270976 2688 270992 2752
rect 271056 2688 271072 2752
rect 271136 2688 271152 2752
rect 271216 2688 271232 2752
rect 271296 2688 271312 2752
rect 271376 2688 271404 2752
rect 270804 2687 271404 2688
rect 306804 2752 307404 2753
rect 306804 2688 306832 2752
rect 306896 2688 306912 2752
rect 306976 2688 306992 2752
rect 307056 2688 307072 2752
rect 307136 2688 307152 2752
rect 307216 2688 307232 2752
rect 307296 2688 307312 2752
rect 307376 2688 307404 2752
rect 306804 2687 307404 2688
rect 342804 2752 343404 2753
rect 342804 2688 342832 2752
rect 342896 2688 342912 2752
rect 342976 2688 342992 2752
rect 343056 2688 343072 2752
rect 343136 2688 343152 2752
rect 343216 2688 343232 2752
rect 343296 2688 343312 2752
rect 343376 2688 343404 2752
rect 342804 2687 343404 2688
rect 378804 2752 379404 2753
rect 378804 2688 378832 2752
rect 378896 2688 378912 2752
rect 378976 2688 378992 2752
rect 379056 2688 379072 2752
rect 379136 2688 379152 2752
rect 379216 2688 379232 2752
rect 379296 2688 379312 2752
rect 379376 2688 379404 2752
rect 378804 2687 379404 2688
rect 414804 2752 415404 2753
rect 414804 2688 414832 2752
rect 414896 2688 414912 2752
rect 414976 2688 414992 2752
rect 415056 2688 415072 2752
rect 415136 2688 415152 2752
rect 415216 2688 415232 2752
rect 415296 2688 415312 2752
rect 415376 2688 415404 2752
rect 414804 2687 415404 2688
rect 450804 2752 451404 2753
rect 450804 2688 450832 2752
rect 450896 2688 450912 2752
rect 450976 2688 450992 2752
rect 451056 2688 451072 2752
rect 451136 2688 451152 2752
rect 451216 2688 451232 2752
rect 451296 2688 451312 2752
rect 451376 2688 451404 2752
rect 450804 2687 451404 2688
rect 486804 2752 487404 2753
rect 486804 2688 486832 2752
rect 486896 2688 486912 2752
rect 486976 2688 486992 2752
rect 487056 2688 487072 2752
rect 487136 2688 487152 2752
rect 487216 2688 487232 2752
rect 487296 2688 487312 2752
rect 487376 2688 487404 2752
rect 486804 2687 487404 2688
rect 522804 2752 523404 2753
rect 522804 2688 522832 2752
rect 522896 2688 522912 2752
rect 522976 2688 522992 2752
rect 523056 2688 523072 2752
rect 523136 2688 523152 2752
rect 523216 2688 523232 2752
rect 523296 2688 523312 2752
rect 523376 2688 523404 2752
rect 522804 2687 523404 2688
rect 558804 2752 559404 2753
rect 558804 2688 558832 2752
rect 558896 2688 558912 2752
rect 558976 2688 558992 2752
rect 559056 2688 559072 2752
rect 559136 2688 559152 2752
rect 559216 2688 559232 2752
rect 559296 2688 559312 2752
rect 559376 2688 559404 2752
rect 558804 2687 559404 2688
rect 36804 2208 37404 2209
rect 36804 2144 36832 2208
rect 36896 2144 36912 2208
rect 36976 2144 36992 2208
rect 37056 2144 37072 2208
rect 37136 2144 37152 2208
rect 37216 2144 37232 2208
rect 37296 2144 37312 2208
rect 37376 2144 37404 2208
rect 36804 2143 37404 2144
rect 72804 2208 73404 2209
rect 72804 2144 72832 2208
rect 72896 2144 72912 2208
rect 72976 2144 72992 2208
rect 73056 2144 73072 2208
rect 73136 2144 73152 2208
rect 73216 2144 73232 2208
rect 73296 2144 73312 2208
rect 73376 2144 73404 2208
rect 72804 2143 73404 2144
rect 108804 2208 109404 2209
rect 108804 2144 108832 2208
rect 108896 2144 108912 2208
rect 108976 2144 108992 2208
rect 109056 2144 109072 2208
rect 109136 2144 109152 2208
rect 109216 2144 109232 2208
rect 109296 2144 109312 2208
rect 109376 2144 109404 2208
rect 108804 2143 109404 2144
rect 144804 2208 145404 2209
rect 144804 2144 144832 2208
rect 144896 2144 144912 2208
rect 144976 2144 144992 2208
rect 145056 2144 145072 2208
rect 145136 2144 145152 2208
rect 145216 2144 145232 2208
rect 145296 2144 145312 2208
rect 145376 2144 145404 2208
rect 144804 2143 145404 2144
rect 180804 2208 181404 2209
rect 180804 2144 180832 2208
rect 180896 2144 180912 2208
rect 180976 2144 180992 2208
rect 181056 2144 181072 2208
rect 181136 2144 181152 2208
rect 181216 2144 181232 2208
rect 181296 2144 181312 2208
rect 181376 2144 181404 2208
rect 180804 2143 181404 2144
rect 216804 2208 217404 2209
rect 216804 2144 216832 2208
rect 216896 2144 216912 2208
rect 216976 2144 216992 2208
rect 217056 2144 217072 2208
rect 217136 2144 217152 2208
rect 217216 2144 217232 2208
rect 217296 2144 217312 2208
rect 217376 2144 217404 2208
rect 216804 2143 217404 2144
rect 252804 2208 253404 2209
rect 252804 2144 252832 2208
rect 252896 2144 252912 2208
rect 252976 2144 252992 2208
rect 253056 2144 253072 2208
rect 253136 2144 253152 2208
rect 253216 2144 253232 2208
rect 253296 2144 253312 2208
rect 253376 2144 253404 2208
rect 252804 2143 253404 2144
rect 288804 2208 289404 2209
rect 288804 2144 288832 2208
rect 288896 2144 288912 2208
rect 288976 2144 288992 2208
rect 289056 2144 289072 2208
rect 289136 2144 289152 2208
rect 289216 2144 289232 2208
rect 289296 2144 289312 2208
rect 289376 2144 289404 2208
rect 288804 2143 289404 2144
rect 324804 2208 325404 2209
rect 324804 2144 324832 2208
rect 324896 2144 324912 2208
rect 324976 2144 324992 2208
rect 325056 2144 325072 2208
rect 325136 2144 325152 2208
rect 325216 2144 325232 2208
rect 325296 2144 325312 2208
rect 325376 2144 325404 2208
rect 324804 2143 325404 2144
rect 360804 2208 361404 2209
rect 360804 2144 360832 2208
rect 360896 2144 360912 2208
rect 360976 2144 360992 2208
rect 361056 2144 361072 2208
rect 361136 2144 361152 2208
rect 361216 2144 361232 2208
rect 361296 2144 361312 2208
rect 361376 2144 361404 2208
rect 360804 2143 361404 2144
rect 396804 2208 397404 2209
rect 396804 2144 396832 2208
rect 396896 2144 396912 2208
rect 396976 2144 396992 2208
rect 397056 2144 397072 2208
rect 397136 2144 397152 2208
rect 397216 2144 397232 2208
rect 397296 2144 397312 2208
rect 397376 2144 397404 2208
rect 396804 2143 397404 2144
rect 432804 2208 433404 2209
rect 432804 2144 432832 2208
rect 432896 2144 432912 2208
rect 432976 2144 432992 2208
rect 433056 2144 433072 2208
rect 433136 2144 433152 2208
rect 433216 2144 433232 2208
rect 433296 2144 433312 2208
rect 433376 2144 433404 2208
rect 432804 2143 433404 2144
rect 468804 2208 469404 2209
rect 468804 2144 468832 2208
rect 468896 2144 468912 2208
rect 468976 2144 468992 2208
rect 469056 2144 469072 2208
rect 469136 2144 469152 2208
rect 469216 2144 469232 2208
rect 469296 2144 469312 2208
rect 469376 2144 469404 2208
rect 468804 2143 469404 2144
rect 504804 2208 505404 2209
rect 504804 2144 504832 2208
rect 504896 2144 504912 2208
rect 504976 2144 504992 2208
rect 505056 2144 505072 2208
rect 505136 2144 505152 2208
rect 505216 2144 505232 2208
rect 505296 2144 505312 2208
rect 505376 2144 505404 2208
rect 504804 2143 505404 2144
rect 540804 2208 541404 2209
rect 540804 2144 540832 2208
rect 540896 2144 540912 2208
rect 540976 2144 540992 2208
rect 541056 2144 541072 2208
rect 541136 2144 541152 2208
rect 541216 2144 541232 2208
rect 541296 2144 541312 2208
rect 541376 2144 541404 2208
rect 540804 2143 541404 2144
rect 576804 2208 577404 2209
rect 576804 2144 576832 2208
rect 576896 2144 576912 2208
rect 576976 2144 576992 2208
rect 577056 2144 577072 2208
rect 577136 2144 577152 2208
rect 577216 2144 577232 2208
rect 577296 2144 577312 2208
rect 577376 2144 577404 2208
rect 576804 2143 577404 2144
<< via3 >>
rect 36832 701788 36896 701792
rect 36832 701732 36836 701788
rect 36836 701732 36892 701788
rect 36892 701732 36896 701788
rect 36832 701728 36896 701732
rect 36912 701788 36976 701792
rect 36912 701732 36916 701788
rect 36916 701732 36972 701788
rect 36972 701732 36976 701788
rect 36912 701728 36976 701732
rect 36992 701788 37056 701792
rect 36992 701732 36996 701788
rect 36996 701732 37052 701788
rect 37052 701732 37056 701788
rect 36992 701728 37056 701732
rect 37072 701788 37136 701792
rect 37072 701732 37076 701788
rect 37076 701732 37132 701788
rect 37132 701732 37136 701788
rect 37072 701728 37136 701732
rect 37152 701788 37216 701792
rect 37152 701732 37156 701788
rect 37156 701732 37212 701788
rect 37212 701732 37216 701788
rect 37152 701728 37216 701732
rect 37232 701788 37296 701792
rect 37232 701732 37236 701788
rect 37236 701732 37292 701788
rect 37292 701732 37296 701788
rect 37232 701728 37296 701732
rect 37312 701788 37376 701792
rect 37312 701732 37316 701788
rect 37316 701732 37372 701788
rect 37372 701732 37376 701788
rect 37312 701728 37376 701732
rect 72832 701788 72896 701792
rect 72832 701732 72836 701788
rect 72836 701732 72892 701788
rect 72892 701732 72896 701788
rect 72832 701728 72896 701732
rect 72912 701788 72976 701792
rect 72912 701732 72916 701788
rect 72916 701732 72972 701788
rect 72972 701732 72976 701788
rect 72912 701728 72976 701732
rect 72992 701788 73056 701792
rect 72992 701732 72996 701788
rect 72996 701732 73052 701788
rect 73052 701732 73056 701788
rect 72992 701728 73056 701732
rect 73072 701788 73136 701792
rect 73072 701732 73076 701788
rect 73076 701732 73132 701788
rect 73132 701732 73136 701788
rect 73072 701728 73136 701732
rect 73152 701788 73216 701792
rect 73152 701732 73156 701788
rect 73156 701732 73212 701788
rect 73212 701732 73216 701788
rect 73152 701728 73216 701732
rect 73232 701788 73296 701792
rect 73232 701732 73236 701788
rect 73236 701732 73292 701788
rect 73292 701732 73296 701788
rect 73232 701728 73296 701732
rect 73312 701788 73376 701792
rect 73312 701732 73316 701788
rect 73316 701732 73372 701788
rect 73372 701732 73376 701788
rect 73312 701728 73376 701732
rect 108832 701788 108896 701792
rect 108832 701732 108836 701788
rect 108836 701732 108892 701788
rect 108892 701732 108896 701788
rect 108832 701728 108896 701732
rect 108912 701788 108976 701792
rect 108912 701732 108916 701788
rect 108916 701732 108972 701788
rect 108972 701732 108976 701788
rect 108912 701728 108976 701732
rect 108992 701788 109056 701792
rect 108992 701732 108996 701788
rect 108996 701732 109052 701788
rect 109052 701732 109056 701788
rect 108992 701728 109056 701732
rect 109072 701788 109136 701792
rect 109072 701732 109076 701788
rect 109076 701732 109132 701788
rect 109132 701732 109136 701788
rect 109072 701728 109136 701732
rect 109152 701788 109216 701792
rect 109152 701732 109156 701788
rect 109156 701732 109212 701788
rect 109212 701732 109216 701788
rect 109152 701728 109216 701732
rect 109232 701788 109296 701792
rect 109232 701732 109236 701788
rect 109236 701732 109292 701788
rect 109292 701732 109296 701788
rect 109232 701728 109296 701732
rect 109312 701788 109376 701792
rect 109312 701732 109316 701788
rect 109316 701732 109372 701788
rect 109372 701732 109376 701788
rect 109312 701728 109376 701732
rect 144832 701788 144896 701792
rect 144832 701732 144836 701788
rect 144836 701732 144892 701788
rect 144892 701732 144896 701788
rect 144832 701728 144896 701732
rect 144912 701788 144976 701792
rect 144912 701732 144916 701788
rect 144916 701732 144972 701788
rect 144972 701732 144976 701788
rect 144912 701728 144976 701732
rect 144992 701788 145056 701792
rect 144992 701732 144996 701788
rect 144996 701732 145052 701788
rect 145052 701732 145056 701788
rect 144992 701728 145056 701732
rect 145072 701788 145136 701792
rect 145072 701732 145076 701788
rect 145076 701732 145132 701788
rect 145132 701732 145136 701788
rect 145072 701728 145136 701732
rect 145152 701788 145216 701792
rect 145152 701732 145156 701788
rect 145156 701732 145212 701788
rect 145212 701732 145216 701788
rect 145152 701728 145216 701732
rect 145232 701788 145296 701792
rect 145232 701732 145236 701788
rect 145236 701732 145292 701788
rect 145292 701732 145296 701788
rect 145232 701728 145296 701732
rect 145312 701788 145376 701792
rect 145312 701732 145316 701788
rect 145316 701732 145372 701788
rect 145372 701732 145376 701788
rect 145312 701728 145376 701732
rect 180832 701788 180896 701792
rect 180832 701732 180836 701788
rect 180836 701732 180892 701788
rect 180892 701732 180896 701788
rect 180832 701728 180896 701732
rect 180912 701788 180976 701792
rect 180912 701732 180916 701788
rect 180916 701732 180972 701788
rect 180972 701732 180976 701788
rect 180912 701728 180976 701732
rect 180992 701788 181056 701792
rect 180992 701732 180996 701788
rect 180996 701732 181052 701788
rect 181052 701732 181056 701788
rect 180992 701728 181056 701732
rect 181072 701788 181136 701792
rect 181072 701732 181076 701788
rect 181076 701732 181132 701788
rect 181132 701732 181136 701788
rect 181072 701728 181136 701732
rect 181152 701788 181216 701792
rect 181152 701732 181156 701788
rect 181156 701732 181212 701788
rect 181212 701732 181216 701788
rect 181152 701728 181216 701732
rect 181232 701788 181296 701792
rect 181232 701732 181236 701788
rect 181236 701732 181292 701788
rect 181292 701732 181296 701788
rect 181232 701728 181296 701732
rect 181312 701788 181376 701792
rect 181312 701732 181316 701788
rect 181316 701732 181372 701788
rect 181372 701732 181376 701788
rect 181312 701728 181376 701732
rect 216832 701788 216896 701792
rect 216832 701732 216836 701788
rect 216836 701732 216892 701788
rect 216892 701732 216896 701788
rect 216832 701728 216896 701732
rect 216912 701788 216976 701792
rect 216912 701732 216916 701788
rect 216916 701732 216972 701788
rect 216972 701732 216976 701788
rect 216912 701728 216976 701732
rect 216992 701788 217056 701792
rect 216992 701732 216996 701788
rect 216996 701732 217052 701788
rect 217052 701732 217056 701788
rect 216992 701728 217056 701732
rect 217072 701788 217136 701792
rect 217072 701732 217076 701788
rect 217076 701732 217132 701788
rect 217132 701732 217136 701788
rect 217072 701728 217136 701732
rect 217152 701788 217216 701792
rect 217152 701732 217156 701788
rect 217156 701732 217212 701788
rect 217212 701732 217216 701788
rect 217152 701728 217216 701732
rect 217232 701788 217296 701792
rect 217232 701732 217236 701788
rect 217236 701732 217292 701788
rect 217292 701732 217296 701788
rect 217232 701728 217296 701732
rect 217312 701788 217376 701792
rect 217312 701732 217316 701788
rect 217316 701732 217372 701788
rect 217372 701732 217376 701788
rect 217312 701728 217376 701732
rect 252832 701788 252896 701792
rect 252832 701732 252836 701788
rect 252836 701732 252892 701788
rect 252892 701732 252896 701788
rect 252832 701728 252896 701732
rect 252912 701788 252976 701792
rect 252912 701732 252916 701788
rect 252916 701732 252972 701788
rect 252972 701732 252976 701788
rect 252912 701728 252976 701732
rect 252992 701788 253056 701792
rect 252992 701732 252996 701788
rect 252996 701732 253052 701788
rect 253052 701732 253056 701788
rect 252992 701728 253056 701732
rect 253072 701788 253136 701792
rect 253072 701732 253076 701788
rect 253076 701732 253132 701788
rect 253132 701732 253136 701788
rect 253072 701728 253136 701732
rect 253152 701788 253216 701792
rect 253152 701732 253156 701788
rect 253156 701732 253212 701788
rect 253212 701732 253216 701788
rect 253152 701728 253216 701732
rect 253232 701788 253296 701792
rect 253232 701732 253236 701788
rect 253236 701732 253292 701788
rect 253292 701732 253296 701788
rect 253232 701728 253296 701732
rect 253312 701788 253376 701792
rect 253312 701732 253316 701788
rect 253316 701732 253372 701788
rect 253372 701732 253376 701788
rect 253312 701728 253376 701732
rect 288832 701788 288896 701792
rect 288832 701732 288836 701788
rect 288836 701732 288892 701788
rect 288892 701732 288896 701788
rect 288832 701728 288896 701732
rect 288912 701788 288976 701792
rect 288912 701732 288916 701788
rect 288916 701732 288972 701788
rect 288972 701732 288976 701788
rect 288912 701728 288976 701732
rect 288992 701788 289056 701792
rect 288992 701732 288996 701788
rect 288996 701732 289052 701788
rect 289052 701732 289056 701788
rect 288992 701728 289056 701732
rect 289072 701788 289136 701792
rect 289072 701732 289076 701788
rect 289076 701732 289132 701788
rect 289132 701732 289136 701788
rect 289072 701728 289136 701732
rect 289152 701788 289216 701792
rect 289152 701732 289156 701788
rect 289156 701732 289212 701788
rect 289212 701732 289216 701788
rect 289152 701728 289216 701732
rect 289232 701788 289296 701792
rect 289232 701732 289236 701788
rect 289236 701732 289292 701788
rect 289292 701732 289296 701788
rect 289232 701728 289296 701732
rect 289312 701788 289376 701792
rect 289312 701732 289316 701788
rect 289316 701732 289372 701788
rect 289372 701732 289376 701788
rect 289312 701728 289376 701732
rect 324832 701788 324896 701792
rect 324832 701732 324836 701788
rect 324836 701732 324892 701788
rect 324892 701732 324896 701788
rect 324832 701728 324896 701732
rect 324912 701788 324976 701792
rect 324912 701732 324916 701788
rect 324916 701732 324972 701788
rect 324972 701732 324976 701788
rect 324912 701728 324976 701732
rect 324992 701788 325056 701792
rect 324992 701732 324996 701788
rect 324996 701732 325052 701788
rect 325052 701732 325056 701788
rect 324992 701728 325056 701732
rect 325072 701788 325136 701792
rect 325072 701732 325076 701788
rect 325076 701732 325132 701788
rect 325132 701732 325136 701788
rect 325072 701728 325136 701732
rect 325152 701788 325216 701792
rect 325152 701732 325156 701788
rect 325156 701732 325212 701788
rect 325212 701732 325216 701788
rect 325152 701728 325216 701732
rect 325232 701788 325296 701792
rect 325232 701732 325236 701788
rect 325236 701732 325292 701788
rect 325292 701732 325296 701788
rect 325232 701728 325296 701732
rect 325312 701788 325376 701792
rect 325312 701732 325316 701788
rect 325316 701732 325372 701788
rect 325372 701732 325376 701788
rect 325312 701728 325376 701732
rect 360832 701788 360896 701792
rect 360832 701732 360836 701788
rect 360836 701732 360892 701788
rect 360892 701732 360896 701788
rect 360832 701728 360896 701732
rect 360912 701788 360976 701792
rect 360912 701732 360916 701788
rect 360916 701732 360972 701788
rect 360972 701732 360976 701788
rect 360912 701728 360976 701732
rect 360992 701788 361056 701792
rect 360992 701732 360996 701788
rect 360996 701732 361052 701788
rect 361052 701732 361056 701788
rect 360992 701728 361056 701732
rect 361072 701788 361136 701792
rect 361072 701732 361076 701788
rect 361076 701732 361132 701788
rect 361132 701732 361136 701788
rect 361072 701728 361136 701732
rect 361152 701788 361216 701792
rect 361152 701732 361156 701788
rect 361156 701732 361212 701788
rect 361212 701732 361216 701788
rect 361152 701728 361216 701732
rect 361232 701788 361296 701792
rect 361232 701732 361236 701788
rect 361236 701732 361292 701788
rect 361292 701732 361296 701788
rect 361232 701728 361296 701732
rect 361312 701788 361376 701792
rect 361312 701732 361316 701788
rect 361316 701732 361372 701788
rect 361372 701732 361376 701788
rect 361312 701728 361376 701732
rect 396832 701788 396896 701792
rect 396832 701732 396836 701788
rect 396836 701732 396892 701788
rect 396892 701732 396896 701788
rect 396832 701728 396896 701732
rect 396912 701788 396976 701792
rect 396912 701732 396916 701788
rect 396916 701732 396972 701788
rect 396972 701732 396976 701788
rect 396912 701728 396976 701732
rect 396992 701788 397056 701792
rect 396992 701732 396996 701788
rect 396996 701732 397052 701788
rect 397052 701732 397056 701788
rect 396992 701728 397056 701732
rect 397072 701788 397136 701792
rect 397072 701732 397076 701788
rect 397076 701732 397132 701788
rect 397132 701732 397136 701788
rect 397072 701728 397136 701732
rect 397152 701788 397216 701792
rect 397152 701732 397156 701788
rect 397156 701732 397212 701788
rect 397212 701732 397216 701788
rect 397152 701728 397216 701732
rect 397232 701788 397296 701792
rect 397232 701732 397236 701788
rect 397236 701732 397292 701788
rect 397292 701732 397296 701788
rect 397232 701728 397296 701732
rect 397312 701788 397376 701792
rect 397312 701732 397316 701788
rect 397316 701732 397372 701788
rect 397372 701732 397376 701788
rect 397312 701728 397376 701732
rect 432832 701788 432896 701792
rect 432832 701732 432836 701788
rect 432836 701732 432892 701788
rect 432892 701732 432896 701788
rect 432832 701728 432896 701732
rect 432912 701788 432976 701792
rect 432912 701732 432916 701788
rect 432916 701732 432972 701788
rect 432972 701732 432976 701788
rect 432912 701728 432976 701732
rect 432992 701788 433056 701792
rect 432992 701732 432996 701788
rect 432996 701732 433052 701788
rect 433052 701732 433056 701788
rect 432992 701728 433056 701732
rect 433072 701788 433136 701792
rect 433072 701732 433076 701788
rect 433076 701732 433132 701788
rect 433132 701732 433136 701788
rect 433072 701728 433136 701732
rect 433152 701788 433216 701792
rect 433152 701732 433156 701788
rect 433156 701732 433212 701788
rect 433212 701732 433216 701788
rect 433152 701728 433216 701732
rect 433232 701788 433296 701792
rect 433232 701732 433236 701788
rect 433236 701732 433292 701788
rect 433292 701732 433296 701788
rect 433232 701728 433296 701732
rect 433312 701788 433376 701792
rect 433312 701732 433316 701788
rect 433316 701732 433372 701788
rect 433372 701732 433376 701788
rect 433312 701728 433376 701732
rect 468832 701788 468896 701792
rect 468832 701732 468836 701788
rect 468836 701732 468892 701788
rect 468892 701732 468896 701788
rect 468832 701728 468896 701732
rect 468912 701788 468976 701792
rect 468912 701732 468916 701788
rect 468916 701732 468972 701788
rect 468972 701732 468976 701788
rect 468912 701728 468976 701732
rect 468992 701788 469056 701792
rect 468992 701732 468996 701788
rect 468996 701732 469052 701788
rect 469052 701732 469056 701788
rect 468992 701728 469056 701732
rect 469072 701788 469136 701792
rect 469072 701732 469076 701788
rect 469076 701732 469132 701788
rect 469132 701732 469136 701788
rect 469072 701728 469136 701732
rect 469152 701788 469216 701792
rect 469152 701732 469156 701788
rect 469156 701732 469212 701788
rect 469212 701732 469216 701788
rect 469152 701728 469216 701732
rect 469232 701788 469296 701792
rect 469232 701732 469236 701788
rect 469236 701732 469292 701788
rect 469292 701732 469296 701788
rect 469232 701728 469296 701732
rect 469312 701788 469376 701792
rect 469312 701732 469316 701788
rect 469316 701732 469372 701788
rect 469372 701732 469376 701788
rect 469312 701728 469376 701732
rect 504832 701788 504896 701792
rect 504832 701732 504836 701788
rect 504836 701732 504892 701788
rect 504892 701732 504896 701788
rect 504832 701728 504896 701732
rect 504912 701788 504976 701792
rect 504912 701732 504916 701788
rect 504916 701732 504972 701788
rect 504972 701732 504976 701788
rect 504912 701728 504976 701732
rect 504992 701788 505056 701792
rect 504992 701732 504996 701788
rect 504996 701732 505052 701788
rect 505052 701732 505056 701788
rect 504992 701728 505056 701732
rect 505072 701788 505136 701792
rect 505072 701732 505076 701788
rect 505076 701732 505132 701788
rect 505132 701732 505136 701788
rect 505072 701728 505136 701732
rect 505152 701788 505216 701792
rect 505152 701732 505156 701788
rect 505156 701732 505212 701788
rect 505212 701732 505216 701788
rect 505152 701728 505216 701732
rect 505232 701788 505296 701792
rect 505232 701732 505236 701788
rect 505236 701732 505292 701788
rect 505292 701732 505296 701788
rect 505232 701728 505296 701732
rect 505312 701788 505376 701792
rect 505312 701732 505316 701788
rect 505316 701732 505372 701788
rect 505372 701732 505376 701788
rect 505312 701728 505376 701732
rect 540832 701788 540896 701792
rect 540832 701732 540836 701788
rect 540836 701732 540892 701788
rect 540892 701732 540896 701788
rect 540832 701728 540896 701732
rect 540912 701788 540976 701792
rect 540912 701732 540916 701788
rect 540916 701732 540972 701788
rect 540972 701732 540976 701788
rect 540912 701728 540976 701732
rect 540992 701788 541056 701792
rect 540992 701732 540996 701788
rect 540996 701732 541052 701788
rect 541052 701732 541056 701788
rect 540992 701728 541056 701732
rect 541072 701788 541136 701792
rect 541072 701732 541076 701788
rect 541076 701732 541132 701788
rect 541132 701732 541136 701788
rect 541072 701728 541136 701732
rect 541152 701788 541216 701792
rect 541152 701732 541156 701788
rect 541156 701732 541212 701788
rect 541212 701732 541216 701788
rect 541152 701728 541216 701732
rect 541232 701788 541296 701792
rect 541232 701732 541236 701788
rect 541236 701732 541292 701788
rect 541292 701732 541296 701788
rect 541232 701728 541296 701732
rect 541312 701788 541376 701792
rect 541312 701732 541316 701788
rect 541316 701732 541372 701788
rect 541372 701732 541376 701788
rect 541312 701728 541376 701732
rect 576832 701788 576896 701792
rect 576832 701732 576836 701788
rect 576836 701732 576892 701788
rect 576892 701732 576896 701788
rect 576832 701728 576896 701732
rect 576912 701788 576976 701792
rect 576912 701732 576916 701788
rect 576916 701732 576972 701788
rect 576972 701732 576976 701788
rect 576912 701728 576976 701732
rect 576992 701788 577056 701792
rect 576992 701732 576996 701788
rect 576996 701732 577052 701788
rect 577052 701732 577056 701788
rect 576992 701728 577056 701732
rect 577072 701788 577136 701792
rect 577072 701732 577076 701788
rect 577076 701732 577132 701788
rect 577132 701732 577136 701788
rect 577072 701728 577136 701732
rect 577152 701788 577216 701792
rect 577152 701732 577156 701788
rect 577156 701732 577212 701788
rect 577212 701732 577216 701788
rect 577152 701728 577216 701732
rect 577232 701788 577296 701792
rect 577232 701732 577236 701788
rect 577236 701732 577292 701788
rect 577292 701732 577296 701788
rect 577232 701728 577296 701732
rect 577312 701788 577376 701792
rect 577312 701732 577316 701788
rect 577316 701732 577372 701788
rect 577372 701732 577376 701788
rect 577312 701728 577376 701732
rect 18832 701244 18896 701248
rect 18832 701188 18836 701244
rect 18836 701188 18892 701244
rect 18892 701188 18896 701244
rect 18832 701184 18896 701188
rect 18912 701244 18976 701248
rect 18912 701188 18916 701244
rect 18916 701188 18972 701244
rect 18972 701188 18976 701244
rect 18912 701184 18976 701188
rect 18992 701244 19056 701248
rect 18992 701188 18996 701244
rect 18996 701188 19052 701244
rect 19052 701188 19056 701244
rect 18992 701184 19056 701188
rect 19072 701244 19136 701248
rect 19072 701188 19076 701244
rect 19076 701188 19132 701244
rect 19132 701188 19136 701244
rect 19072 701184 19136 701188
rect 19152 701244 19216 701248
rect 19152 701188 19156 701244
rect 19156 701188 19212 701244
rect 19212 701188 19216 701244
rect 19152 701184 19216 701188
rect 19232 701244 19296 701248
rect 19232 701188 19236 701244
rect 19236 701188 19292 701244
rect 19292 701188 19296 701244
rect 19232 701184 19296 701188
rect 19312 701244 19376 701248
rect 19312 701188 19316 701244
rect 19316 701188 19372 701244
rect 19372 701188 19376 701244
rect 19312 701184 19376 701188
rect 54832 701244 54896 701248
rect 54832 701188 54836 701244
rect 54836 701188 54892 701244
rect 54892 701188 54896 701244
rect 54832 701184 54896 701188
rect 54912 701244 54976 701248
rect 54912 701188 54916 701244
rect 54916 701188 54972 701244
rect 54972 701188 54976 701244
rect 54912 701184 54976 701188
rect 54992 701244 55056 701248
rect 54992 701188 54996 701244
rect 54996 701188 55052 701244
rect 55052 701188 55056 701244
rect 54992 701184 55056 701188
rect 55072 701244 55136 701248
rect 55072 701188 55076 701244
rect 55076 701188 55132 701244
rect 55132 701188 55136 701244
rect 55072 701184 55136 701188
rect 55152 701244 55216 701248
rect 55152 701188 55156 701244
rect 55156 701188 55212 701244
rect 55212 701188 55216 701244
rect 55152 701184 55216 701188
rect 55232 701244 55296 701248
rect 55232 701188 55236 701244
rect 55236 701188 55292 701244
rect 55292 701188 55296 701244
rect 55232 701184 55296 701188
rect 55312 701244 55376 701248
rect 55312 701188 55316 701244
rect 55316 701188 55372 701244
rect 55372 701188 55376 701244
rect 55312 701184 55376 701188
rect 90832 701244 90896 701248
rect 90832 701188 90836 701244
rect 90836 701188 90892 701244
rect 90892 701188 90896 701244
rect 90832 701184 90896 701188
rect 90912 701244 90976 701248
rect 90912 701188 90916 701244
rect 90916 701188 90972 701244
rect 90972 701188 90976 701244
rect 90912 701184 90976 701188
rect 90992 701244 91056 701248
rect 90992 701188 90996 701244
rect 90996 701188 91052 701244
rect 91052 701188 91056 701244
rect 90992 701184 91056 701188
rect 91072 701244 91136 701248
rect 91072 701188 91076 701244
rect 91076 701188 91132 701244
rect 91132 701188 91136 701244
rect 91072 701184 91136 701188
rect 91152 701244 91216 701248
rect 91152 701188 91156 701244
rect 91156 701188 91212 701244
rect 91212 701188 91216 701244
rect 91152 701184 91216 701188
rect 91232 701244 91296 701248
rect 91232 701188 91236 701244
rect 91236 701188 91292 701244
rect 91292 701188 91296 701244
rect 91232 701184 91296 701188
rect 91312 701244 91376 701248
rect 91312 701188 91316 701244
rect 91316 701188 91372 701244
rect 91372 701188 91376 701244
rect 91312 701184 91376 701188
rect 126832 701244 126896 701248
rect 126832 701188 126836 701244
rect 126836 701188 126892 701244
rect 126892 701188 126896 701244
rect 126832 701184 126896 701188
rect 126912 701244 126976 701248
rect 126912 701188 126916 701244
rect 126916 701188 126972 701244
rect 126972 701188 126976 701244
rect 126912 701184 126976 701188
rect 126992 701244 127056 701248
rect 126992 701188 126996 701244
rect 126996 701188 127052 701244
rect 127052 701188 127056 701244
rect 126992 701184 127056 701188
rect 127072 701244 127136 701248
rect 127072 701188 127076 701244
rect 127076 701188 127132 701244
rect 127132 701188 127136 701244
rect 127072 701184 127136 701188
rect 127152 701244 127216 701248
rect 127152 701188 127156 701244
rect 127156 701188 127212 701244
rect 127212 701188 127216 701244
rect 127152 701184 127216 701188
rect 127232 701244 127296 701248
rect 127232 701188 127236 701244
rect 127236 701188 127292 701244
rect 127292 701188 127296 701244
rect 127232 701184 127296 701188
rect 127312 701244 127376 701248
rect 127312 701188 127316 701244
rect 127316 701188 127372 701244
rect 127372 701188 127376 701244
rect 127312 701184 127376 701188
rect 162832 701244 162896 701248
rect 162832 701188 162836 701244
rect 162836 701188 162892 701244
rect 162892 701188 162896 701244
rect 162832 701184 162896 701188
rect 162912 701244 162976 701248
rect 162912 701188 162916 701244
rect 162916 701188 162972 701244
rect 162972 701188 162976 701244
rect 162912 701184 162976 701188
rect 162992 701244 163056 701248
rect 162992 701188 162996 701244
rect 162996 701188 163052 701244
rect 163052 701188 163056 701244
rect 162992 701184 163056 701188
rect 163072 701244 163136 701248
rect 163072 701188 163076 701244
rect 163076 701188 163132 701244
rect 163132 701188 163136 701244
rect 163072 701184 163136 701188
rect 163152 701244 163216 701248
rect 163152 701188 163156 701244
rect 163156 701188 163212 701244
rect 163212 701188 163216 701244
rect 163152 701184 163216 701188
rect 163232 701244 163296 701248
rect 163232 701188 163236 701244
rect 163236 701188 163292 701244
rect 163292 701188 163296 701244
rect 163232 701184 163296 701188
rect 163312 701244 163376 701248
rect 163312 701188 163316 701244
rect 163316 701188 163372 701244
rect 163372 701188 163376 701244
rect 163312 701184 163376 701188
rect 198832 701244 198896 701248
rect 198832 701188 198836 701244
rect 198836 701188 198892 701244
rect 198892 701188 198896 701244
rect 198832 701184 198896 701188
rect 198912 701244 198976 701248
rect 198912 701188 198916 701244
rect 198916 701188 198972 701244
rect 198972 701188 198976 701244
rect 198912 701184 198976 701188
rect 198992 701244 199056 701248
rect 198992 701188 198996 701244
rect 198996 701188 199052 701244
rect 199052 701188 199056 701244
rect 198992 701184 199056 701188
rect 199072 701244 199136 701248
rect 199072 701188 199076 701244
rect 199076 701188 199132 701244
rect 199132 701188 199136 701244
rect 199072 701184 199136 701188
rect 199152 701244 199216 701248
rect 199152 701188 199156 701244
rect 199156 701188 199212 701244
rect 199212 701188 199216 701244
rect 199152 701184 199216 701188
rect 199232 701244 199296 701248
rect 199232 701188 199236 701244
rect 199236 701188 199292 701244
rect 199292 701188 199296 701244
rect 199232 701184 199296 701188
rect 199312 701244 199376 701248
rect 199312 701188 199316 701244
rect 199316 701188 199372 701244
rect 199372 701188 199376 701244
rect 199312 701184 199376 701188
rect 234832 701244 234896 701248
rect 234832 701188 234836 701244
rect 234836 701188 234892 701244
rect 234892 701188 234896 701244
rect 234832 701184 234896 701188
rect 234912 701244 234976 701248
rect 234912 701188 234916 701244
rect 234916 701188 234972 701244
rect 234972 701188 234976 701244
rect 234912 701184 234976 701188
rect 234992 701244 235056 701248
rect 234992 701188 234996 701244
rect 234996 701188 235052 701244
rect 235052 701188 235056 701244
rect 234992 701184 235056 701188
rect 235072 701244 235136 701248
rect 235072 701188 235076 701244
rect 235076 701188 235132 701244
rect 235132 701188 235136 701244
rect 235072 701184 235136 701188
rect 235152 701244 235216 701248
rect 235152 701188 235156 701244
rect 235156 701188 235212 701244
rect 235212 701188 235216 701244
rect 235152 701184 235216 701188
rect 235232 701244 235296 701248
rect 235232 701188 235236 701244
rect 235236 701188 235292 701244
rect 235292 701188 235296 701244
rect 235232 701184 235296 701188
rect 235312 701244 235376 701248
rect 235312 701188 235316 701244
rect 235316 701188 235372 701244
rect 235372 701188 235376 701244
rect 235312 701184 235376 701188
rect 270832 701244 270896 701248
rect 270832 701188 270836 701244
rect 270836 701188 270892 701244
rect 270892 701188 270896 701244
rect 270832 701184 270896 701188
rect 270912 701244 270976 701248
rect 270912 701188 270916 701244
rect 270916 701188 270972 701244
rect 270972 701188 270976 701244
rect 270912 701184 270976 701188
rect 270992 701244 271056 701248
rect 270992 701188 270996 701244
rect 270996 701188 271052 701244
rect 271052 701188 271056 701244
rect 270992 701184 271056 701188
rect 271072 701244 271136 701248
rect 271072 701188 271076 701244
rect 271076 701188 271132 701244
rect 271132 701188 271136 701244
rect 271072 701184 271136 701188
rect 271152 701244 271216 701248
rect 271152 701188 271156 701244
rect 271156 701188 271212 701244
rect 271212 701188 271216 701244
rect 271152 701184 271216 701188
rect 271232 701244 271296 701248
rect 271232 701188 271236 701244
rect 271236 701188 271292 701244
rect 271292 701188 271296 701244
rect 271232 701184 271296 701188
rect 271312 701244 271376 701248
rect 271312 701188 271316 701244
rect 271316 701188 271372 701244
rect 271372 701188 271376 701244
rect 271312 701184 271376 701188
rect 306832 701244 306896 701248
rect 306832 701188 306836 701244
rect 306836 701188 306892 701244
rect 306892 701188 306896 701244
rect 306832 701184 306896 701188
rect 306912 701244 306976 701248
rect 306912 701188 306916 701244
rect 306916 701188 306972 701244
rect 306972 701188 306976 701244
rect 306912 701184 306976 701188
rect 306992 701244 307056 701248
rect 306992 701188 306996 701244
rect 306996 701188 307052 701244
rect 307052 701188 307056 701244
rect 306992 701184 307056 701188
rect 307072 701244 307136 701248
rect 307072 701188 307076 701244
rect 307076 701188 307132 701244
rect 307132 701188 307136 701244
rect 307072 701184 307136 701188
rect 307152 701244 307216 701248
rect 307152 701188 307156 701244
rect 307156 701188 307212 701244
rect 307212 701188 307216 701244
rect 307152 701184 307216 701188
rect 307232 701244 307296 701248
rect 307232 701188 307236 701244
rect 307236 701188 307292 701244
rect 307292 701188 307296 701244
rect 307232 701184 307296 701188
rect 307312 701244 307376 701248
rect 307312 701188 307316 701244
rect 307316 701188 307372 701244
rect 307372 701188 307376 701244
rect 307312 701184 307376 701188
rect 342832 701244 342896 701248
rect 342832 701188 342836 701244
rect 342836 701188 342892 701244
rect 342892 701188 342896 701244
rect 342832 701184 342896 701188
rect 342912 701244 342976 701248
rect 342912 701188 342916 701244
rect 342916 701188 342972 701244
rect 342972 701188 342976 701244
rect 342912 701184 342976 701188
rect 342992 701244 343056 701248
rect 342992 701188 342996 701244
rect 342996 701188 343052 701244
rect 343052 701188 343056 701244
rect 342992 701184 343056 701188
rect 343072 701244 343136 701248
rect 343072 701188 343076 701244
rect 343076 701188 343132 701244
rect 343132 701188 343136 701244
rect 343072 701184 343136 701188
rect 343152 701244 343216 701248
rect 343152 701188 343156 701244
rect 343156 701188 343212 701244
rect 343212 701188 343216 701244
rect 343152 701184 343216 701188
rect 343232 701244 343296 701248
rect 343232 701188 343236 701244
rect 343236 701188 343292 701244
rect 343292 701188 343296 701244
rect 343232 701184 343296 701188
rect 343312 701244 343376 701248
rect 343312 701188 343316 701244
rect 343316 701188 343372 701244
rect 343372 701188 343376 701244
rect 343312 701184 343376 701188
rect 378832 701244 378896 701248
rect 378832 701188 378836 701244
rect 378836 701188 378892 701244
rect 378892 701188 378896 701244
rect 378832 701184 378896 701188
rect 378912 701244 378976 701248
rect 378912 701188 378916 701244
rect 378916 701188 378972 701244
rect 378972 701188 378976 701244
rect 378912 701184 378976 701188
rect 378992 701244 379056 701248
rect 378992 701188 378996 701244
rect 378996 701188 379052 701244
rect 379052 701188 379056 701244
rect 378992 701184 379056 701188
rect 379072 701244 379136 701248
rect 379072 701188 379076 701244
rect 379076 701188 379132 701244
rect 379132 701188 379136 701244
rect 379072 701184 379136 701188
rect 379152 701244 379216 701248
rect 379152 701188 379156 701244
rect 379156 701188 379212 701244
rect 379212 701188 379216 701244
rect 379152 701184 379216 701188
rect 379232 701244 379296 701248
rect 379232 701188 379236 701244
rect 379236 701188 379292 701244
rect 379292 701188 379296 701244
rect 379232 701184 379296 701188
rect 379312 701244 379376 701248
rect 379312 701188 379316 701244
rect 379316 701188 379372 701244
rect 379372 701188 379376 701244
rect 379312 701184 379376 701188
rect 414832 701244 414896 701248
rect 414832 701188 414836 701244
rect 414836 701188 414892 701244
rect 414892 701188 414896 701244
rect 414832 701184 414896 701188
rect 414912 701244 414976 701248
rect 414912 701188 414916 701244
rect 414916 701188 414972 701244
rect 414972 701188 414976 701244
rect 414912 701184 414976 701188
rect 414992 701244 415056 701248
rect 414992 701188 414996 701244
rect 414996 701188 415052 701244
rect 415052 701188 415056 701244
rect 414992 701184 415056 701188
rect 415072 701244 415136 701248
rect 415072 701188 415076 701244
rect 415076 701188 415132 701244
rect 415132 701188 415136 701244
rect 415072 701184 415136 701188
rect 415152 701244 415216 701248
rect 415152 701188 415156 701244
rect 415156 701188 415212 701244
rect 415212 701188 415216 701244
rect 415152 701184 415216 701188
rect 415232 701244 415296 701248
rect 415232 701188 415236 701244
rect 415236 701188 415292 701244
rect 415292 701188 415296 701244
rect 415232 701184 415296 701188
rect 415312 701244 415376 701248
rect 415312 701188 415316 701244
rect 415316 701188 415372 701244
rect 415372 701188 415376 701244
rect 415312 701184 415376 701188
rect 450832 701244 450896 701248
rect 450832 701188 450836 701244
rect 450836 701188 450892 701244
rect 450892 701188 450896 701244
rect 450832 701184 450896 701188
rect 450912 701244 450976 701248
rect 450912 701188 450916 701244
rect 450916 701188 450972 701244
rect 450972 701188 450976 701244
rect 450912 701184 450976 701188
rect 450992 701244 451056 701248
rect 450992 701188 450996 701244
rect 450996 701188 451052 701244
rect 451052 701188 451056 701244
rect 450992 701184 451056 701188
rect 451072 701244 451136 701248
rect 451072 701188 451076 701244
rect 451076 701188 451132 701244
rect 451132 701188 451136 701244
rect 451072 701184 451136 701188
rect 451152 701244 451216 701248
rect 451152 701188 451156 701244
rect 451156 701188 451212 701244
rect 451212 701188 451216 701244
rect 451152 701184 451216 701188
rect 451232 701244 451296 701248
rect 451232 701188 451236 701244
rect 451236 701188 451292 701244
rect 451292 701188 451296 701244
rect 451232 701184 451296 701188
rect 451312 701244 451376 701248
rect 451312 701188 451316 701244
rect 451316 701188 451372 701244
rect 451372 701188 451376 701244
rect 451312 701184 451376 701188
rect 486832 701244 486896 701248
rect 486832 701188 486836 701244
rect 486836 701188 486892 701244
rect 486892 701188 486896 701244
rect 486832 701184 486896 701188
rect 486912 701244 486976 701248
rect 486912 701188 486916 701244
rect 486916 701188 486972 701244
rect 486972 701188 486976 701244
rect 486912 701184 486976 701188
rect 486992 701244 487056 701248
rect 486992 701188 486996 701244
rect 486996 701188 487052 701244
rect 487052 701188 487056 701244
rect 486992 701184 487056 701188
rect 487072 701244 487136 701248
rect 487072 701188 487076 701244
rect 487076 701188 487132 701244
rect 487132 701188 487136 701244
rect 487072 701184 487136 701188
rect 487152 701244 487216 701248
rect 487152 701188 487156 701244
rect 487156 701188 487212 701244
rect 487212 701188 487216 701244
rect 487152 701184 487216 701188
rect 487232 701244 487296 701248
rect 487232 701188 487236 701244
rect 487236 701188 487292 701244
rect 487292 701188 487296 701244
rect 487232 701184 487296 701188
rect 487312 701244 487376 701248
rect 487312 701188 487316 701244
rect 487316 701188 487372 701244
rect 487372 701188 487376 701244
rect 487312 701184 487376 701188
rect 522832 701244 522896 701248
rect 522832 701188 522836 701244
rect 522836 701188 522892 701244
rect 522892 701188 522896 701244
rect 522832 701184 522896 701188
rect 522912 701244 522976 701248
rect 522912 701188 522916 701244
rect 522916 701188 522972 701244
rect 522972 701188 522976 701244
rect 522912 701184 522976 701188
rect 522992 701244 523056 701248
rect 522992 701188 522996 701244
rect 522996 701188 523052 701244
rect 523052 701188 523056 701244
rect 522992 701184 523056 701188
rect 523072 701244 523136 701248
rect 523072 701188 523076 701244
rect 523076 701188 523132 701244
rect 523132 701188 523136 701244
rect 523072 701184 523136 701188
rect 523152 701244 523216 701248
rect 523152 701188 523156 701244
rect 523156 701188 523212 701244
rect 523212 701188 523216 701244
rect 523152 701184 523216 701188
rect 523232 701244 523296 701248
rect 523232 701188 523236 701244
rect 523236 701188 523292 701244
rect 523292 701188 523296 701244
rect 523232 701184 523296 701188
rect 523312 701244 523376 701248
rect 523312 701188 523316 701244
rect 523316 701188 523372 701244
rect 523372 701188 523376 701244
rect 523312 701184 523376 701188
rect 558832 701244 558896 701248
rect 558832 701188 558836 701244
rect 558836 701188 558892 701244
rect 558892 701188 558896 701244
rect 558832 701184 558896 701188
rect 558912 701244 558976 701248
rect 558912 701188 558916 701244
rect 558916 701188 558972 701244
rect 558972 701188 558976 701244
rect 558912 701184 558976 701188
rect 558992 701244 559056 701248
rect 558992 701188 558996 701244
rect 558996 701188 559052 701244
rect 559052 701188 559056 701244
rect 558992 701184 559056 701188
rect 559072 701244 559136 701248
rect 559072 701188 559076 701244
rect 559076 701188 559132 701244
rect 559132 701188 559136 701244
rect 559072 701184 559136 701188
rect 559152 701244 559216 701248
rect 559152 701188 559156 701244
rect 559156 701188 559212 701244
rect 559212 701188 559216 701244
rect 559152 701184 559216 701188
rect 559232 701244 559296 701248
rect 559232 701188 559236 701244
rect 559236 701188 559292 701244
rect 559292 701188 559296 701244
rect 559232 701184 559296 701188
rect 559312 701244 559376 701248
rect 559312 701188 559316 701244
rect 559316 701188 559372 701244
rect 559372 701188 559376 701244
rect 559312 701184 559376 701188
rect 36832 700700 36896 700704
rect 36832 700644 36836 700700
rect 36836 700644 36892 700700
rect 36892 700644 36896 700700
rect 36832 700640 36896 700644
rect 36912 700700 36976 700704
rect 36912 700644 36916 700700
rect 36916 700644 36972 700700
rect 36972 700644 36976 700700
rect 36912 700640 36976 700644
rect 36992 700700 37056 700704
rect 36992 700644 36996 700700
rect 36996 700644 37052 700700
rect 37052 700644 37056 700700
rect 36992 700640 37056 700644
rect 37072 700700 37136 700704
rect 37072 700644 37076 700700
rect 37076 700644 37132 700700
rect 37132 700644 37136 700700
rect 37072 700640 37136 700644
rect 37152 700700 37216 700704
rect 37152 700644 37156 700700
rect 37156 700644 37212 700700
rect 37212 700644 37216 700700
rect 37152 700640 37216 700644
rect 37232 700700 37296 700704
rect 37232 700644 37236 700700
rect 37236 700644 37292 700700
rect 37292 700644 37296 700700
rect 37232 700640 37296 700644
rect 37312 700700 37376 700704
rect 37312 700644 37316 700700
rect 37316 700644 37372 700700
rect 37372 700644 37376 700700
rect 37312 700640 37376 700644
rect 72832 700700 72896 700704
rect 72832 700644 72836 700700
rect 72836 700644 72892 700700
rect 72892 700644 72896 700700
rect 72832 700640 72896 700644
rect 72912 700700 72976 700704
rect 72912 700644 72916 700700
rect 72916 700644 72972 700700
rect 72972 700644 72976 700700
rect 72912 700640 72976 700644
rect 72992 700700 73056 700704
rect 72992 700644 72996 700700
rect 72996 700644 73052 700700
rect 73052 700644 73056 700700
rect 72992 700640 73056 700644
rect 73072 700700 73136 700704
rect 73072 700644 73076 700700
rect 73076 700644 73132 700700
rect 73132 700644 73136 700700
rect 73072 700640 73136 700644
rect 73152 700700 73216 700704
rect 73152 700644 73156 700700
rect 73156 700644 73212 700700
rect 73212 700644 73216 700700
rect 73152 700640 73216 700644
rect 73232 700700 73296 700704
rect 73232 700644 73236 700700
rect 73236 700644 73292 700700
rect 73292 700644 73296 700700
rect 73232 700640 73296 700644
rect 73312 700700 73376 700704
rect 73312 700644 73316 700700
rect 73316 700644 73372 700700
rect 73372 700644 73376 700700
rect 73312 700640 73376 700644
rect 108832 700700 108896 700704
rect 108832 700644 108836 700700
rect 108836 700644 108892 700700
rect 108892 700644 108896 700700
rect 108832 700640 108896 700644
rect 108912 700700 108976 700704
rect 108912 700644 108916 700700
rect 108916 700644 108972 700700
rect 108972 700644 108976 700700
rect 108912 700640 108976 700644
rect 108992 700700 109056 700704
rect 108992 700644 108996 700700
rect 108996 700644 109052 700700
rect 109052 700644 109056 700700
rect 108992 700640 109056 700644
rect 109072 700700 109136 700704
rect 109072 700644 109076 700700
rect 109076 700644 109132 700700
rect 109132 700644 109136 700700
rect 109072 700640 109136 700644
rect 109152 700700 109216 700704
rect 109152 700644 109156 700700
rect 109156 700644 109212 700700
rect 109212 700644 109216 700700
rect 109152 700640 109216 700644
rect 109232 700700 109296 700704
rect 109232 700644 109236 700700
rect 109236 700644 109292 700700
rect 109292 700644 109296 700700
rect 109232 700640 109296 700644
rect 109312 700700 109376 700704
rect 109312 700644 109316 700700
rect 109316 700644 109372 700700
rect 109372 700644 109376 700700
rect 109312 700640 109376 700644
rect 144832 700700 144896 700704
rect 144832 700644 144836 700700
rect 144836 700644 144892 700700
rect 144892 700644 144896 700700
rect 144832 700640 144896 700644
rect 144912 700700 144976 700704
rect 144912 700644 144916 700700
rect 144916 700644 144972 700700
rect 144972 700644 144976 700700
rect 144912 700640 144976 700644
rect 144992 700700 145056 700704
rect 144992 700644 144996 700700
rect 144996 700644 145052 700700
rect 145052 700644 145056 700700
rect 144992 700640 145056 700644
rect 145072 700700 145136 700704
rect 145072 700644 145076 700700
rect 145076 700644 145132 700700
rect 145132 700644 145136 700700
rect 145072 700640 145136 700644
rect 145152 700700 145216 700704
rect 145152 700644 145156 700700
rect 145156 700644 145212 700700
rect 145212 700644 145216 700700
rect 145152 700640 145216 700644
rect 145232 700700 145296 700704
rect 145232 700644 145236 700700
rect 145236 700644 145292 700700
rect 145292 700644 145296 700700
rect 145232 700640 145296 700644
rect 145312 700700 145376 700704
rect 145312 700644 145316 700700
rect 145316 700644 145372 700700
rect 145372 700644 145376 700700
rect 145312 700640 145376 700644
rect 180832 700700 180896 700704
rect 180832 700644 180836 700700
rect 180836 700644 180892 700700
rect 180892 700644 180896 700700
rect 180832 700640 180896 700644
rect 180912 700700 180976 700704
rect 180912 700644 180916 700700
rect 180916 700644 180972 700700
rect 180972 700644 180976 700700
rect 180912 700640 180976 700644
rect 180992 700700 181056 700704
rect 180992 700644 180996 700700
rect 180996 700644 181052 700700
rect 181052 700644 181056 700700
rect 180992 700640 181056 700644
rect 181072 700700 181136 700704
rect 181072 700644 181076 700700
rect 181076 700644 181132 700700
rect 181132 700644 181136 700700
rect 181072 700640 181136 700644
rect 181152 700700 181216 700704
rect 181152 700644 181156 700700
rect 181156 700644 181212 700700
rect 181212 700644 181216 700700
rect 181152 700640 181216 700644
rect 181232 700700 181296 700704
rect 181232 700644 181236 700700
rect 181236 700644 181292 700700
rect 181292 700644 181296 700700
rect 181232 700640 181296 700644
rect 181312 700700 181376 700704
rect 181312 700644 181316 700700
rect 181316 700644 181372 700700
rect 181372 700644 181376 700700
rect 181312 700640 181376 700644
rect 216832 700700 216896 700704
rect 216832 700644 216836 700700
rect 216836 700644 216892 700700
rect 216892 700644 216896 700700
rect 216832 700640 216896 700644
rect 216912 700700 216976 700704
rect 216912 700644 216916 700700
rect 216916 700644 216972 700700
rect 216972 700644 216976 700700
rect 216912 700640 216976 700644
rect 216992 700700 217056 700704
rect 216992 700644 216996 700700
rect 216996 700644 217052 700700
rect 217052 700644 217056 700700
rect 216992 700640 217056 700644
rect 217072 700700 217136 700704
rect 217072 700644 217076 700700
rect 217076 700644 217132 700700
rect 217132 700644 217136 700700
rect 217072 700640 217136 700644
rect 217152 700700 217216 700704
rect 217152 700644 217156 700700
rect 217156 700644 217212 700700
rect 217212 700644 217216 700700
rect 217152 700640 217216 700644
rect 217232 700700 217296 700704
rect 217232 700644 217236 700700
rect 217236 700644 217292 700700
rect 217292 700644 217296 700700
rect 217232 700640 217296 700644
rect 217312 700700 217376 700704
rect 217312 700644 217316 700700
rect 217316 700644 217372 700700
rect 217372 700644 217376 700700
rect 217312 700640 217376 700644
rect 252832 700700 252896 700704
rect 252832 700644 252836 700700
rect 252836 700644 252892 700700
rect 252892 700644 252896 700700
rect 252832 700640 252896 700644
rect 252912 700700 252976 700704
rect 252912 700644 252916 700700
rect 252916 700644 252972 700700
rect 252972 700644 252976 700700
rect 252912 700640 252976 700644
rect 252992 700700 253056 700704
rect 252992 700644 252996 700700
rect 252996 700644 253052 700700
rect 253052 700644 253056 700700
rect 252992 700640 253056 700644
rect 253072 700700 253136 700704
rect 253072 700644 253076 700700
rect 253076 700644 253132 700700
rect 253132 700644 253136 700700
rect 253072 700640 253136 700644
rect 253152 700700 253216 700704
rect 253152 700644 253156 700700
rect 253156 700644 253212 700700
rect 253212 700644 253216 700700
rect 253152 700640 253216 700644
rect 253232 700700 253296 700704
rect 253232 700644 253236 700700
rect 253236 700644 253292 700700
rect 253292 700644 253296 700700
rect 253232 700640 253296 700644
rect 253312 700700 253376 700704
rect 253312 700644 253316 700700
rect 253316 700644 253372 700700
rect 253372 700644 253376 700700
rect 253312 700640 253376 700644
rect 288832 700700 288896 700704
rect 288832 700644 288836 700700
rect 288836 700644 288892 700700
rect 288892 700644 288896 700700
rect 288832 700640 288896 700644
rect 288912 700700 288976 700704
rect 288912 700644 288916 700700
rect 288916 700644 288972 700700
rect 288972 700644 288976 700700
rect 288912 700640 288976 700644
rect 288992 700700 289056 700704
rect 288992 700644 288996 700700
rect 288996 700644 289052 700700
rect 289052 700644 289056 700700
rect 288992 700640 289056 700644
rect 289072 700700 289136 700704
rect 289072 700644 289076 700700
rect 289076 700644 289132 700700
rect 289132 700644 289136 700700
rect 289072 700640 289136 700644
rect 289152 700700 289216 700704
rect 289152 700644 289156 700700
rect 289156 700644 289212 700700
rect 289212 700644 289216 700700
rect 289152 700640 289216 700644
rect 289232 700700 289296 700704
rect 289232 700644 289236 700700
rect 289236 700644 289292 700700
rect 289292 700644 289296 700700
rect 289232 700640 289296 700644
rect 289312 700700 289376 700704
rect 289312 700644 289316 700700
rect 289316 700644 289372 700700
rect 289372 700644 289376 700700
rect 289312 700640 289376 700644
rect 324832 700700 324896 700704
rect 324832 700644 324836 700700
rect 324836 700644 324892 700700
rect 324892 700644 324896 700700
rect 324832 700640 324896 700644
rect 324912 700700 324976 700704
rect 324912 700644 324916 700700
rect 324916 700644 324972 700700
rect 324972 700644 324976 700700
rect 324912 700640 324976 700644
rect 324992 700700 325056 700704
rect 324992 700644 324996 700700
rect 324996 700644 325052 700700
rect 325052 700644 325056 700700
rect 324992 700640 325056 700644
rect 325072 700700 325136 700704
rect 325072 700644 325076 700700
rect 325076 700644 325132 700700
rect 325132 700644 325136 700700
rect 325072 700640 325136 700644
rect 325152 700700 325216 700704
rect 325152 700644 325156 700700
rect 325156 700644 325212 700700
rect 325212 700644 325216 700700
rect 325152 700640 325216 700644
rect 325232 700700 325296 700704
rect 325232 700644 325236 700700
rect 325236 700644 325292 700700
rect 325292 700644 325296 700700
rect 325232 700640 325296 700644
rect 325312 700700 325376 700704
rect 325312 700644 325316 700700
rect 325316 700644 325372 700700
rect 325372 700644 325376 700700
rect 325312 700640 325376 700644
rect 360832 700700 360896 700704
rect 360832 700644 360836 700700
rect 360836 700644 360892 700700
rect 360892 700644 360896 700700
rect 360832 700640 360896 700644
rect 360912 700700 360976 700704
rect 360912 700644 360916 700700
rect 360916 700644 360972 700700
rect 360972 700644 360976 700700
rect 360912 700640 360976 700644
rect 360992 700700 361056 700704
rect 360992 700644 360996 700700
rect 360996 700644 361052 700700
rect 361052 700644 361056 700700
rect 360992 700640 361056 700644
rect 361072 700700 361136 700704
rect 361072 700644 361076 700700
rect 361076 700644 361132 700700
rect 361132 700644 361136 700700
rect 361072 700640 361136 700644
rect 361152 700700 361216 700704
rect 361152 700644 361156 700700
rect 361156 700644 361212 700700
rect 361212 700644 361216 700700
rect 361152 700640 361216 700644
rect 361232 700700 361296 700704
rect 361232 700644 361236 700700
rect 361236 700644 361292 700700
rect 361292 700644 361296 700700
rect 361232 700640 361296 700644
rect 361312 700700 361376 700704
rect 361312 700644 361316 700700
rect 361316 700644 361372 700700
rect 361372 700644 361376 700700
rect 361312 700640 361376 700644
rect 396832 700700 396896 700704
rect 396832 700644 396836 700700
rect 396836 700644 396892 700700
rect 396892 700644 396896 700700
rect 396832 700640 396896 700644
rect 396912 700700 396976 700704
rect 396912 700644 396916 700700
rect 396916 700644 396972 700700
rect 396972 700644 396976 700700
rect 396912 700640 396976 700644
rect 396992 700700 397056 700704
rect 396992 700644 396996 700700
rect 396996 700644 397052 700700
rect 397052 700644 397056 700700
rect 396992 700640 397056 700644
rect 397072 700700 397136 700704
rect 397072 700644 397076 700700
rect 397076 700644 397132 700700
rect 397132 700644 397136 700700
rect 397072 700640 397136 700644
rect 397152 700700 397216 700704
rect 397152 700644 397156 700700
rect 397156 700644 397212 700700
rect 397212 700644 397216 700700
rect 397152 700640 397216 700644
rect 397232 700700 397296 700704
rect 397232 700644 397236 700700
rect 397236 700644 397292 700700
rect 397292 700644 397296 700700
rect 397232 700640 397296 700644
rect 397312 700700 397376 700704
rect 397312 700644 397316 700700
rect 397316 700644 397372 700700
rect 397372 700644 397376 700700
rect 397312 700640 397376 700644
rect 432832 700700 432896 700704
rect 432832 700644 432836 700700
rect 432836 700644 432892 700700
rect 432892 700644 432896 700700
rect 432832 700640 432896 700644
rect 432912 700700 432976 700704
rect 432912 700644 432916 700700
rect 432916 700644 432972 700700
rect 432972 700644 432976 700700
rect 432912 700640 432976 700644
rect 432992 700700 433056 700704
rect 432992 700644 432996 700700
rect 432996 700644 433052 700700
rect 433052 700644 433056 700700
rect 432992 700640 433056 700644
rect 433072 700700 433136 700704
rect 433072 700644 433076 700700
rect 433076 700644 433132 700700
rect 433132 700644 433136 700700
rect 433072 700640 433136 700644
rect 433152 700700 433216 700704
rect 433152 700644 433156 700700
rect 433156 700644 433212 700700
rect 433212 700644 433216 700700
rect 433152 700640 433216 700644
rect 433232 700700 433296 700704
rect 433232 700644 433236 700700
rect 433236 700644 433292 700700
rect 433292 700644 433296 700700
rect 433232 700640 433296 700644
rect 433312 700700 433376 700704
rect 433312 700644 433316 700700
rect 433316 700644 433372 700700
rect 433372 700644 433376 700700
rect 433312 700640 433376 700644
rect 468832 700700 468896 700704
rect 468832 700644 468836 700700
rect 468836 700644 468892 700700
rect 468892 700644 468896 700700
rect 468832 700640 468896 700644
rect 468912 700700 468976 700704
rect 468912 700644 468916 700700
rect 468916 700644 468972 700700
rect 468972 700644 468976 700700
rect 468912 700640 468976 700644
rect 468992 700700 469056 700704
rect 468992 700644 468996 700700
rect 468996 700644 469052 700700
rect 469052 700644 469056 700700
rect 468992 700640 469056 700644
rect 469072 700700 469136 700704
rect 469072 700644 469076 700700
rect 469076 700644 469132 700700
rect 469132 700644 469136 700700
rect 469072 700640 469136 700644
rect 469152 700700 469216 700704
rect 469152 700644 469156 700700
rect 469156 700644 469212 700700
rect 469212 700644 469216 700700
rect 469152 700640 469216 700644
rect 469232 700700 469296 700704
rect 469232 700644 469236 700700
rect 469236 700644 469292 700700
rect 469292 700644 469296 700700
rect 469232 700640 469296 700644
rect 469312 700700 469376 700704
rect 469312 700644 469316 700700
rect 469316 700644 469372 700700
rect 469372 700644 469376 700700
rect 469312 700640 469376 700644
rect 504832 700700 504896 700704
rect 504832 700644 504836 700700
rect 504836 700644 504892 700700
rect 504892 700644 504896 700700
rect 504832 700640 504896 700644
rect 504912 700700 504976 700704
rect 504912 700644 504916 700700
rect 504916 700644 504972 700700
rect 504972 700644 504976 700700
rect 504912 700640 504976 700644
rect 504992 700700 505056 700704
rect 504992 700644 504996 700700
rect 504996 700644 505052 700700
rect 505052 700644 505056 700700
rect 504992 700640 505056 700644
rect 505072 700700 505136 700704
rect 505072 700644 505076 700700
rect 505076 700644 505132 700700
rect 505132 700644 505136 700700
rect 505072 700640 505136 700644
rect 505152 700700 505216 700704
rect 505152 700644 505156 700700
rect 505156 700644 505212 700700
rect 505212 700644 505216 700700
rect 505152 700640 505216 700644
rect 505232 700700 505296 700704
rect 505232 700644 505236 700700
rect 505236 700644 505292 700700
rect 505292 700644 505296 700700
rect 505232 700640 505296 700644
rect 505312 700700 505376 700704
rect 505312 700644 505316 700700
rect 505316 700644 505372 700700
rect 505372 700644 505376 700700
rect 505312 700640 505376 700644
rect 540832 700700 540896 700704
rect 540832 700644 540836 700700
rect 540836 700644 540892 700700
rect 540892 700644 540896 700700
rect 540832 700640 540896 700644
rect 540912 700700 540976 700704
rect 540912 700644 540916 700700
rect 540916 700644 540972 700700
rect 540972 700644 540976 700700
rect 540912 700640 540976 700644
rect 540992 700700 541056 700704
rect 540992 700644 540996 700700
rect 540996 700644 541052 700700
rect 541052 700644 541056 700700
rect 540992 700640 541056 700644
rect 541072 700700 541136 700704
rect 541072 700644 541076 700700
rect 541076 700644 541132 700700
rect 541132 700644 541136 700700
rect 541072 700640 541136 700644
rect 541152 700700 541216 700704
rect 541152 700644 541156 700700
rect 541156 700644 541212 700700
rect 541212 700644 541216 700700
rect 541152 700640 541216 700644
rect 541232 700700 541296 700704
rect 541232 700644 541236 700700
rect 541236 700644 541292 700700
rect 541292 700644 541296 700700
rect 541232 700640 541296 700644
rect 541312 700700 541376 700704
rect 541312 700644 541316 700700
rect 541316 700644 541372 700700
rect 541372 700644 541376 700700
rect 541312 700640 541376 700644
rect 576832 700700 576896 700704
rect 576832 700644 576836 700700
rect 576836 700644 576892 700700
rect 576892 700644 576896 700700
rect 576832 700640 576896 700644
rect 576912 700700 576976 700704
rect 576912 700644 576916 700700
rect 576916 700644 576972 700700
rect 576972 700644 576976 700700
rect 576912 700640 576976 700644
rect 576992 700700 577056 700704
rect 576992 700644 576996 700700
rect 576996 700644 577052 700700
rect 577052 700644 577056 700700
rect 576992 700640 577056 700644
rect 577072 700700 577136 700704
rect 577072 700644 577076 700700
rect 577076 700644 577132 700700
rect 577132 700644 577136 700700
rect 577072 700640 577136 700644
rect 577152 700700 577216 700704
rect 577152 700644 577156 700700
rect 577156 700644 577212 700700
rect 577212 700644 577216 700700
rect 577152 700640 577216 700644
rect 577232 700700 577296 700704
rect 577232 700644 577236 700700
rect 577236 700644 577292 700700
rect 577292 700644 577296 700700
rect 577232 700640 577296 700644
rect 577312 700700 577376 700704
rect 577312 700644 577316 700700
rect 577316 700644 577372 700700
rect 577372 700644 577376 700700
rect 577312 700640 577376 700644
rect 18832 700156 18896 700160
rect 18832 700100 18836 700156
rect 18836 700100 18892 700156
rect 18892 700100 18896 700156
rect 18832 700096 18896 700100
rect 18912 700156 18976 700160
rect 18912 700100 18916 700156
rect 18916 700100 18972 700156
rect 18972 700100 18976 700156
rect 18912 700096 18976 700100
rect 18992 700156 19056 700160
rect 18992 700100 18996 700156
rect 18996 700100 19052 700156
rect 19052 700100 19056 700156
rect 18992 700096 19056 700100
rect 19072 700156 19136 700160
rect 19072 700100 19076 700156
rect 19076 700100 19132 700156
rect 19132 700100 19136 700156
rect 19072 700096 19136 700100
rect 19152 700156 19216 700160
rect 19152 700100 19156 700156
rect 19156 700100 19212 700156
rect 19212 700100 19216 700156
rect 19152 700096 19216 700100
rect 19232 700156 19296 700160
rect 19232 700100 19236 700156
rect 19236 700100 19292 700156
rect 19292 700100 19296 700156
rect 19232 700096 19296 700100
rect 19312 700156 19376 700160
rect 19312 700100 19316 700156
rect 19316 700100 19372 700156
rect 19372 700100 19376 700156
rect 19312 700096 19376 700100
rect 54832 700156 54896 700160
rect 54832 700100 54836 700156
rect 54836 700100 54892 700156
rect 54892 700100 54896 700156
rect 54832 700096 54896 700100
rect 54912 700156 54976 700160
rect 54912 700100 54916 700156
rect 54916 700100 54972 700156
rect 54972 700100 54976 700156
rect 54912 700096 54976 700100
rect 54992 700156 55056 700160
rect 54992 700100 54996 700156
rect 54996 700100 55052 700156
rect 55052 700100 55056 700156
rect 54992 700096 55056 700100
rect 55072 700156 55136 700160
rect 55072 700100 55076 700156
rect 55076 700100 55132 700156
rect 55132 700100 55136 700156
rect 55072 700096 55136 700100
rect 55152 700156 55216 700160
rect 55152 700100 55156 700156
rect 55156 700100 55212 700156
rect 55212 700100 55216 700156
rect 55152 700096 55216 700100
rect 55232 700156 55296 700160
rect 55232 700100 55236 700156
rect 55236 700100 55292 700156
rect 55292 700100 55296 700156
rect 55232 700096 55296 700100
rect 55312 700156 55376 700160
rect 55312 700100 55316 700156
rect 55316 700100 55372 700156
rect 55372 700100 55376 700156
rect 55312 700096 55376 700100
rect 90832 700156 90896 700160
rect 90832 700100 90836 700156
rect 90836 700100 90892 700156
rect 90892 700100 90896 700156
rect 90832 700096 90896 700100
rect 90912 700156 90976 700160
rect 90912 700100 90916 700156
rect 90916 700100 90972 700156
rect 90972 700100 90976 700156
rect 90912 700096 90976 700100
rect 90992 700156 91056 700160
rect 90992 700100 90996 700156
rect 90996 700100 91052 700156
rect 91052 700100 91056 700156
rect 90992 700096 91056 700100
rect 91072 700156 91136 700160
rect 91072 700100 91076 700156
rect 91076 700100 91132 700156
rect 91132 700100 91136 700156
rect 91072 700096 91136 700100
rect 91152 700156 91216 700160
rect 91152 700100 91156 700156
rect 91156 700100 91212 700156
rect 91212 700100 91216 700156
rect 91152 700096 91216 700100
rect 91232 700156 91296 700160
rect 91232 700100 91236 700156
rect 91236 700100 91292 700156
rect 91292 700100 91296 700156
rect 91232 700096 91296 700100
rect 91312 700156 91376 700160
rect 91312 700100 91316 700156
rect 91316 700100 91372 700156
rect 91372 700100 91376 700156
rect 91312 700096 91376 700100
rect 126832 700156 126896 700160
rect 126832 700100 126836 700156
rect 126836 700100 126892 700156
rect 126892 700100 126896 700156
rect 126832 700096 126896 700100
rect 126912 700156 126976 700160
rect 126912 700100 126916 700156
rect 126916 700100 126972 700156
rect 126972 700100 126976 700156
rect 126912 700096 126976 700100
rect 126992 700156 127056 700160
rect 126992 700100 126996 700156
rect 126996 700100 127052 700156
rect 127052 700100 127056 700156
rect 126992 700096 127056 700100
rect 127072 700156 127136 700160
rect 127072 700100 127076 700156
rect 127076 700100 127132 700156
rect 127132 700100 127136 700156
rect 127072 700096 127136 700100
rect 127152 700156 127216 700160
rect 127152 700100 127156 700156
rect 127156 700100 127212 700156
rect 127212 700100 127216 700156
rect 127152 700096 127216 700100
rect 127232 700156 127296 700160
rect 127232 700100 127236 700156
rect 127236 700100 127292 700156
rect 127292 700100 127296 700156
rect 127232 700096 127296 700100
rect 127312 700156 127376 700160
rect 127312 700100 127316 700156
rect 127316 700100 127372 700156
rect 127372 700100 127376 700156
rect 127312 700096 127376 700100
rect 162832 700156 162896 700160
rect 162832 700100 162836 700156
rect 162836 700100 162892 700156
rect 162892 700100 162896 700156
rect 162832 700096 162896 700100
rect 162912 700156 162976 700160
rect 162912 700100 162916 700156
rect 162916 700100 162972 700156
rect 162972 700100 162976 700156
rect 162912 700096 162976 700100
rect 162992 700156 163056 700160
rect 162992 700100 162996 700156
rect 162996 700100 163052 700156
rect 163052 700100 163056 700156
rect 162992 700096 163056 700100
rect 163072 700156 163136 700160
rect 163072 700100 163076 700156
rect 163076 700100 163132 700156
rect 163132 700100 163136 700156
rect 163072 700096 163136 700100
rect 163152 700156 163216 700160
rect 163152 700100 163156 700156
rect 163156 700100 163212 700156
rect 163212 700100 163216 700156
rect 163152 700096 163216 700100
rect 163232 700156 163296 700160
rect 163232 700100 163236 700156
rect 163236 700100 163292 700156
rect 163292 700100 163296 700156
rect 163232 700096 163296 700100
rect 163312 700156 163376 700160
rect 163312 700100 163316 700156
rect 163316 700100 163372 700156
rect 163372 700100 163376 700156
rect 163312 700096 163376 700100
rect 198832 700156 198896 700160
rect 198832 700100 198836 700156
rect 198836 700100 198892 700156
rect 198892 700100 198896 700156
rect 198832 700096 198896 700100
rect 198912 700156 198976 700160
rect 198912 700100 198916 700156
rect 198916 700100 198972 700156
rect 198972 700100 198976 700156
rect 198912 700096 198976 700100
rect 198992 700156 199056 700160
rect 198992 700100 198996 700156
rect 198996 700100 199052 700156
rect 199052 700100 199056 700156
rect 198992 700096 199056 700100
rect 199072 700156 199136 700160
rect 199072 700100 199076 700156
rect 199076 700100 199132 700156
rect 199132 700100 199136 700156
rect 199072 700096 199136 700100
rect 199152 700156 199216 700160
rect 199152 700100 199156 700156
rect 199156 700100 199212 700156
rect 199212 700100 199216 700156
rect 199152 700096 199216 700100
rect 199232 700156 199296 700160
rect 199232 700100 199236 700156
rect 199236 700100 199292 700156
rect 199292 700100 199296 700156
rect 199232 700096 199296 700100
rect 199312 700156 199376 700160
rect 199312 700100 199316 700156
rect 199316 700100 199372 700156
rect 199372 700100 199376 700156
rect 199312 700096 199376 700100
rect 234832 700156 234896 700160
rect 234832 700100 234836 700156
rect 234836 700100 234892 700156
rect 234892 700100 234896 700156
rect 234832 700096 234896 700100
rect 234912 700156 234976 700160
rect 234912 700100 234916 700156
rect 234916 700100 234972 700156
rect 234972 700100 234976 700156
rect 234912 700096 234976 700100
rect 234992 700156 235056 700160
rect 234992 700100 234996 700156
rect 234996 700100 235052 700156
rect 235052 700100 235056 700156
rect 234992 700096 235056 700100
rect 235072 700156 235136 700160
rect 235072 700100 235076 700156
rect 235076 700100 235132 700156
rect 235132 700100 235136 700156
rect 235072 700096 235136 700100
rect 235152 700156 235216 700160
rect 235152 700100 235156 700156
rect 235156 700100 235212 700156
rect 235212 700100 235216 700156
rect 235152 700096 235216 700100
rect 235232 700156 235296 700160
rect 235232 700100 235236 700156
rect 235236 700100 235292 700156
rect 235292 700100 235296 700156
rect 235232 700096 235296 700100
rect 235312 700156 235376 700160
rect 235312 700100 235316 700156
rect 235316 700100 235372 700156
rect 235372 700100 235376 700156
rect 235312 700096 235376 700100
rect 270832 700156 270896 700160
rect 270832 700100 270836 700156
rect 270836 700100 270892 700156
rect 270892 700100 270896 700156
rect 270832 700096 270896 700100
rect 270912 700156 270976 700160
rect 270912 700100 270916 700156
rect 270916 700100 270972 700156
rect 270972 700100 270976 700156
rect 270912 700096 270976 700100
rect 270992 700156 271056 700160
rect 270992 700100 270996 700156
rect 270996 700100 271052 700156
rect 271052 700100 271056 700156
rect 270992 700096 271056 700100
rect 271072 700156 271136 700160
rect 271072 700100 271076 700156
rect 271076 700100 271132 700156
rect 271132 700100 271136 700156
rect 271072 700096 271136 700100
rect 271152 700156 271216 700160
rect 271152 700100 271156 700156
rect 271156 700100 271212 700156
rect 271212 700100 271216 700156
rect 271152 700096 271216 700100
rect 271232 700156 271296 700160
rect 271232 700100 271236 700156
rect 271236 700100 271292 700156
rect 271292 700100 271296 700156
rect 271232 700096 271296 700100
rect 271312 700156 271376 700160
rect 271312 700100 271316 700156
rect 271316 700100 271372 700156
rect 271372 700100 271376 700156
rect 271312 700096 271376 700100
rect 306832 700156 306896 700160
rect 306832 700100 306836 700156
rect 306836 700100 306892 700156
rect 306892 700100 306896 700156
rect 306832 700096 306896 700100
rect 306912 700156 306976 700160
rect 306912 700100 306916 700156
rect 306916 700100 306972 700156
rect 306972 700100 306976 700156
rect 306912 700096 306976 700100
rect 306992 700156 307056 700160
rect 306992 700100 306996 700156
rect 306996 700100 307052 700156
rect 307052 700100 307056 700156
rect 306992 700096 307056 700100
rect 307072 700156 307136 700160
rect 307072 700100 307076 700156
rect 307076 700100 307132 700156
rect 307132 700100 307136 700156
rect 307072 700096 307136 700100
rect 307152 700156 307216 700160
rect 307152 700100 307156 700156
rect 307156 700100 307212 700156
rect 307212 700100 307216 700156
rect 307152 700096 307216 700100
rect 307232 700156 307296 700160
rect 307232 700100 307236 700156
rect 307236 700100 307292 700156
rect 307292 700100 307296 700156
rect 307232 700096 307296 700100
rect 307312 700156 307376 700160
rect 307312 700100 307316 700156
rect 307316 700100 307372 700156
rect 307372 700100 307376 700156
rect 307312 700096 307376 700100
rect 342832 700156 342896 700160
rect 342832 700100 342836 700156
rect 342836 700100 342892 700156
rect 342892 700100 342896 700156
rect 342832 700096 342896 700100
rect 342912 700156 342976 700160
rect 342912 700100 342916 700156
rect 342916 700100 342972 700156
rect 342972 700100 342976 700156
rect 342912 700096 342976 700100
rect 342992 700156 343056 700160
rect 342992 700100 342996 700156
rect 342996 700100 343052 700156
rect 343052 700100 343056 700156
rect 342992 700096 343056 700100
rect 343072 700156 343136 700160
rect 343072 700100 343076 700156
rect 343076 700100 343132 700156
rect 343132 700100 343136 700156
rect 343072 700096 343136 700100
rect 343152 700156 343216 700160
rect 343152 700100 343156 700156
rect 343156 700100 343212 700156
rect 343212 700100 343216 700156
rect 343152 700096 343216 700100
rect 343232 700156 343296 700160
rect 343232 700100 343236 700156
rect 343236 700100 343292 700156
rect 343292 700100 343296 700156
rect 343232 700096 343296 700100
rect 343312 700156 343376 700160
rect 343312 700100 343316 700156
rect 343316 700100 343372 700156
rect 343372 700100 343376 700156
rect 343312 700096 343376 700100
rect 378832 700156 378896 700160
rect 378832 700100 378836 700156
rect 378836 700100 378892 700156
rect 378892 700100 378896 700156
rect 378832 700096 378896 700100
rect 378912 700156 378976 700160
rect 378912 700100 378916 700156
rect 378916 700100 378972 700156
rect 378972 700100 378976 700156
rect 378912 700096 378976 700100
rect 378992 700156 379056 700160
rect 378992 700100 378996 700156
rect 378996 700100 379052 700156
rect 379052 700100 379056 700156
rect 378992 700096 379056 700100
rect 379072 700156 379136 700160
rect 379072 700100 379076 700156
rect 379076 700100 379132 700156
rect 379132 700100 379136 700156
rect 379072 700096 379136 700100
rect 379152 700156 379216 700160
rect 379152 700100 379156 700156
rect 379156 700100 379212 700156
rect 379212 700100 379216 700156
rect 379152 700096 379216 700100
rect 379232 700156 379296 700160
rect 379232 700100 379236 700156
rect 379236 700100 379292 700156
rect 379292 700100 379296 700156
rect 379232 700096 379296 700100
rect 379312 700156 379376 700160
rect 379312 700100 379316 700156
rect 379316 700100 379372 700156
rect 379372 700100 379376 700156
rect 379312 700096 379376 700100
rect 414832 700156 414896 700160
rect 414832 700100 414836 700156
rect 414836 700100 414892 700156
rect 414892 700100 414896 700156
rect 414832 700096 414896 700100
rect 414912 700156 414976 700160
rect 414912 700100 414916 700156
rect 414916 700100 414972 700156
rect 414972 700100 414976 700156
rect 414912 700096 414976 700100
rect 414992 700156 415056 700160
rect 414992 700100 414996 700156
rect 414996 700100 415052 700156
rect 415052 700100 415056 700156
rect 414992 700096 415056 700100
rect 415072 700156 415136 700160
rect 415072 700100 415076 700156
rect 415076 700100 415132 700156
rect 415132 700100 415136 700156
rect 415072 700096 415136 700100
rect 415152 700156 415216 700160
rect 415152 700100 415156 700156
rect 415156 700100 415212 700156
rect 415212 700100 415216 700156
rect 415152 700096 415216 700100
rect 415232 700156 415296 700160
rect 415232 700100 415236 700156
rect 415236 700100 415292 700156
rect 415292 700100 415296 700156
rect 415232 700096 415296 700100
rect 415312 700156 415376 700160
rect 415312 700100 415316 700156
rect 415316 700100 415372 700156
rect 415372 700100 415376 700156
rect 415312 700096 415376 700100
rect 450832 700156 450896 700160
rect 450832 700100 450836 700156
rect 450836 700100 450892 700156
rect 450892 700100 450896 700156
rect 450832 700096 450896 700100
rect 450912 700156 450976 700160
rect 450912 700100 450916 700156
rect 450916 700100 450972 700156
rect 450972 700100 450976 700156
rect 450912 700096 450976 700100
rect 450992 700156 451056 700160
rect 450992 700100 450996 700156
rect 450996 700100 451052 700156
rect 451052 700100 451056 700156
rect 450992 700096 451056 700100
rect 451072 700156 451136 700160
rect 451072 700100 451076 700156
rect 451076 700100 451132 700156
rect 451132 700100 451136 700156
rect 451072 700096 451136 700100
rect 451152 700156 451216 700160
rect 451152 700100 451156 700156
rect 451156 700100 451212 700156
rect 451212 700100 451216 700156
rect 451152 700096 451216 700100
rect 451232 700156 451296 700160
rect 451232 700100 451236 700156
rect 451236 700100 451292 700156
rect 451292 700100 451296 700156
rect 451232 700096 451296 700100
rect 451312 700156 451376 700160
rect 451312 700100 451316 700156
rect 451316 700100 451372 700156
rect 451372 700100 451376 700156
rect 451312 700096 451376 700100
rect 486832 700156 486896 700160
rect 486832 700100 486836 700156
rect 486836 700100 486892 700156
rect 486892 700100 486896 700156
rect 486832 700096 486896 700100
rect 486912 700156 486976 700160
rect 486912 700100 486916 700156
rect 486916 700100 486972 700156
rect 486972 700100 486976 700156
rect 486912 700096 486976 700100
rect 486992 700156 487056 700160
rect 486992 700100 486996 700156
rect 486996 700100 487052 700156
rect 487052 700100 487056 700156
rect 486992 700096 487056 700100
rect 487072 700156 487136 700160
rect 487072 700100 487076 700156
rect 487076 700100 487132 700156
rect 487132 700100 487136 700156
rect 487072 700096 487136 700100
rect 487152 700156 487216 700160
rect 487152 700100 487156 700156
rect 487156 700100 487212 700156
rect 487212 700100 487216 700156
rect 487152 700096 487216 700100
rect 487232 700156 487296 700160
rect 487232 700100 487236 700156
rect 487236 700100 487292 700156
rect 487292 700100 487296 700156
rect 487232 700096 487296 700100
rect 487312 700156 487376 700160
rect 487312 700100 487316 700156
rect 487316 700100 487372 700156
rect 487372 700100 487376 700156
rect 487312 700096 487376 700100
rect 522832 700156 522896 700160
rect 522832 700100 522836 700156
rect 522836 700100 522892 700156
rect 522892 700100 522896 700156
rect 522832 700096 522896 700100
rect 522912 700156 522976 700160
rect 522912 700100 522916 700156
rect 522916 700100 522972 700156
rect 522972 700100 522976 700156
rect 522912 700096 522976 700100
rect 522992 700156 523056 700160
rect 522992 700100 522996 700156
rect 522996 700100 523052 700156
rect 523052 700100 523056 700156
rect 522992 700096 523056 700100
rect 523072 700156 523136 700160
rect 523072 700100 523076 700156
rect 523076 700100 523132 700156
rect 523132 700100 523136 700156
rect 523072 700096 523136 700100
rect 523152 700156 523216 700160
rect 523152 700100 523156 700156
rect 523156 700100 523212 700156
rect 523212 700100 523216 700156
rect 523152 700096 523216 700100
rect 523232 700156 523296 700160
rect 523232 700100 523236 700156
rect 523236 700100 523292 700156
rect 523292 700100 523296 700156
rect 523232 700096 523296 700100
rect 523312 700156 523376 700160
rect 523312 700100 523316 700156
rect 523316 700100 523372 700156
rect 523372 700100 523376 700156
rect 523312 700096 523376 700100
rect 558832 700156 558896 700160
rect 558832 700100 558836 700156
rect 558836 700100 558892 700156
rect 558892 700100 558896 700156
rect 558832 700096 558896 700100
rect 558912 700156 558976 700160
rect 558912 700100 558916 700156
rect 558916 700100 558972 700156
rect 558972 700100 558976 700156
rect 558912 700096 558976 700100
rect 558992 700156 559056 700160
rect 558992 700100 558996 700156
rect 558996 700100 559052 700156
rect 559052 700100 559056 700156
rect 558992 700096 559056 700100
rect 559072 700156 559136 700160
rect 559072 700100 559076 700156
rect 559076 700100 559132 700156
rect 559132 700100 559136 700156
rect 559072 700096 559136 700100
rect 559152 700156 559216 700160
rect 559152 700100 559156 700156
rect 559156 700100 559212 700156
rect 559212 700100 559216 700156
rect 559152 700096 559216 700100
rect 559232 700156 559296 700160
rect 559232 700100 559236 700156
rect 559236 700100 559292 700156
rect 559292 700100 559296 700156
rect 559232 700096 559296 700100
rect 559312 700156 559376 700160
rect 559312 700100 559316 700156
rect 559316 700100 559372 700156
rect 559372 700100 559376 700156
rect 559312 700096 559376 700100
rect 269068 699756 269132 699820
rect 36832 699612 36896 699616
rect 36832 699556 36836 699612
rect 36836 699556 36892 699612
rect 36892 699556 36896 699612
rect 36832 699552 36896 699556
rect 36912 699612 36976 699616
rect 36912 699556 36916 699612
rect 36916 699556 36972 699612
rect 36972 699556 36976 699612
rect 36912 699552 36976 699556
rect 36992 699612 37056 699616
rect 36992 699556 36996 699612
rect 36996 699556 37052 699612
rect 37052 699556 37056 699612
rect 36992 699552 37056 699556
rect 37072 699612 37136 699616
rect 37072 699556 37076 699612
rect 37076 699556 37132 699612
rect 37132 699556 37136 699612
rect 37072 699552 37136 699556
rect 37152 699612 37216 699616
rect 37152 699556 37156 699612
rect 37156 699556 37212 699612
rect 37212 699556 37216 699612
rect 37152 699552 37216 699556
rect 37232 699612 37296 699616
rect 37232 699556 37236 699612
rect 37236 699556 37292 699612
rect 37292 699556 37296 699612
rect 37232 699552 37296 699556
rect 37312 699612 37376 699616
rect 37312 699556 37316 699612
rect 37316 699556 37372 699612
rect 37372 699556 37376 699612
rect 37312 699552 37376 699556
rect 72832 699612 72896 699616
rect 72832 699556 72836 699612
rect 72836 699556 72892 699612
rect 72892 699556 72896 699612
rect 72832 699552 72896 699556
rect 72912 699612 72976 699616
rect 72912 699556 72916 699612
rect 72916 699556 72972 699612
rect 72972 699556 72976 699612
rect 72912 699552 72976 699556
rect 72992 699612 73056 699616
rect 72992 699556 72996 699612
rect 72996 699556 73052 699612
rect 73052 699556 73056 699612
rect 72992 699552 73056 699556
rect 73072 699612 73136 699616
rect 73072 699556 73076 699612
rect 73076 699556 73132 699612
rect 73132 699556 73136 699612
rect 73072 699552 73136 699556
rect 73152 699612 73216 699616
rect 73152 699556 73156 699612
rect 73156 699556 73212 699612
rect 73212 699556 73216 699612
rect 73152 699552 73216 699556
rect 73232 699612 73296 699616
rect 73232 699556 73236 699612
rect 73236 699556 73292 699612
rect 73292 699556 73296 699612
rect 73232 699552 73296 699556
rect 73312 699612 73376 699616
rect 73312 699556 73316 699612
rect 73316 699556 73372 699612
rect 73372 699556 73376 699612
rect 73312 699552 73376 699556
rect 108832 699612 108896 699616
rect 108832 699556 108836 699612
rect 108836 699556 108892 699612
rect 108892 699556 108896 699612
rect 108832 699552 108896 699556
rect 108912 699612 108976 699616
rect 108912 699556 108916 699612
rect 108916 699556 108972 699612
rect 108972 699556 108976 699612
rect 108912 699552 108976 699556
rect 108992 699612 109056 699616
rect 108992 699556 108996 699612
rect 108996 699556 109052 699612
rect 109052 699556 109056 699612
rect 108992 699552 109056 699556
rect 109072 699612 109136 699616
rect 109072 699556 109076 699612
rect 109076 699556 109132 699612
rect 109132 699556 109136 699612
rect 109072 699552 109136 699556
rect 109152 699612 109216 699616
rect 109152 699556 109156 699612
rect 109156 699556 109212 699612
rect 109212 699556 109216 699612
rect 109152 699552 109216 699556
rect 109232 699612 109296 699616
rect 109232 699556 109236 699612
rect 109236 699556 109292 699612
rect 109292 699556 109296 699612
rect 109232 699552 109296 699556
rect 109312 699612 109376 699616
rect 109312 699556 109316 699612
rect 109316 699556 109372 699612
rect 109372 699556 109376 699612
rect 109312 699552 109376 699556
rect 144832 699612 144896 699616
rect 144832 699556 144836 699612
rect 144836 699556 144892 699612
rect 144892 699556 144896 699612
rect 144832 699552 144896 699556
rect 144912 699612 144976 699616
rect 144912 699556 144916 699612
rect 144916 699556 144972 699612
rect 144972 699556 144976 699612
rect 144912 699552 144976 699556
rect 144992 699612 145056 699616
rect 144992 699556 144996 699612
rect 144996 699556 145052 699612
rect 145052 699556 145056 699612
rect 144992 699552 145056 699556
rect 145072 699612 145136 699616
rect 145072 699556 145076 699612
rect 145076 699556 145132 699612
rect 145132 699556 145136 699612
rect 145072 699552 145136 699556
rect 145152 699612 145216 699616
rect 145152 699556 145156 699612
rect 145156 699556 145212 699612
rect 145212 699556 145216 699612
rect 145152 699552 145216 699556
rect 145232 699612 145296 699616
rect 145232 699556 145236 699612
rect 145236 699556 145292 699612
rect 145292 699556 145296 699612
rect 145232 699552 145296 699556
rect 145312 699612 145376 699616
rect 145312 699556 145316 699612
rect 145316 699556 145372 699612
rect 145372 699556 145376 699612
rect 145312 699552 145376 699556
rect 180832 699612 180896 699616
rect 180832 699556 180836 699612
rect 180836 699556 180892 699612
rect 180892 699556 180896 699612
rect 180832 699552 180896 699556
rect 180912 699612 180976 699616
rect 180912 699556 180916 699612
rect 180916 699556 180972 699612
rect 180972 699556 180976 699612
rect 180912 699552 180976 699556
rect 180992 699612 181056 699616
rect 180992 699556 180996 699612
rect 180996 699556 181052 699612
rect 181052 699556 181056 699612
rect 180992 699552 181056 699556
rect 181072 699612 181136 699616
rect 181072 699556 181076 699612
rect 181076 699556 181132 699612
rect 181132 699556 181136 699612
rect 181072 699552 181136 699556
rect 181152 699612 181216 699616
rect 181152 699556 181156 699612
rect 181156 699556 181212 699612
rect 181212 699556 181216 699612
rect 181152 699552 181216 699556
rect 181232 699612 181296 699616
rect 181232 699556 181236 699612
rect 181236 699556 181292 699612
rect 181292 699556 181296 699612
rect 181232 699552 181296 699556
rect 181312 699612 181376 699616
rect 181312 699556 181316 699612
rect 181316 699556 181372 699612
rect 181372 699556 181376 699612
rect 181312 699552 181376 699556
rect 216832 699612 216896 699616
rect 216832 699556 216836 699612
rect 216836 699556 216892 699612
rect 216892 699556 216896 699612
rect 216832 699552 216896 699556
rect 216912 699612 216976 699616
rect 216912 699556 216916 699612
rect 216916 699556 216972 699612
rect 216972 699556 216976 699612
rect 216912 699552 216976 699556
rect 216992 699612 217056 699616
rect 216992 699556 216996 699612
rect 216996 699556 217052 699612
rect 217052 699556 217056 699612
rect 216992 699552 217056 699556
rect 217072 699612 217136 699616
rect 217072 699556 217076 699612
rect 217076 699556 217132 699612
rect 217132 699556 217136 699612
rect 217072 699552 217136 699556
rect 217152 699612 217216 699616
rect 217152 699556 217156 699612
rect 217156 699556 217212 699612
rect 217212 699556 217216 699612
rect 217152 699552 217216 699556
rect 217232 699612 217296 699616
rect 217232 699556 217236 699612
rect 217236 699556 217292 699612
rect 217292 699556 217296 699612
rect 217232 699552 217296 699556
rect 217312 699612 217376 699616
rect 217312 699556 217316 699612
rect 217316 699556 217372 699612
rect 217372 699556 217376 699612
rect 217312 699552 217376 699556
rect 252832 699612 252896 699616
rect 252832 699556 252836 699612
rect 252836 699556 252892 699612
rect 252892 699556 252896 699612
rect 252832 699552 252896 699556
rect 252912 699612 252976 699616
rect 252912 699556 252916 699612
rect 252916 699556 252972 699612
rect 252972 699556 252976 699612
rect 252912 699552 252976 699556
rect 252992 699612 253056 699616
rect 252992 699556 252996 699612
rect 252996 699556 253052 699612
rect 253052 699556 253056 699612
rect 252992 699552 253056 699556
rect 253072 699612 253136 699616
rect 253072 699556 253076 699612
rect 253076 699556 253132 699612
rect 253132 699556 253136 699612
rect 253072 699552 253136 699556
rect 253152 699612 253216 699616
rect 253152 699556 253156 699612
rect 253156 699556 253212 699612
rect 253212 699556 253216 699612
rect 253152 699552 253216 699556
rect 253232 699612 253296 699616
rect 253232 699556 253236 699612
rect 253236 699556 253292 699612
rect 253292 699556 253296 699612
rect 253232 699552 253296 699556
rect 253312 699612 253376 699616
rect 253312 699556 253316 699612
rect 253316 699556 253372 699612
rect 253372 699556 253376 699612
rect 253312 699552 253376 699556
rect 288832 699612 288896 699616
rect 288832 699556 288836 699612
rect 288836 699556 288892 699612
rect 288892 699556 288896 699612
rect 288832 699552 288896 699556
rect 288912 699612 288976 699616
rect 288912 699556 288916 699612
rect 288916 699556 288972 699612
rect 288972 699556 288976 699612
rect 288912 699552 288976 699556
rect 288992 699612 289056 699616
rect 288992 699556 288996 699612
rect 288996 699556 289052 699612
rect 289052 699556 289056 699612
rect 288992 699552 289056 699556
rect 289072 699612 289136 699616
rect 289072 699556 289076 699612
rect 289076 699556 289132 699612
rect 289132 699556 289136 699612
rect 289072 699552 289136 699556
rect 289152 699612 289216 699616
rect 289152 699556 289156 699612
rect 289156 699556 289212 699612
rect 289212 699556 289216 699612
rect 289152 699552 289216 699556
rect 289232 699612 289296 699616
rect 289232 699556 289236 699612
rect 289236 699556 289292 699612
rect 289292 699556 289296 699612
rect 289232 699552 289296 699556
rect 289312 699612 289376 699616
rect 289312 699556 289316 699612
rect 289316 699556 289372 699612
rect 289372 699556 289376 699612
rect 289312 699552 289376 699556
rect 324832 699612 324896 699616
rect 324832 699556 324836 699612
rect 324836 699556 324892 699612
rect 324892 699556 324896 699612
rect 324832 699552 324896 699556
rect 324912 699612 324976 699616
rect 324912 699556 324916 699612
rect 324916 699556 324972 699612
rect 324972 699556 324976 699612
rect 324912 699552 324976 699556
rect 324992 699612 325056 699616
rect 324992 699556 324996 699612
rect 324996 699556 325052 699612
rect 325052 699556 325056 699612
rect 324992 699552 325056 699556
rect 325072 699612 325136 699616
rect 325072 699556 325076 699612
rect 325076 699556 325132 699612
rect 325132 699556 325136 699612
rect 325072 699552 325136 699556
rect 325152 699612 325216 699616
rect 325152 699556 325156 699612
rect 325156 699556 325212 699612
rect 325212 699556 325216 699612
rect 325152 699552 325216 699556
rect 325232 699612 325296 699616
rect 325232 699556 325236 699612
rect 325236 699556 325292 699612
rect 325292 699556 325296 699612
rect 325232 699552 325296 699556
rect 325312 699612 325376 699616
rect 325312 699556 325316 699612
rect 325316 699556 325372 699612
rect 325372 699556 325376 699612
rect 325312 699552 325376 699556
rect 360832 699612 360896 699616
rect 360832 699556 360836 699612
rect 360836 699556 360892 699612
rect 360892 699556 360896 699612
rect 360832 699552 360896 699556
rect 360912 699612 360976 699616
rect 360912 699556 360916 699612
rect 360916 699556 360972 699612
rect 360972 699556 360976 699612
rect 360912 699552 360976 699556
rect 360992 699612 361056 699616
rect 360992 699556 360996 699612
rect 360996 699556 361052 699612
rect 361052 699556 361056 699612
rect 360992 699552 361056 699556
rect 361072 699612 361136 699616
rect 361072 699556 361076 699612
rect 361076 699556 361132 699612
rect 361132 699556 361136 699612
rect 361072 699552 361136 699556
rect 361152 699612 361216 699616
rect 361152 699556 361156 699612
rect 361156 699556 361212 699612
rect 361212 699556 361216 699612
rect 361152 699552 361216 699556
rect 361232 699612 361296 699616
rect 361232 699556 361236 699612
rect 361236 699556 361292 699612
rect 361292 699556 361296 699612
rect 361232 699552 361296 699556
rect 361312 699612 361376 699616
rect 361312 699556 361316 699612
rect 361316 699556 361372 699612
rect 361372 699556 361376 699612
rect 361312 699552 361376 699556
rect 396832 699612 396896 699616
rect 396832 699556 396836 699612
rect 396836 699556 396892 699612
rect 396892 699556 396896 699612
rect 396832 699552 396896 699556
rect 396912 699612 396976 699616
rect 396912 699556 396916 699612
rect 396916 699556 396972 699612
rect 396972 699556 396976 699612
rect 396912 699552 396976 699556
rect 396992 699612 397056 699616
rect 396992 699556 396996 699612
rect 396996 699556 397052 699612
rect 397052 699556 397056 699612
rect 396992 699552 397056 699556
rect 397072 699612 397136 699616
rect 397072 699556 397076 699612
rect 397076 699556 397132 699612
rect 397132 699556 397136 699612
rect 397072 699552 397136 699556
rect 397152 699612 397216 699616
rect 397152 699556 397156 699612
rect 397156 699556 397212 699612
rect 397212 699556 397216 699612
rect 397152 699552 397216 699556
rect 397232 699612 397296 699616
rect 397232 699556 397236 699612
rect 397236 699556 397292 699612
rect 397292 699556 397296 699612
rect 397232 699552 397296 699556
rect 397312 699612 397376 699616
rect 397312 699556 397316 699612
rect 397316 699556 397372 699612
rect 397372 699556 397376 699612
rect 397312 699552 397376 699556
rect 432832 699612 432896 699616
rect 432832 699556 432836 699612
rect 432836 699556 432892 699612
rect 432892 699556 432896 699612
rect 432832 699552 432896 699556
rect 432912 699612 432976 699616
rect 432912 699556 432916 699612
rect 432916 699556 432972 699612
rect 432972 699556 432976 699612
rect 432912 699552 432976 699556
rect 432992 699612 433056 699616
rect 432992 699556 432996 699612
rect 432996 699556 433052 699612
rect 433052 699556 433056 699612
rect 432992 699552 433056 699556
rect 433072 699612 433136 699616
rect 433072 699556 433076 699612
rect 433076 699556 433132 699612
rect 433132 699556 433136 699612
rect 433072 699552 433136 699556
rect 433152 699612 433216 699616
rect 433152 699556 433156 699612
rect 433156 699556 433212 699612
rect 433212 699556 433216 699612
rect 433152 699552 433216 699556
rect 433232 699612 433296 699616
rect 433232 699556 433236 699612
rect 433236 699556 433292 699612
rect 433292 699556 433296 699612
rect 433232 699552 433296 699556
rect 433312 699612 433376 699616
rect 433312 699556 433316 699612
rect 433316 699556 433372 699612
rect 433372 699556 433376 699612
rect 433312 699552 433376 699556
rect 468832 699612 468896 699616
rect 468832 699556 468836 699612
rect 468836 699556 468892 699612
rect 468892 699556 468896 699612
rect 468832 699552 468896 699556
rect 468912 699612 468976 699616
rect 468912 699556 468916 699612
rect 468916 699556 468972 699612
rect 468972 699556 468976 699612
rect 468912 699552 468976 699556
rect 468992 699612 469056 699616
rect 468992 699556 468996 699612
rect 468996 699556 469052 699612
rect 469052 699556 469056 699612
rect 468992 699552 469056 699556
rect 469072 699612 469136 699616
rect 469072 699556 469076 699612
rect 469076 699556 469132 699612
rect 469132 699556 469136 699612
rect 469072 699552 469136 699556
rect 469152 699612 469216 699616
rect 469152 699556 469156 699612
rect 469156 699556 469212 699612
rect 469212 699556 469216 699612
rect 469152 699552 469216 699556
rect 469232 699612 469296 699616
rect 469232 699556 469236 699612
rect 469236 699556 469292 699612
rect 469292 699556 469296 699612
rect 469232 699552 469296 699556
rect 469312 699612 469376 699616
rect 469312 699556 469316 699612
rect 469316 699556 469372 699612
rect 469372 699556 469376 699612
rect 469312 699552 469376 699556
rect 504832 699612 504896 699616
rect 504832 699556 504836 699612
rect 504836 699556 504892 699612
rect 504892 699556 504896 699612
rect 504832 699552 504896 699556
rect 504912 699612 504976 699616
rect 504912 699556 504916 699612
rect 504916 699556 504972 699612
rect 504972 699556 504976 699612
rect 504912 699552 504976 699556
rect 504992 699612 505056 699616
rect 504992 699556 504996 699612
rect 504996 699556 505052 699612
rect 505052 699556 505056 699612
rect 504992 699552 505056 699556
rect 505072 699612 505136 699616
rect 505072 699556 505076 699612
rect 505076 699556 505132 699612
rect 505132 699556 505136 699612
rect 505072 699552 505136 699556
rect 505152 699612 505216 699616
rect 505152 699556 505156 699612
rect 505156 699556 505212 699612
rect 505212 699556 505216 699612
rect 505152 699552 505216 699556
rect 505232 699612 505296 699616
rect 505232 699556 505236 699612
rect 505236 699556 505292 699612
rect 505292 699556 505296 699612
rect 505232 699552 505296 699556
rect 505312 699612 505376 699616
rect 505312 699556 505316 699612
rect 505316 699556 505372 699612
rect 505372 699556 505376 699612
rect 505312 699552 505376 699556
rect 540832 699612 540896 699616
rect 540832 699556 540836 699612
rect 540836 699556 540892 699612
rect 540892 699556 540896 699612
rect 540832 699552 540896 699556
rect 540912 699612 540976 699616
rect 540912 699556 540916 699612
rect 540916 699556 540972 699612
rect 540972 699556 540976 699612
rect 540912 699552 540976 699556
rect 540992 699612 541056 699616
rect 540992 699556 540996 699612
rect 540996 699556 541052 699612
rect 541052 699556 541056 699612
rect 540992 699552 541056 699556
rect 541072 699612 541136 699616
rect 541072 699556 541076 699612
rect 541076 699556 541132 699612
rect 541132 699556 541136 699612
rect 541072 699552 541136 699556
rect 541152 699612 541216 699616
rect 541152 699556 541156 699612
rect 541156 699556 541212 699612
rect 541212 699556 541216 699612
rect 541152 699552 541216 699556
rect 541232 699612 541296 699616
rect 541232 699556 541236 699612
rect 541236 699556 541292 699612
rect 541292 699556 541296 699612
rect 541232 699552 541296 699556
rect 541312 699612 541376 699616
rect 541312 699556 541316 699612
rect 541316 699556 541372 699612
rect 541372 699556 541376 699612
rect 541312 699552 541376 699556
rect 576832 699612 576896 699616
rect 576832 699556 576836 699612
rect 576836 699556 576892 699612
rect 576892 699556 576896 699612
rect 576832 699552 576896 699556
rect 576912 699612 576976 699616
rect 576912 699556 576916 699612
rect 576916 699556 576972 699612
rect 576972 699556 576976 699612
rect 576912 699552 576976 699556
rect 576992 699612 577056 699616
rect 576992 699556 576996 699612
rect 576996 699556 577052 699612
rect 577052 699556 577056 699612
rect 576992 699552 577056 699556
rect 577072 699612 577136 699616
rect 577072 699556 577076 699612
rect 577076 699556 577132 699612
rect 577132 699556 577136 699612
rect 577072 699552 577136 699556
rect 577152 699612 577216 699616
rect 577152 699556 577156 699612
rect 577156 699556 577212 699612
rect 577212 699556 577216 699612
rect 577152 699552 577216 699556
rect 577232 699612 577296 699616
rect 577232 699556 577236 699612
rect 577236 699556 577292 699612
rect 577292 699556 577296 699612
rect 577232 699552 577296 699556
rect 577312 699612 577376 699616
rect 577312 699556 577316 699612
rect 577316 699556 577372 699612
rect 577372 699556 577376 699612
rect 577312 699552 577376 699556
rect 269068 699484 269132 699548
rect 18832 699068 18896 699072
rect 18832 699012 18836 699068
rect 18836 699012 18892 699068
rect 18892 699012 18896 699068
rect 18832 699008 18896 699012
rect 18912 699068 18976 699072
rect 18912 699012 18916 699068
rect 18916 699012 18972 699068
rect 18972 699012 18976 699068
rect 18912 699008 18976 699012
rect 18992 699068 19056 699072
rect 18992 699012 18996 699068
rect 18996 699012 19052 699068
rect 19052 699012 19056 699068
rect 18992 699008 19056 699012
rect 19072 699068 19136 699072
rect 19072 699012 19076 699068
rect 19076 699012 19132 699068
rect 19132 699012 19136 699068
rect 19072 699008 19136 699012
rect 19152 699068 19216 699072
rect 19152 699012 19156 699068
rect 19156 699012 19212 699068
rect 19212 699012 19216 699068
rect 19152 699008 19216 699012
rect 19232 699068 19296 699072
rect 19232 699012 19236 699068
rect 19236 699012 19292 699068
rect 19292 699012 19296 699068
rect 19232 699008 19296 699012
rect 19312 699068 19376 699072
rect 19312 699012 19316 699068
rect 19316 699012 19372 699068
rect 19372 699012 19376 699068
rect 19312 699008 19376 699012
rect 54832 699068 54896 699072
rect 54832 699012 54836 699068
rect 54836 699012 54892 699068
rect 54892 699012 54896 699068
rect 54832 699008 54896 699012
rect 54912 699068 54976 699072
rect 54912 699012 54916 699068
rect 54916 699012 54972 699068
rect 54972 699012 54976 699068
rect 54912 699008 54976 699012
rect 54992 699068 55056 699072
rect 54992 699012 54996 699068
rect 54996 699012 55052 699068
rect 55052 699012 55056 699068
rect 54992 699008 55056 699012
rect 55072 699068 55136 699072
rect 55072 699012 55076 699068
rect 55076 699012 55132 699068
rect 55132 699012 55136 699068
rect 55072 699008 55136 699012
rect 55152 699068 55216 699072
rect 55152 699012 55156 699068
rect 55156 699012 55212 699068
rect 55212 699012 55216 699068
rect 55152 699008 55216 699012
rect 55232 699068 55296 699072
rect 55232 699012 55236 699068
rect 55236 699012 55292 699068
rect 55292 699012 55296 699068
rect 55232 699008 55296 699012
rect 55312 699068 55376 699072
rect 55312 699012 55316 699068
rect 55316 699012 55372 699068
rect 55372 699012 55376 699068
rect 55312 699008 55376 699012
rect 90832 699068 90896 699072
rect 90832 699012 90836 699068
rect 90836 699012 90892 699068
rect 90892 699012 90896 699068
rect 90832 699008 90896 699012
rect 90912 699068 90976 699072
rect 90912 699012 90916 699068
rect 90916 699012 90972 699068
rect 90972 699012 90976 699068
rect 90912 699008 90976 699012
rect 90992 699068 91056 699072
rect 90992 699012 90996 699068
rect 90996 699012 91052 699068
rect 91052 699012 91056 699068
rect 90992 699008 91056 699012
rect 91072 699068 91136 699072
rect 91072 699012 91076 699068
rect 91076 699012 91132 699068
rect 91132 699012 91136 699068
rect 91072 699008 91136 699012
rect 91152 699068 91216 699072
rect 91152 699012 91156 699068
rect 91156 699012 91212 699068
rect 91212 699012 91216 699068
rect 91152 699008 91216 699012
rect 91232 699068 91296 699072
rect 91232 699012 91236 699068
rect 91236 699012 91292 699068
rect 91292 699012 91296 699068
rect 91232 699008 91296 699012
rect 91312 699068 91376 699072
rect 91312 699012 91316 699068
rect 91316 699012 91372 699068
rect 91372 699012 91376 699068
rect 91312 699008 91376 699012
rect 126832 699068 126896 699072
rect 126832 699012 126836 699068
rect 126836 699012 126892 699068
rect 126892 699012 126896 699068
rect 126832 699008 126896 699012
rect 126912 699068 126976 699072
rect 126912 699012 126916 699068
rect 126916 699012 126972 699068
rect 126972 699012 126976 699068
rect 126912 699008 126976 699012
rect 126992 699068 127056 699072
rect 126992 699012 126996 699068
rect 126996 699012 127052 699068
rect 127052 699012 127056 699068
rect 126992 699008 127056 699012
rect 127072 699068 127136 699072
rect 127072 699012 127076 699068
rect 127076 699012 127132 699068
rect 127132 699012 127136 699068
rect 127072 699008 127136 699012
rect 127152 699068 127216 699072
rect 127152 699012 127156 699068
rect 127156 699012 127212 699068
rect 127212 699012 127216 699068
rect 127152 699008 127216 699012
rect 127232 699068 127296 699072
rect 127232 699012 127236 699068
rect 127236 699012 127292 699068
rect 127292 699012 127296 699068
rect 127232 699008 127296 699012
rect 127312 699068 127376 699072
rect 127312 699012 127316 699068
rect 127316 699012 127372 699068
rect 127372 699012 127376 699068
rect 127312 699008 127376 699012
rect 162832 699068 162896 699072
rect 162832 699012 162836 699068
rect 162836 699012 162892 699068
rect 162892 699012 162896 699068
rect 162832 699008 162896 699012
rect 162912 699068 162976 699072
rect 162912 699012 162916 699068
rect 162916 699012 162972 699068
rect 162972 699012 162976 699068
rect 162912 699008 162976 699012
rect 162992 699068 163056 699072
rect 162992 699012 162996 699068
rect 162996 699012 163052 699068
rect 163052 699012 163056 699068
rect 162992 699008 163056 699012
rect 163072 699068 163136 699072
rect 163072 699012 163076 699068
rect 163076 699012 163132 699068
rect 163132 699012 163136 699068
rect 163072 699008 163136 699012
rect 163152 699068 163216 699072
rect 163152 699012 163156 699068
rect 163156 699012 163212 699068
rect 163212 699012 163216 699068
rect 163152 699008 163216 699012
rect 163232 699068 163296 699072
rect 163232 699012 163236 699068
rect 163236 699012 163292 699068
rect 163292 699012 163296 699068
rect 163232 699008 163296 699012
rect 163312 699068 163376 699072
rect 163312 699012 163316 699068
rect 163316 699012 163372 699068
rect 163372 699012 163376 699068
rect 163312 699008 163376 699012
rect 198832 699068 198896 699072
rect 198832 699012 198836 699068
rect 198836 699012 198892 699068
rect 198892 699012 198896 699068
rect 198832 699008 198896 699012
rect 198912 699068 198976 699072
rect 198912 699012 198916 699068
rect 198916 699012 198972 699068
rect 198972 699012 198976 699068
rect 198912 699008 198976 699012
rect 198992 699068 199056 699072
rect 198992 699012 198996 699068
rect 198996 699012 199052 699068
rect 199052 699012 199056 699068
rect 198992 699008 199056 699012
rect 199072 699068 199136 699072
rect 199072 699012 199076 699068
rect 199076 699012 199132 699068
rect 199132 699012 199136 699068
rect 199072 699008 199136 699012
rect 199152 699068 199216 699072
rect 199152 699012 199156 699068
rect 199156 699012 199212 699068
rect 199212 699012 199216 699068
rect 199152 699008 199216 699012
rect 199232 699068 199296 699072
rect 199232 699012 199236 699068
rect 199236 699012 199292 699068
rect 199292 699012 199296 699068
rect 199232 699008 199296 699012
rect 199312 699068 199376 699072
rect 199312 699012 199316 699068
rect 199316 699012 199372 699068
rect 199372 699012 199376 699068
rect 199312 699008 199376 699012
rect 234832 699068 234896 699072
rect 234832 699012 234836 699068
rect 234836 699012 234892 699068
rect 234892 699012 234896 699068
rect 234832 699008 234896 699012
rect 234912 699068 234976 699072
rect 234912 699012 234916 699068
rect 234916 699012 234972 699068
rect 234972 699012 234976 699068
rect 234912 699008 234976 699012
rect 234992 699068 235056 699072
rect 234992 699012 234996 699068
rect 234996 699012 235052 699068
rect 235052 699012 235056 699068
rect 234992 699008 235056 699012
rect 235072 699068 235136 699072
rect 235072 699012 235076 699068
rect 235076 699012 235132 699068
rect 235132 699012 235136 699068
rect 235072 699008 235136 699012
rect 235152 699068 235216 699072
rect 235152 699012 235156 699068
rect 235156 699012 235212 699068
rect 235212 699012 235216 699068
rect 235152 699008 235216 699012
rect 235232 699068 235296 699072
rect 235232 699012 235236 699068
rect 235236 699012 235292 699068
rect 235292 699012 235296 699068
rect 235232 699008 235296 699012
rect 235312 699068 235376 699072
rect 235312 699012 235316 699068
rect 235316 699012 235372 699068
rect 235372 699012 235376 699068
rect 235312 699008 235376 699012
rect 503484 699212 503548 699276
rect 270832 699068 270896 699072
rect 270832 699012 270836 699068
rect 270836 699012 270892 699068
rect 270892 699012 270896 699068
rect 270832 699008 270896 699012
rect 270912 699068 270976 699072
rect 270912 699012 270916 699068
rect 270916 699012 270972 699068
rect 270972 699012 270976 699068
rect 270912 699008 270976 699012
rect 270992 699068 271056 699072
rect 270992 699012 270996 699068
rect 270996 699012 271052 699068
rect 271052 699012 271056 699068
rect 270992 699008 271056 699012
rect 271072 699068 271136 699072
rect 271072 699012 271076 699068
rect 271076 699012 271132 699068
rect 271132 699012 271136 699068
rect 271072 699008 271136 699012
rect 271152 699068 271216 699072
rect 271152 699012 271156 699068
rect 271156 699012 271212 699068
rect 271212 699012 271216 699068
rect 271152 699008 271216 699012
rect 271232 699068 271296 699072
rect 271232 699012 271236 699068
rect 271236 699012 271292 699068
rect 271292 699012 271296 699068
rect 271232 699008 271296 699012
rect 271312 699068 271376 699072
rect 271312 699012 271316 699068
rect 271316 699012 271372 699068
rect 271372 699012 271376 699068
rect 271312 699008 271376 699012
rect 306832 699068 306896 699072
rect 306832 699012 306836 699068
rect 306836 699012 306892 699068
rect 306892 699012 306896 699068
rect 306832 699008 306896 699012
rect 306912 699068 306976 699072
rect 306912 699012 306916 699068
rect 306916 699012 306972 699068
rect 306972 699012 306976 699068
rect 306912 699008 306976 699012
rect 306992 699068 307056 699072
rect 306992 699012 306996 699068
rect 306996 699012 307052 699068
rect 307052 699012 307056 699068
rect 306992 699008 307056 699012
rect 307072 699068 307136 699072
rect 307072 699012 307076 699068
rect 307076 699012 307132 699068
rect 307132 699012 307136 699068
rect 307072 699008 307136 699012
rect 307152 699068 307216 699072
rect 307152 699012 307156 699068
rect 307156 699012 307212 699068
rect 307212 699012 307216 699068
rect 307152 699008 307216 699012
rect 307232 699068 307296 699072
rect 307232 699012 307236 699068
rect 307236 699012 307292 699068
rect 307292 699012 307296 699068
rect 307232 699008 307296 699012
rect 307312 699068 307376 699072
rect 307312 699012 307316 699068
rect 307316 699012 307372 699068
rect 307372 699012 307376 699068
rect 307312 699008 307376 699012
rect 342832 699068 342896 699072
rect 342832 699012 342836 699068
rect 342836 699012 342892 699068
rect 342892 699012 342896 699068
rect 342832 699008 342896 699012
rect 342912 699068 342976 699072
rect 342912 699012 342916 699068
rect 342916 699012 342972 699068
rect 342972 699012 342976 699068
rect 342912 699008 342976 699012
rect 342992 699068 343056 699072
rect 342992 699012 342996 699068
rect 342996 699012 343052 699068
rect 343052 699012 343056 699068
rect 342992 699008 343056 699012
rect 343072 699068 343136 699072
rect 343072 699012 343076 699068
rect 343076 699012 343132 699068
rect 343132 699012 343136 699068
rect 343072 699008 343136 699012
rect 343152 699068 343216 699072
rect 343152 699012 343156 699068
rect 343156 699012 343212 699068
rect 343212 699012 343216 699068
rect 343152 699008 343216 699012
rect 343232 699068 343296 699072
rect 343232 699012 343236 699068
rect 343236 699012 343292 699068
rect 343292 699012 343296 699068
rect 343232 699008 343296 699012
rect 343312 699068 343376 699072
rect 343312 699012 343316 699068
rect 343316 699012 343372 699068
rect 343372 699012 343376 699068
rect 343312 699008 343376 699012
rect 378832 699068 378896 699072
rect 378832 699012 378836 699068
rect 378836 699012 378892 699068
rect 378892 699012 378896 699068
rect 378832 699008 378896 699012
rect 378912 699068 378976 699072
rect 378912 699012 378916 699068
rect 378916 699012 378972 699068
rect 378972 699012 378976 699068
rect 378912 699008 378976 699012
rect 378992 699068 379056 699072
rect 378992 699012 378996 699068
rect 378996 699012 379052 699068
rect 379052 699012 379056 699068
rect 378992 699008 379056 699012
rect 379072 699068 379136 699072
rect 379072 699012 379076 699068
rect 379076 699012 379132 699068
rect 379132 699012 379136 699068
rect 379072 699008 379136 699012
rect 379152 699068 379216 699072
rect 379152 699012 379156 699068
rect 379156 699012 379212 699068
rect 379212 699012 379216 699068
rect 379152 699008 379216 699012
rect 379232 699068 379296 699072
rect 379232 699012 379236 699068
rect 379236 699012 379292 699068
rect 379292 699012 379296 699068
rect 379232 699008 379296 699012
rect 379312 699068 379376 699072
rect 379312 699012 379316 699068
rect 379316 699012 379372 699068
rect 379372 699012 379376 699068
rect 379312 699008 379376 699012
rect 414832 699068 414896 699072
rect 414832 699012 414836 699068
rect 414836 699012 414892 699068
rect 414892 699012 414896 699068
rect 414832 699008 414896 699012
rect 414912 699068 414976 699072
rect 414912 699012 414916 699068
rect 414916 699012 414972 699068
rect 414972 699012 414976 699068
rect 414912 699008 414976 699012
rect 414992 699068 415056 699072
rect 414992 699012 414996 699068
rect 414996 699012 415052 699068
rect 415052 699012 415056 699068
rect 414992 699008 415056 699012
rect 415072 699068 415136 699072
rect 415072 699012 415076 699068
rect 415076 699012 415132 699068
rect 415132 699012 415136 699068
rect 415072 699008 415136 699012
rect 415152 699068 415216 699072
rect 415152 699012 415156 699068
rect 415156 699012 415212 699068
rect 415212 699012 415216 699068
rect 415152 699008 415216 699012
rect 415232 699068 415296 699072
rect 415232 699012 415236 699068
rect 415236 699012 415292 699068
rect 415292 699012 415296 699068
rect 415232 699008 415296 699012
rect 415312 699068 415376 699072
rect 415312 699012 415316 699068
rect 415316 699012 415372 699068
rect 415372 699012 415376 699068
rect 415312 699008 415376 699012
rect 450832 699068 450896 699072
rect 450832 699012 450836 699068
rect 450836 699012 450892 699068
rect 450892 699012 450896 699068
rect 450832 699008 450896 699012
rect 450912 699068 450976 699072
rect 450912 699012 450916 699068
rect 450916 699012 450972 699068
rect 450972 699012 450976 699068
rect 450912 699008 450976 699012
rect 450992 699068 451056 699072
rect 450992 699012 450996 699068
rect 450996 699012 451052 699068
rect 451052 699012 451056 699068
rect 450992 699008 451056 699012
rect 451072 699068 451136 699072
rect 451072 699012 451076 699068
rect 451076 699012 451132 699068
rect 451132 699012 451136 699068
rect 451072 699008 451136 699012
rect 451152 699068 451216 699072
rect 451152 699012 451156 699068
rect 451156 699012 451212 699068
rect 451212 699012 451216 699068
rect 451152 699008 451216 699012
rect 451232 699068 451296 699072
rect 451232 699012 451236 699068
rect 451236 699012 451292 699068
rect 451292 699012 451296 699068
rect 451232 699008 451296 699012
rect 451312 699068 451376 699072
rect 451312 699012 451316 699068
rect 451316 699012 451372 699068
rect 451372 699012 451376 699068
rect 451312 699008 451376 699012
rect 486832 699068 486896 699072
rect 486832 699012 486836 699068
rect 486836 699012 486892 699068
rect 486892 699012 486896 699068
rect 486832 699008 486896 699012
rect 486912 699068 486976 699072
rect 486912 699012 486916 699068
rect 486916 699012 486972 699068
rect 486972 699012 486976 699068
rect 486912 699008 486976 699012
rect 486992 699068 487056 699072
rect 486992 699012 486996 699068
rect 486996 699012 487052 699068
rect 487052 699012 487056 699068
rect 486992 699008 487056 699012
rect 487072 699068 487136 699072
rect 487072 699012 487076 699068
rect 487076 699012 487132 699068
rect 487132 699012 487136 699068
rect 487072 699008 487136 699012
rect 487152 699068 487216 699072
rect 487152 699012 487156 699068
rect 487156 699012 487212 699068
rect 487212 699012 487216 699068
rect 487152 699008 487216 699012
rect 487232 699068 487296 699072
rect 487232 699012 487236 699068
rect 487236 699012 487292 699068
rect 487292 699012 487296 699068
rect 487232 699008 487296 699012
rect 487312 699068 487376 699072
rect 487312 699012 487316 699068
rect 487316 699012 487372 699068
rect 487372 699012 487376 699068
rect 487312 699008 487376 699012
rect 522832 699068 522896 699072
rect 522832 699012 522836 699068
rect 522836 699012 522892 699068
rect 522892 699012 522896 699068
rect 522832 699008 522896 699012
rect 522912 699068 522976 699072
rect 522912 699012 522916 699068
rect 522916 699012 522972 699068
rect 522972 699012 522976 699068
rect 522912 699008 522976 699012
rect 522992 699068 523056 699072
rect 522992 699012 522996 699068
rect 522996 699012 523052 699068
rect 523052 699012 523056 699068
rect 522992 699008 523056 699012
rect 523072 699068 523136 699072
rect 523072 699012 523076 699068
rect 523076 699012 523132 699068
rect 523132 699012 523136 699068
rect 523072 699008 523136 699012
rect 523152 699068 523216 699072
rect 523152 699012 523156 699068
rect 523156 699012 523212 699068
rect 523212 699012 523216 699068
rect 523152 699008 523216 699012
rect 523232 699068 523296 699072
rect 523232 699012 523236 699068
rect 523236 699012 523292 699068
rect 523292 699012 523296 699068
rect 523232 699008 523296 699012
rect 523312 699068 523376 699072
rect 523312 699012 523316 699068
rect 523316 699012 523372 699068
rect 523372 699012 523376 699068
rect 523312 699008 523376 699012
rect 558832 699068 558896 699072
rect 558832 699012 558836 699068
rect 558836 699012 558892 699068
rect 558892 699012 558896 699068
rect 558832 699008 558896 699012
rect 558912 699068 558976 699072
rect 558912 699012 558916 699068
rect 558916 699012 558972 699068
rect 558972 699012 558976 699068
rect 558912 699008 558976 699012
rect 558992 699068 559056 699072
rect 558992 699012 558996 699068
rect 558996 699012 559052 699068
rect 559052 699012 559056 699068
rect 558992 699008 559056 699012
rect 559072 699068 559136 699072
rect 559072 699012 559076 699068
rect 559076 699012 559132 699068
rect 559132 699012 559136 699068
rect 559072 699008 559136 699012
rect 559152 699068 559216 699072
rect 559152 699012 559156 699068
rect 559156 699012 559212 699068
rect 559212 699012 559216 699068
rect 559152 699008 559216 699012
rect 559232 699068 559296 699072
rect 559232 699012 559236 699068
rect 559236 699012 559292 699068
rect 559292 699012 559296 699068
rect 559232 699008 559296 699012
rect 559312 699068 559376 699072
rect 559312 699012 559316 699068
rect 559316 699012 559372 699068
rect 559372 699012 559376 699068
rect 559312 699008 559376 699012
rect 36832 698524 36896 698528
rect 36832 698468 36836 698524
rect 36836 698468 36892 698524
rect 36892 698468 36896 698524
rect 36832 698464 36896 698468
rect 36912 698524 36976 698528
rect 36912 698468 36916 698524
rect 36916 698468 36972 698524
rect 36972 698468 36976 698524
rect 36912 698464 36976 698468
rect 36992 698524 37056 698528
rect 36992 698468 36996 698524
rect 36996 698468 37052 698524
rect 37052 698468 37056 698524
rect 36992 698464 37056 698468
rect 37072 698524 37136 698528
rect 37072 698468 37076 698524
rect 37076 698468 37132 698524
rect 37132 698468 37136 698524
rect 37072 698464 37136 698468
rect 37152 698524 37216 698528
rect 37152 698468 37156 698524
rect 37156 698468 37212 698524
rect 37212 698468 37216 698524
rect 37152 698464 37216 698468
rect 37232 698524 37296 698528
rect 37232 698468 37236 698524
rect 37236 698468 37292 698524
rect 37292 698468 37296 698524
rect 37232 698464 37296 698468
rect 37312 698524 37376 698528
rect 37312 698468 37316 698524
rect 37316 698468 37372 698524
rect 37372 698468 37376 698524
rect 37312 698464 37376 698468
rect 72832 698524 72896 698528
rect 72832 698468 72836 698524
rect 72836 698468 72892 698524
rect 72892 698468 72896 698524
rect 72832 698464 72896 698468
rect 72912 698524 72976 698528
rect 72912 698468 72916 698524
rect 72916 698468 72972 698524
rect 72972 698468 72976 698524
rect 72912 698464 72976 698468
rect 72992 698524 73056 698528
rect 72992 698468 72996 698524
rect 72996 698468 73052 698524
rect 73052 698468 73056 698524
rect 72992 698464 73056 698468
rect 73072 698524 73136 698528
rect 73072 698468 73076 698524
rect 73076 698468 73132 698524
rect 73132 698468 73136 698524
rect 73072 698464 73136 698468
rect 73152 698524 73216 698528
rect 73152 698468 73156 698524
rect 73156 698468 73212 698524
rect 73212 698468 73216 698524
rect 73152 698464 73216 698468
rect 73232 698524 73296 698528
rect 73232 698468 73236 698524
rect 73236 698468 73292 698524
rect 73292 698468 73296 698524
rect 73232 698464 73296 698468
rect 73312 698524 73376 698528
rect 73312 698468 73316 698524
rect 73316 698468 73372 698524
rect 73372 698468 73376 698524
rect 73312 698464 73376 698468
rect 108832 698524 108896 698528
rect 108832 698468 108836 698524
rect 108836 698468 108892 698524
rect 108892 698468 108896 698524
rect 108832 698464 108896 698468
rect 108912 698524 108976 698528
rect 108912 698468 108916 698524
rect 108916 698468 108972 698524
rect 108972 698468 108976 698524
rect 108912 698464 108976 698468
rect 108992 698524 109056 698528
rect 108992 698468 108996 698524
rect 108996 698468 109052 698524
rect 109052 698468 109056 698524
rect 108992 698464 109056 698468
rect 109072 698524 109136 698528
rect 109072 698468 109076 698524
rect 109076 698468 109132 698524
rect 109132 698468 109136 698524
rect 109072 698464 109136 698468
rect 109152 698524 109216 698528
rect 109152 698468 109156 698524
rect 109156 698468 109212 698524
rect 109212 698468 109216 698524
rect 109152 698464 109216 698468
rect 109232 698524 109296 698528
rect 109232 698468 109236 698524
rect 109236 698468 109292 698524
rect 109292 698468 109296 698524
rect 109232 698464 109296 698468
rect 109312 698524 109376 698528
rect 109312 698468 109316 698524
rect 109316 698468 109372 698524
rect 109372 698468 109376 698524
rect 109312 698464 109376 698468
rect 144832 698524 144896 698528
rect 144832 698468 144836 698524
rect 144836 698468 144892 698524
rect 144892 698468 144896 698524
rect 144832 698464 144896 698468
rect 144912 698524 144976 698528
rect 144912 698468 144916 698524
rect 144916 698468 144972 698524
rect 144972 698468 144976 698524
rect 144912 698464 144976 698468
rect 144992 698524 145056 698528
rect 144992 698468 144996 698524
rect 144996 698468 145052 698524
rect 145052 698468 145056 698524
rect 144992 698464 145056 698468
rect 145072 698524 145136 698528
rect 145072 698468 145076 698524
rect 145076 698468 145132 698524
rect 145132 698468 145136 698524
rect 145072 698464 145136 698468
rect 145152 698524 145216 698528
rect 145152 698468 145156 698524
rect 145156 698468 145212 698524
rect 145212 698468 145216 698524
rect 145152 698464 145216 698468
rect 145232 698524 145296 698528
rect 145232 698468 145236 698524
rect 145236 698468 145292 698524
rect 145292 698468 145296 698524
rect 145232 698464 145296 698468
rect 145312 698524 145376 698528
rect 145312 698468 145316 698524
rect 145316 698468 145372 698524
rect 145372 698468 145376 698524
rect 145312 698464 145376 698468
rect 180832 698524 180896 698528
rect 180832 698468 180836 698524
rect 180836 698468 180892 698524
rect 180892 698468 180896 698524
rect 180832 698464 180896 698468
rect 180912 698524 180976 698528
rect 180912 698468 180916 698524
rect 180916 698468 180972 698524
rect 180972 698468 180976 698524
rect 180912 698464 180976 698468
rect 180992 698524 181056 698528
rect 180992 698468 180996 698524
rect 180996 698468 181052 698524
rect 181052 698468 181056 698524
rect 180992 698464 181056 698468
rect 181072 698524 181136 698528
rect 181072 698468 181076 698524
rect 181076 698468 181132 698524
rect 181132 698468 181136 698524
rect 181072 698464 181136 698468
rect 181152 698524 181216 698528
rect 181152 698468 181156 698524
rect 181156 698468 181212 698524
rect 181212 698468 181216 698524
rect 181152 698464 181216 698468
rect 181232 698524 181296 698528
rect 181232 698468 181236 698524
rect 181236 698468 181292 698524
rect 181292 698468 181296 698524
rect 181232 698464 181296 698468
rect 181312 698524 181376 698528
rect 181312 698468 181316 698524
rect 181316 698468 181372 698524
rect 181372 698468 181376 698524
rect 181312 698464 181376 698468
rect 216832 698524 216896 698528
rect 216832 698468 216836 698524
rect 216836 698468 216892 698524
rect 216892 698468 216896 698524
rect 216832 698464 216896 698468
rect 216912 698524 216976 698528
rect 216912 698468 216916 698524
rect 216916 698468 216972 698524
rect 216972 698468 216976 698524
rect 216912 698464 216976 698468
rect 216992 698524 217056 698528
rect 216992 698468 216996 698524
rect 216996 698468 217052 698524
rect 217052 698468 217056 698524
rect 216992 698464 217056 698468
rect 217072 698524 217136 698528
rect 217072 698468 217076 698524
rect 217076 698468 217132 698524
rect 217132 698468 217136 698524
rect 217072 698464 217136 698468
rect 217152 698524 217216 698528
rect 217152 698468 217156 698524
rect 217156 698468 217212 698524
rect 217212 698468 217216 698524
rect 217152 698464 217216 698468
rect 217232 698524 217296 698528
rect 217232 698468 217236 698524
rect 217236 698468 217292 698524
rect 217292 698468 217296 698524
rect 217232 698464 217296 698468
rect 217312 698524 217376 698528
rect 217312 698468 217316 698524
rect 217316 698468 217372 698524
rect 217372 698468 217376 698524
rect 217312 698464 217376 698468
rect 252832 698524 252896 698528
rect 252832 698468 252836 698524
rect 252836 698468 252892 698524
rect 252892 698468 252896 698524
rect 252832 698464 252896 698468
rect 252912 698524 252976 698528
rect 252912 698468 252916 698524
rect 252916 698468 252972 698524
rect 252972 698468 252976 698524
rect 252912 698464 252976 698468
rect 252992 698524 253056 698528
rect 252992 698468 252996 698524
rect 252996 698468 253052 698524
rect 253052 698468 253056 698524
rect 252992 698464 253056 698468
rect 253072 698524 253136 698528
rect 253072 698468 253076 698524
rect 253076 698468 253132 698524
rect 253132 698468 253136 698524
rect 253072 698464 253136 698468
rect 253152 698524 253216 698528
rect 253152 698468 253156 698524
rect 253156 698468 253212 698524
rect 253212 698468 253216 698524
rect 253152 698464 253216 698468
rect 253232 698524 253296 698528
rect 253232 698468 253236 698524
rect 253236 698468 253292 698524
rect 253292 698468 253296 698524
rect 253232 698464 253296 698468
rect 253312 698524 253376 698528
rect 253312 698468 253316 698524
rect 253316 698468 253372 698524
rect 253372 698468 253376 698524
rect 253312 698464 253376 698468
rect 288832 698524 288896 698528
rect 288832 698468 288836 698524
rect 288836 698468 288892 698524
rect 288892 698468 288896 698524
rect 288832 698464 288896 698468
rect 288912 698524 288976 698528
rect 288912 698468 288916 698524
rect 288916 698468 288972 698524
rect 288972 698468 288976 698524
rect 288912 698464 288976 698468
rect 288992 698524 289056 698528
rect 288992 698468 288996 698524
rect 288996 698468 289052 698524
rect 289052 698468 289056 698524
rect 288992 698464 289056 698468
rect 289072 698524 289136 698528
rect 289072 698468 289076 698524
rect 289076 698468 289132 698524
rect 289132 698468 289136 698524
rect 289072 698464 289136 698468
rect 289152 698524 289216 698528
rect 289152 698468 289156 698524
rect 289156 698468 289212 698524
rect 289212 698468 289216 698524
rect 289152 698464 289216 698468
rect 289232 698524 289296 698528
rect 289232 698468 289236 698524
rect 289236 698468 289292 698524
rect 289292 698468 289296 698524
rect 289232 698464 289296 698468
rect 289312 698524 289376 698528
rect 289312 698468 289316 698524
rect 289316 698468 289372 698524
rect 289372 698468 289376 698524
rect 289312 698464 289376 698468
rect 324832 698524 324896 698528
rect 324832 698468 324836 698524
rect 324836 698468 324892 698524
rect 324892 698468 324896 698524
rect 324832 698464 324896 698468
rect 324912 698524 324976 698528
rect 324912 698468 324916 698524
rect 324916 698468 324972 698524
rect 324972 698468 324976 698524
rect 324912 698464 324976 698468
rect 324992 698524 325056 698528
rect 324992 698468 324996 698524
rect 324996 698468 325052 698524
rect 325052 698468 325056 698524
rect 324992 698464 325056 698468
rect 325072 698524 325136 698528
rect 325072 698468 325076 698524
rect 325076 698468 325132 698524
rect 325132 698468 325136 698524
rect 325072 698464 325136 698468
rect 325152 698524 325216 698528
rect 325152 698468 325156 698524
rect 325156 698468 325212 698524
rect 325212 698468 325216 698524
rect 325152 698464 325216 698468
rect 325232 698524 325296 698528
rect 325232 698468 325236 698524
rect 325236 698468 325292 698524
rect 325292 698468 325296 698524
rect 325232 698464 325296 698468
rect 325312 698524 325376 698528
rect 325312 698468 325316 698524
rect 325316 698468 325372 698524
rect 325372 698468 325376 698524
rect 325312 698464 325376 698468
rect 360832 698524 360896 698528
rect 360832 698468 360836 698524
rect 360836 698468 360892 698524
rect 360892 698468 360896 698524
rect 360832 698464 360896 698468
rect 360912 698524 360976 698528
rect 360912 698468 360916 698524
rect 360916 698468 360972 698524
rect 360972 698468 360976 698524
rect 360912 698464 360976 698468
rect 360992 698524 361056 698528
rect 360992 698468 360996 698524
rect 360996 698468 361052 698524
rect 361052 698468 361056 698524
rect 360992 698464 361056 698468
rect 361072 698524 361136 698528
rect 361072 698468 361076 698524
rect 361076 698468 361132 698524
rect 361132 698468 361136 698524
rect 361072 698464 361136 698468
rect 361152 698524 361216 698528
rect 361152 698468 361156 698524
rect 361156 698468 361212 698524
rect 361212 698468 361216 698524
rect 361152 698464 361216 698468
rect 361232 698524 361296 698528
rect 361232 698468 361236 698524
rect 361236 698468 361292 698524
rect 361292 698468 361296 698524
rect 361232 698464 361296 698468
rect 361312 698524 361376 698528
rect 361312 698468 361316 698524
rect 361316 698468 361372 698524
rect 361372 698468 361376 698524
rect 361312 698464 361376 698468
rect 396832 698524 396896 698528
rect 396832 698468 396836 698524
rect 396836 698468 396892 698524
rect 396892 698468 396896 698524
rect 396832 698464 396896 698468
rect 396912 698524 396976 698528
rect 396912 698468 396916 698524
rect 396916 698468 396972 698524
rect 396972 698468 396976 698524
rect 396912 698464 396976 698468
rect 396992 698524 397056 698528
rect 396992 698468 396996 698524
rect 396996 698468 397052 698524
rect 397052 698468 397056 698524
rect 396992 698464 397056 698468
rect 397072 698524 397136 698528
rect 397072 698468 397076 698524
rect 397076 698468 397132 698524
rect 397132 698468 397136 698524
rect 397072 698464 397136 698468
rect 397152 698524 397216 698528
rect 397152 698468 397156 698524
rect 397156 698468 397212 698524
rect 397212 698468 397216 698524
rect 397152 698464 397216 698468
rect 397232 698524 397296 698528
rect 397232 698468 397236 698524
rect 397236 698468 397292 698524
rect 397292 698468 397296 698524
rect 397232 698464 397296 698468
rect 397312 698524 397376 698528
rect 397312 698468 397316 698524
rect 397316 698468 397372 698524
rect 397372 698468 397376 698524
rect 397312 698464 397376 698468
rect 432832 698524 432896 698528
rect 432832 698468 432836 698524
rect 432836 698468 432892 698524
rect 432892 698468 432896 698524
rect 432832 698464 432896 698468
rect 432912 698524 432976 698528
rect 432912 698468 432916 698524
rect 432916 698468 432972 698524
rect 432972 698468 432976 698524
rect 432912 698464 432976 698468
rect 432992 698524 433056 698528
rect 432992 698468 432996 698524
rect 432996 698468 433052 698524
rect 433052 698468 433056 698524
rect 432992 698464 433056 698468
rect 433072 698524 433136 698528
rect 433072 698468 433076 698524
rect 433076 698468 433132 698524
rect 433132 698468 433136 698524
rect 433072 698464 433136 698468
rect 433152 698524 433216 698528
rect 433152 698468 433156 698524
rect 433156 698468 433212 698524
rect 433212 698468 433216 698524
rect 433152 698464 433216 698468
rect 433232 698524 433296 698528
rect 433232 698468 433236 698524
rect 433236 698468 433292 698524
rect 433292 698468 433296 698524
rect 433232 698464 433296 698468
rect 433312 698524 433376 698528
rect 433312 698468 433316 698524
rect 433316 698468 433372 698524
rect 433372 698468 433376 698524
rect 433312 698464 433376 698468
rect 468832 698524 468896 698528
rect 468832 698468 468836 698524
rect 468836 698468 468892 698524
rect 468892 698468 468896 698524
rect 468832 698464 468896 698468
rect 468912 698524 468976 698528
rect 468912 698468 468916 698524
rect 468916 698468 468972 698524
rect 468972 698468 468976 698524
rect 468912 698464 468976 698468
rect 468992 698524 469056 698528
rect 468992 698468 468996 698524
rect 468996 698468 469052 698524
rect 469052 698468 469056 698524
rect 468992 698464 469056 698468
rect 469072 698524 469136 698528
rect 469072 698468 469076 698524
rect 469076 698468 469132 698524
rect 469132 698468 469136 698524
rect 469072 698464 469136 698468
rect 469152 698524 469216 698528
rect 469152 698468 469156 698524
rect 469156 698468 469212 698524
rect 469212 698468 469216 698524
rect 469152 698464 469216 698468
rect 469232 698524 469296 698528
rect 469232 698468 469236 698524
rect 469236 698468 469292 698524
rect 469292 698468 469296 698524
rect 469232 698464 469296 698468
rect 469312 698524 469376 698528
rect 469312 698468 469316 698524
rect 469316 698468 469372 698524
rect 469372 698468 469376 698524
rect 469312 698464 469376 698468
rect 504832 698524 504896 698528
rect 504832 698468 504836 698524
rect 504836 698468 504892 698524
rect 504892 698468 504896 698524
rect 504832 698464 504896 698468
rect 504912 698524 504976 698528
rect 504912 698468 504916 698524
rect 504916 698468 504972 698524
rect 504972 698468 504976 698524
rect 504912 698464 504976 698468
rect 504992 698524 505056 698528
rect 504992 698468 504996 698524
rect 504996 698468 505052 698524
rect 505052 698468 505056 698524
rect 504992 698464 505056 698468
rect 505072 698524 505136 698528
rect 505072 698468 505076 698524
rect 505076 698468 505132 698524
rect 505132 698468 505136 698524
rect 505072 698464 505136 698468
rect 505152 698524 505216 698528
rect 505152 698468 505156 698524
rect 505156 698468 505212 698524
rect 505212 698468 505216 698524
rect 505152 698464 505216 698468
rect 505232 698524 505296 698528
rect 505232 698468 505236 698524
rect 505236 698468 505292 698524
rect 505292 698468 505296 698524
rect 505232 698464 505296 698468
rect 505312 698524 505376 698528
rect 505312 698468 505316 698524
rect 505316 698468 505372 698524
rect 505372 698468 505376 698524
rect 505312 698464 505376 698468
rect 540832 698524 540896 698528
rect 540832 698468 540836 698524
rect 540836 698468 540892 698524
rect 540892 698468 540896 698524
rect 540832 698464 540896 698468
rect 540912 698524 540976 698528
rect 540912 698468 540916 698524
rect 540916 698468 540972 698524
rect 540972 698468 540976 698524
rect 540912 698464 540976 698468
rect 540992 698524 541056 698528
rect 540992 698468 540996 698524
rect 540996 698468 541052 698524
rect 541052 698468 541056 698524
rect 540992 698464 541056 698468
rect 541072 698524 541136 698528
rect 541072 698468 541076 698524
rect 541076 698468 541132 698524
rect 541132 698468 541136 698524
rect 541072 698464 541136 698468
rect 541152 698524 541216 698528
rect 541152 698468 541156 698524
rect 541156 698468 541212 698524
rect 541212 698468 541216 698524
rect 541152 698464 541216 698468
rect 541232 698524 541296 698528
rect 541232 698468 541236 698524
rect 541236 698468 541292 698524
rect 541292 698468 541296 698524
rect 541232 698464 541296 698468
rect 541312 698524 541376 698528
rect 541312 698468 541316 698524
rect 541316 698468 541372 698524
rect 541372 698468 541376 698524
rect 541312 698464 541376 698468
rect 576832 698524 576896 698528
rect 576832 698468 576836 698524
rect 576836 698468 576892 698524
rect 576892 698468 576896 698524
rect 576832 698464 576896 698468
rect 576912 698524 576976 698528
rect 576912 698468 576916 698524
rect 576916 698468 576972 698524
rect 576972 698468 576976 698524
rect 576912 698464 576976 698468
rect 576992 698524 577056 698528
rect 576992 698468 576996 698524
rect 576996 698468 577052 698524
rect 577052 698468 577056 698524
rect 576992 698464 577056 698468
rect 577072 698524 577136 698528
rect 577072 698468 577076 698524
rect 577076 698468 577132 698524
rect 577132 698468 577136 698524
rect 577072 698464 577136 698468
rect 577152 698524 577216 698528
rect 577152 698468 577156 698524
rect 577156 698468 577212 698524
rect 577212 698468 577216 698524
rect 577152 698464 577216 698468
rect 577232 698524 577296 698528
rect 577232 698468 577236 698524
rect 577236 698468 577292 698524
rect 577292 698468 577296 698524
rect 577232 698464 577296 698468
rect 577312 698524 577376 698528
rect 577312 698468 577316 698524
rect 577316 698468 577372 698524
rect 577372 698468 577376 698524
rect 577312 698464 577376 698468
rect 241468 695948 241532 696012
rect 260788 695948 260852 696012
rect 318748 695948 318812 696012
rect 144868 695812 144932 695876
rect 144868 695540 144932 695604
rect 176516 695540 176580 695604
rect 241468 695676 241532 695740
rect 260788 695676 260852 695740
rect 318748 695676 318812 695740
rect 347636 695812 347700 695876
rect 367140 695812 367204 695876
rect 434668 695812 434732 695876
rect 473308 695948 473372 696012
rect 442948 695812 443012 695876
rect 463740 695812 463804 695876
rect 367140 695676 367204 695740
rect 412588 695676 412652 695740
rect 463740 695676 463804 695740
rect 347636 695540 347700 695604
rect 426388 695540 426452 695604
rect 434668 695540 434732 695604
rect 473308 695540 473372 695604
rect 442948 695404 443012 695468
rect 17172 695268 17236 695332
rect 157012 695328 157076 695332
rect 157012 695272 157062 695328
rect 157062 695272 157076 695328
rect 157012 695268 157076 695272
rect 412588 695268 412652 695332
rect 521332 695328 521396 695332
rect 521332 695272 521382 695328
rect 521382 695272 521396 695328
rect 521332 695268 521396 695272
rect 176516 694860 176580 694924
rect 178908 694860 178972 694924
rect 311572 694860 311636 694924
rect 124260 694724 124324 694788
rect 133644 694724 133708 694788
rect 153332 694724 153396 694788
rect 111012 694452 111076 694516
rect 115612 694452 115676 694516
rect 273300 694724 273364 694788
rect 279924 694724 279988 694788
rect 299796 694724 299860 694788
rect 311204 694724 311268 694788
rect 321508 694860 321572 694924
rect 323716 694860 323780 694924
rect 489684 694860 489748 694924
rect 318748 694724 318812 694788
rect 186268 694588 186332 694652
rect 256004 694588 256068 694652
rect 275324 694588 275388 694652
rect 284892 694588 284956 694652
rect 17172 694180 17236 694244
rect 133644 694316 133708 694380
rect 153148 694316 153212 694380
rect 160876 694316 160940 694380
rect 164188 694316 164252 694380
rect 185900 694316 185964 694380
rect 196020 694452 196084 694516
rect 124260 694180 124324 694244
rect 178908 694180 178972 694244
rect 9628 694044 9692 694108
rect 9812 693908 9876 693972
rect 31524 694044 31588 694108
rect 89852 694044 89916 694108
rect 96660 694044 96724 694108
rect 140820 694044 140884 694108
rect 143580 694044 143644 694108
rect 152964 694044 153028 694108
rect 160876 694044 160940 694108
rect 164188 694044 164252 694108
rect 185900 694044 185964 694108
rect 186268 694044 186332 694108
rect 195836 694316 195900 694380
rect 215340 694452 215404 694516
rect 215156 694316 215220 694380
rect 263548 694452 263612 694516
rect 273668 694452 273732 694516
rect 283052 694452 283116 694516
rect 311756 694588 311820 694652
rect 318932 694588 318996 694652
rect 331076 694724 331140 694788
rect 331260 694588 331324 694652
rect 253796 694316 253860 694380
rect 254348 694316 254412 694380
rect 256004 694180 256068 694244
rect 280062 694316 280126 694380
rect 282684 694316 282748 694380
rect 283236 694316 283300 694380
rect 195836 694044 195900 694108
rect 196020 694044 196084 694108
rect 205404 694044 205468 694108
rect 205956 694044 206020 694108
rect 215156 694044 215220 694108
rect 215340 694044 215404 694108
rect 224724 694044 224788 694108
rect 225276 694044 225340 694108
rect 244044 694044 244108 694108
rect 244596 694044 244660 694108
rect 263548 694044 263612 694108
rect 273300 694180 273364 694244
rect 275324 694180 275388 694244
rect 311572 694316 311636 694380
rect 311756 694316 311820 694380
rect 323532 694452 323596 694516
rect 323716 694452 323780 694516
rect 330708 694452 330772 694516
rect 340828 694588 340892 694652
rect 371924 694588 371988 694652
rect 379100 694588 379164 694652
rect 391244 694588 391308 694652
rect 398420 694588 398484 694652
rect 424916 694724 424980 694788
rect 425100 694724 425164 694788
rect 434300 694724 434364 694788
rect 461164 694724 461228 694788
rect 470364 694724 470428 694788
rect 470548 694588 470612 694652
rect 359964 694452 360028 694516
rect 369900 694452 369964 694516
rect 273668 694044 273732 694108
rect 282868 694044 282932 694108
rect 284892 694044 284956 694108
rect 299244 694044 299308 694108
rect 311204 694044 311268 694108
rect 321508 694044 321572 694108
rect 323532 694044 323596 694108
rect 330708 694044 330772 694108
rect 340828 694044 340892 694108
rect 360332 694316 360396 694380
rect 369716 694316 369780 694380
rect 390140 694452 390204 694516
rect 389220 694316 389284 694380
rect 420132 694452 420196 694516
rect 426388 694452 426452 694516
rect 371924 694180 371988 694244
rect 379100 694180 379164 694244
rect 391244 694180 391308 694244
rect 398420 694180 398484 694244
rect 420316 694180 420380 694244
rect 424732 694180 424796 694244
rect 424916 694180 424980 694244
rect 470364 694316 470428 694380
rect 470548 694316 470612 694380
rect 531268 694724 531332 694788
rect 511948 694588 512012 694652
rect 521516 694588 521580 694652
rect 489500 694316 489564 694380
rect 460980 694180 461044 694244
rect 500908 694452 500972 694516
rect 500908 694180 500972 694244
rect 521700 694452 521764 694516
rect 531268 694452 531332 694516
rect 550588 694452 550652 694516
rect 521700 694180 521764 694244
rect 550588 694180 550652 694244
rect 359964 694044 360028 694108
rect 360332 694044 360396 694108
rect 369716 694044 369780 694108
rect 369900 694044 369964 694108
rect 420132 694044 420196 694108
rect 425100 694044 425164 694108
rect 434484 694044 434548 694108
rect 434668 694044 434732 694108
rect 435036 694044 435100 694108
rect 511948 694044 512012 694108
rect 521516 694044 521580 694108
rect 521700 694044 521764 694108
rect 524460 694044 524524 694108
rect 539548 694044 539612 694108
rect 31892 693908 31956 693972
rect 37228 693908 37292 693972
rect 46796 693908 46860 693972
rect 56548 693908 56612 693972
rect 66116 693908 66180 693972
rect 75868 693908 75932 693972
rect 85436 693908 85500 693972
rect 89484 693908 89548 693972
rect 96844 693908 96908 693972
rect 111012 693908 111076 693972
rect 115612 693908 115676 693972
rect 124260 693908 124324 693972
rect 133644 693908 133708 693972
rect 140636 693908 140700 693972
rect 157012 693908 157076 693972
rect 173940 693908 174004 693972
rect 174124 693908 174188 693972
rect 420316 693908 420380 693972
rect 424916 693908 424980 693972
rect 434668 693908 434732 693972
rect 435036 693908 435100 693972
rect 543596 693908 543660 693972
rect 543780 693908 543844 693972
rect 562916 693908 562980 693972
rect 563100 693908 563164 693972
rect 55628 693772 55692 693836
rect 56364 693772 56428 693836
rect 74948 693772 75012 693836
rect 75684 693772 75748 693836
rect 108804 693772 108868 693836
rect 114140 693772 114204 693836
rect 162900 693772 162964 693836
rect 163820 693772 163884 693836
rect 424180 693772 424244 693836
rect 424916 693772 424980 693836
rect 434116 693772 434180 693836
rect 434484 693772 434548 693836
rect 434668 693772 434732 693836
rect 435220 693772 435284 693836
rect 503484 693772 503548 693836
rect 521700 693772 521764 693836
rect 524460 693772 524524 693836
rect 549116 693772 549180 693836
rect 123708 693636 123772 693700
rect 124076 693636 124140 693700
rect 163084 693636 163148 693700
rect 163636 693636 163700 693700
rect 423996 693636 424060 693700
rect 424732 693636 424796 693700
rect 433932 693636 433996 693700
rect 434484 693636 434548 693700
rect 473492 693636 473556 693700
rect 474044 693636 474108 693700
rect 521332 693636 521396 693700
rect 550588 693636 550652 693700
rect 550772 693636 550836 693700
rect 558868 693636 558932 693700
rect 565676 693364 565740 693428
rect 18832 6012 18896 6016
rect 18832 5956 18836 6012
rect 18836 5956 18892 6012
rect 18892 5956 18896 6012
rect 18832 5952 18896 5956
rect 18912 6012 18976 6016
rect 18912 5956 18916 6012
rect 18916 5956 18972 6012
rect 18972 5956 18976 6012
rect 18912 5952 18976 5956
rect 18992 6012 19056 6016
rect 18992 5956 18996 6012
rect 18996 5956 19052 6012
rect 19052 5956 19056 6012
rect 18992 5952 19056 5956
rect 19072 6012 19136 6016
rect 19072 5956 19076 6012
rect 19076 5956 19132 6012
rect 19132 5956 19136 6012
rect 19072 5952 19136 5956
rect 19152 6012 19216 6016
rect 19152 5956 19156 6012
rect 19156 5956 19212 6012
rect 19212 5956 19216 6012
rect 19152 5952 19216 5956
rect 19232 6012 19296 6016
rect 19232 5956 19236 6012
rect 19236 5956 19292 6012
rect 19292 5956 19296 6012
rect 19232 5952 19296 5956
rect 19312 6012 19376 6016
rect 19312 5956 19316 6012
rect 19316 5956 19372 6012
rect 19372 5956 19376 6012
rect 19312 5952 19376 5956
rect 54832 6012 54896 6016
rect 54832 5956 54836 6012
rect 54836 5956 54892 6012
rect 54892 5956 54896 6012
rect 54832 5952 54896 5956
rect 54912 6012 54976 6016
rect 54912 5956 54916 6012
rect 54916 5956 54972 6012
rect 54972 5956 54976 6012
rect 54912 5952 54976 5956
rect 54992 6012 55056 6016
rect 54992 5956 54996 6012
rect 54996 5956 55052 6012
rect 55052 5956 55056 6012
rect 54992 5952 55056 5956
rect 55072 6012 55136 6016
rect 55072 5956 55076 6012
rect 55076 5956 55132 6012
rect 55132 5956 55136 6012
rect 55072 5952 55136 5956
rect 55152 6012 55216 6016
rect 55152 5956 55156 6012
rect 55156 5956 55212 6012
rect 55212 5956 55216 6012
rect 55152 5952 55216 5956
rect 55232 6012 55296 6016
rect 55232 5956 55236 6012
rect 55236 5956 55292 6012
rect 55292 5956 55296 6012
rect 55232 5952 55296 5956
rect 55312 6012 55376 6016
rect 55312 5956 55316 6012
rect 55316 5956 55372 6012
rect 55372 5956 55376 6012
rect 55312 5952 55376 5956
rect 90832 6012 90896 6016
rect 90832 5956 90836 6012
rect 90836 5956 90892 6012
rect 90892 5956 90896 6012
rect 90832 5952 90896 5956
rect 90912 6012 90976 6016
rect 90912 5956 90916 6012
rect 90916 5956 90972 6012
rect 90972 5956 90976 6012
rect 90912 5952 90976 5956
rect 90992 6012 91056 6016
rect 90992 5956 90996 6012
rect 90996 5956 91052 6012
rect 91052 5956 91056 6012
rect 90992 5952 91056 5956
rect 91072 6012 91136 6016
rect 91072 5956 91076 6012
rect 91076 5956 91132 6012
rect 91132 5956 91136 6012
rect 91072 5952 91136 5956
rect 91152 6012 91216 6016
rect 91152 5956 91156 6012
rect 91156 5956 91212 6012
rect 91212 5956 91216 6012
rect 91152 5952 91216 5956
rect 91232 6012 91296 6016
rect 91232 5956 91236 6012
rect 91236 5956 91292 6012
rect 91292 5956 91296 6012
rect 91232 5952 91296 5956
rect 91312 6012 91376 6016
rect 91312 5956 91316 6012
rect 91316 5956 91372 6012
rect 91372 5956 91376 6012
rect 91312 5952 91376 5956
rect 126832 6012 126896 6016
rect 126832 5956 126836 6012
rect 126836 5956 126892 6012
rect 126892 5956 126896 6012
rect 126832 5952 126896 5956
rect 126912 6012 126976 6016
rect 126912 5956 126916 6012
rect 126916 5956 126972 6012
rect 126972 5956 126976 6012
rect 126912 5952 126976 5956
rect 126992 6012 127056 6016
rect 126992 5956 126996 6012
rect 126996 5956 127052 6012
rect 127052 5956 127056 6012
rect 126992 5952 127056 5956
rect 127072 6012 127136 6016
rect 127072 5956 127076 6012
rect 127076 5956 127132 6012
rect 127132 5956 127136 6012
rect 127072 5952 127136 5956
rect 127152 6012 127216 6016
rect 127152 5956 127156 6012
rect 127156 5956 127212 6012
rect 127212 5956 127216 6012
rect 127152 5952 127216 5956
rect 127232 6012 127296 6016
rect 127232 5956 127236 6012
rect 127236 5956 127292 6012
rect 127292 5956 127296 6012
rect 127232 5952 127296 5956
rect 127312 6012 127376 6016
rect 127312 5956 127316 6012
rect 127316 5956 127372 6012
rect 127372 5956 127376 6012
rect 127312 5952 127376 5956
rect 162832 6012 162896 6016
rect 162832 5956 162836 6012
rect 162836 5956 162892 6012
rect 162892 5956 162896 6012
rect 162832 5952 162896 5956
rect 162912 6012 162976 6016
rect 162912 5956 162916 6012
rect 162916 5956 162972 6012
rect 162972 5956 162976 6012
rect 162912 5952 162976 5956
rect 162992 6012 163056 6016
rect 162992 5956 162996 6012
rect 162996 5956 163052 6012
rect 163052 5956 163056 6012
rect 162992 5952 163056 5956
rect 163072 6012 163136 6016
rect 163072 5956 163076 6012
rect 163076 5956 163132 6012
rect 163132 5956 163136 6012
rect 163072 5952 163136 5956
rect 163152 6012 163216 6016
rect 163152 5956 163156 6012
rect 163156 5956 163212 6012
rect 163212 5956 163216 6012
rect 163152 5952 163216 5956
rect 163232 6012 163296 6016
rect 163232 5956 163236 6012
rect 163236 5956 163292 6012
rect 163292 5956 163296 6012
rect 163232 5952 163296 5956
rect 163312 6012 163376 6016
rect 163312 5956 163316 6012
rect 163316 5956 163372 6012
rect 163372 5956 163376 6012
rect 163312 5952 163376 5956
rect 198832 6012 198896 6016
rect 198832 5956 198836 6012
rect 198836 5956 198892 6012
rect 198892 5956 198896 6012
rect 198832 5952 198896 5956
rect 198912 6012 198976 6016
rect 198912 5956 198916 6012
rect 198916 5956 198972 6012
rect 198972 5956 198976 6012
rect 198912 5952 198976 5956
rect 198992 6012 199056 6016
rect 198992 5956 198996 6012
rect 198996 5956 199052 6012
rect 199052 5956 199056 6012
rect 198992 5952 199056 5956
rect 199072 6012 199136 6016
rect 199072 5956 199076 6012
rect 199076 5956 199132 6012
rect 199132 5956 199136 6012
rect 199072 5952 199136 5956
rect 199152 6012 199216 6016
rect 199152 5956 199156 6012
rect 199156 5956 199212 6012
rect 199212 5956 199216 6012
rect 199152 5952 199216 5956
rect 199232 6012 199296 6016
rect 199232 5956 199236 6012
rect 199236 5956 199292 6012
rect 199292 5956 199296 6012
rect 199232 5952 199296 5956
rect 199312 6012 199376 6016
rect 199312 5956 199316 6012
rect 199316 5956 199372 6012
rect 199372 5956 199376 6012
rect 199312 5952 199376 5956
rect 234832 6012 234896 6016
rect 234832 5956 234836 6012
rect 234836 5956 234892 6012
rect 234892 5956 234896 6012
rect 234832 5952 234896 5956
rect 234912 6012 234976 6016
rect 234912 5956 234916 6012
rect 234916 5956 234972 6012
rect 234972 5956 234976 6012
rect 234912 5952 234976 5956
rect 234992 6012 235056 6016
rect 234992 5956 234996 6012
rect 234996 5956 235052 6012
rect 235052 5956 235056 6012
rect 234992 5952 235056 5956
rect 235072 6012 235136 6016
rect 235072 5956 235076 6012
rect 235076 5956 235132 6012
rect 235132 5956 235136 6012
rect 235072 5952 235136 5956
rect 235152 6012 235216 6016
rect 235152 5956 235156 6012
rect 235156 5956 235212 6012
rect 235212 5956 235216 6012
rect 235152 5952 235216 5956
rect 235232 6012 235296 6016
rect 235232 5956 235236 6012
rect 235236 5956 235292 6012
rect 235292 5956 235296 6012
rect 235232 5952 235296 5956
rect 235312 6012 235376 6016
rect 235312 5956 235316 6012
rect 235316 5956 235372 6012
rect 235372 5956 235376 6012
rect 235312 5952 235376 5956
rect 270832 6012 270896 6016
rect 270832 5956 270836 6012
rect 270836 5956 270892 6012
rect 270892 5956 270896 6012
rect 270832 5952 270896 5956
rect 270912 6012 270976 6016
rect 270912 5956 270916 6012
rect 270916 5956 270972 6012
rect 270972 5956 270976 6012
rect 270912 5952 270976 5956
rect 270992 6012 271056 6016
rect 270992 5956 270996 6012
rect 270996 5956 271052 6012
rect 271052 5956 271056 6012
rect 270992 5952 271056 5956
rect 271072 6012 271136 6016
rect 271072 5956 271076 6012
rect 271076 5956 271132 6012
rect 271132 5956 271136 6012
rect 271072 5952 271136 5956
rect 271152 6012 271216 6016
rect 271152 5956 271156 6012
rect 271156 5956 271212 6012
rect 271212 5956 271216 6012
rect 271152 5952 271216 5956
rect 271232 6012 271296 6016
rect 271232 5956 271236 6012
rect 271236 5956 271292 6012
rect 271292 5956 271296 6012
rect 271232 5952 271296 5956
rect 271312 6012 271376 6016
rect 271312 5956 271316 6012
rect 271316 5956 271372 6012
rect 271372 5956 271376 6012
rect 271312 5952 271376 5956
rect 306832 6012 306896 6016
rect 306832 5956 306836 6012
rect 306836 5956 306892 6012
rect 306892 5956 306896 6012
rect 306832 5952 306896 5956
rect 306912 6012 306976 6016
rect 306912 5956 306916 6012
rect 306916 5956 306972 6012
rect 306972 5956 306976 6012
rect 306912 5952 306976 5956
rect 306992 6012 307056 6016
rect 306992 5956 306996 6012
rect 306996 5956 307052 6012
rect 307052 5956 307056 6012
rect 306992 5952 307056 5956
rect 307072 6012 307136 6016
rect 307072 5956 307076 6012
rect 307076 5956 307132 6012
rect 307132 5956 307136 6012
rect 307072 5952 307136 5956
rect 307152 6012 307216 6016
rect 307152 5956 307156 6012
rect 307156 5956 307212 6012
rect 307212 5956 307216 6012
rect 307152 5952 307216 5956
rect 307232 6012 307296 6016
rect 307232 5956 307236 6012
rect 307236 5956 307292 6012
rect 307292 5956 307296 6012
rect 307232 5952 307296 5956
rect 307312 6012 307376 6016
rect 307312 5956 307316 6012
rect 307316 5956 307372 6012
rect 307372 5956 307376 6012
rect 307312 5952 307376 5956
rect 342832 6012 342896 6016
rect 342832 5956 342836 6012
rect 342836 5956 342892 6012
rect 342892 5956 342896 6012
rect 342832 5952 342896 5956
rect 342912 6012 342976 6016
rect 342912 5956 342916 6012
rect 342916 5956 342972 6012
rect 342972 5956 342976 6012
rect 342912 5952 342976 5956
rect 342992 6012 343056 6016
rect 342992 5956 342996 6012
rect 342996 5956 343052 6012
rect 343052 5956 343056 6012
rect 342992 5952 343056 5956
rect 343072 6012 343136 6016
rect 343072 5956 343076 6012
rect 343076 5956 343132 6012
rect 343132 5956 343136 6012
rect 343072 5952 343136 5956
rect 343152 6012 343216 6016
rect 343152 5956 343156 6012
rect 343156 5956 343212 6012
rect 343212 5956 343216 6012
rect 343152 5952 343216 5956
rect 343232 6012 343296 6016
rect 343232 5956 343236 6012
rect 343236 5956 343292 6012
rect 343292 5956 343296 6012
rect 343232 5952 343296 5956
rect 343312 6012 343376 6016
rect 343312 5956 343316 6012
rect 343316 5956 343372 6012
rect 343372 5956 343376 6012
rect 343312 5952 343376 5956
rect 378832 6012 378896 6016
rect 378832 5956 378836 6012
rect 378836 5956 378892 6012
rect 378892 5956 378896 6012
rect 378832 5952 378896 5956
rect 378912 6012 378976 6016
rect 378912 5956 378916 6012
rect 378916 5956 378972 6012
rect 378972 5956 378976 6012
rect 378912 5952 378976 5956
rect 378992 6012 379056 6016
rect 378992 5956 378996 6012
rect 378996 5956 379052 6012
rect 379052 5956 379056 6012
rect 378992 5952 379056 5956
rect 379072 6012 379136 6016
rect 379072 5956 379076 6012
rect 379076 5956 379132 6012
rect 379132 5956 379136 6012
rect 379072 5952 379136 5956
rect 379152 6012 379216 6016
rect 379152 5956 379156 6012
rect 379156 5956 379212 6012
rect 379212 5956 379216 6012
rect 379152 5952 379216 5956
rect 379232 6012 379296 6016
rect 379232 5956 379236 6012
rect 379236 5956 379292 6012
rect 379292 5956 379296 6012
rect 379232 5952 379296 5956
rect 379312 6012 379376 6016
rect 379312 5956 379316 6012
rect 379316 5956 379372 6012
rect 379372 5956 379376 6012
rect 379312 5952 379376 5956
rect 414832 6012 414896 6016
rect 414832 5956 414836 6012
rect 414836 5956 414892 6012
rect 414892 5956 414896 6012
rect 414832 5952 414896 5956
rect 414912 6012 414976 6016
rect 414912 5956 414916 6012
rect 414916 5956 414972 6012
rect 414972 5956 414976 6012
rect 414912 5952 414976 5956
rect 414992 6012 415056 6016
rect 414992 5956 414996 6012
rect 414996 5956 415052 6012
rect 415052 5956 415056 6012
rect 414992 5952 415056 5956
rect 415072 6012 415136 6016
rect 415072 5956 415076 6012
rect 415076 5956 415132 6012
rect 415132 5956 415136 6012
rect 415072 5952 415136 5956
rect 415152 6012 415216 6016
rect 415152 5956 415156 6012
rect 415156 5956 415212 6012
rect 415212 5956 415216 6012
rect 415152 5952 415216 5956
rect 415232 6012 415296 6016
rect 415232 5956 415236 6012
rect 415236 5956 415292 6012
rect 415292 5956 415296 6012
rect 415232 5952 415296 5956
rect 415312 6012 415376 6016
rect 415312 5956 415316 6012
rect 415316 5956 415372 6012
rect 415372 5956 415376 6012
rect 415312 5952 415376 5956
rect 450832 6012 450896 6016
rect 450832 5956 450836 6012
rect 450836 5956 450892 6012
rect 450892 5956 450896 6012
rect 450832 5952 450896 5956
rect 450912 6012 450976 6016
rect 450912 5956 450916 6012
rect 450916 5956 450972 6012
rect 450972 5956 450976 6012
rect 450912 5952 450976 5956
rect 450992 6012 451056 6016
rect 450992 5956 450996 6012
rect 450996 5956 451052 6012
rect 451052 5956 451056 6012
rect 450992 5952 451056 5956
rect 451072 6012 451136 6016
rect 451072 5956 451076 6012
rect 451076 5956 451132 6012
rect 451132 5956 451136 6012
rect 451072 5952 451136 5956
rect 451152 6012 451216 6016
rect 451152 5956 451156 6012
rect 451156 5956 451212 6012
rect 451212 5956 451216 6012
rect 451152 5952 451216 5956
rect 451232 6012 451296 6016
rect 451232 5956 451236 6012
rect 451236 5956 451292 6012
rect 451292 5956 451296 6012
rect 451232 5952 451296 5956
rect 451312 6012 451376 6016
rect 451312 5956 451316 6012
rect 451316 5956 451372 6012
rect 451372 5956 451376 6012
rect 451312 5952 451376 5956
rect 486832 6012 486896 6016
rect 486832 5956 486836 6012
rect 486836 5956 486892 6012
rect 486892 5956 486896 6012
rect 486832 5952 486896 5956
rect 486912 6012 486976 6016
rect 486912 5956 486916 6012
rect 486916 5956 486972 6012
rect 486972 5956 486976 6012
rect 486912 5952 486976 5956
rect 486992 6012 487056 6016
rect 486992 5956 486996 6012
rect 486996 5956 487052 6012
rect 487052 5956 487056 6012
rect 486992 5952 487056 5956
rect 487072 6012 487136 6016
rect 487072 5956 487076 6012
rect 487076 5956 487132 6012
rect 487132 5956 487136 6012
rect 487072 5952 487136 5956
rect 487152 6012 487216 6016
rect 487152 5956 487156 6012
rect 487156 5956 487212 6012
rect 487212 5956 487216 6012
rect 487152 5952 487216 5956
rect 487232 6012 487296 6016
rect 487232 5956 487236 6012
rect 487236 5956 487292 6012
rect 487292 5956 487296 6012
rect 487232 5952 487296 5956
rect 487312 6012 487376 6016
rect 487312 5956 487316 6012
rect 487316 5956 487372 6012
rect 487372 5956 487376 6012
rect 487312 5952 487376 5956
rect 522832 6012 522896 6016
rect 522832 5956 522836 6012
rect 522836 5956 522892 6012
rect 522892 5956 522896 6012
rect 522832 5952 522896 5956
rect 522912 6012 522976 6016
rect 522912 5956 522916 6012
rect 522916 5956 522972 6012
rect 522972 5956 522976 6012
rect 522912 5952 522976 5956
rect 522992 6012 523056 6016
rect 522992 5956 522996 6012
rect 522996 5956 523052 6012
rect 523052 5956 523056 6012
rect 522992 5952 523056 5956
rect 523072 6012 523136 6016
rect 523072 5956 523076 6012
rect 523076 5956 523132 6012
rect 523132 5956 523136 6012
rect 523072 5952 523136 5956
rect 523152 6012 523216 6016
rect 523152 5956 523156 6012
rect 523156 5956 523212 6012
rect 523212 5956 523216 6012
rect 523152 5952 523216 5956
rect 523232 6012 523296 6016
rect 523232 5956 523236 6012
rect 523236 5956 523292 6012
rect 523292 5956 523296 6012
rect 523232 5952 523296 5956
rect 523312 6012 523376 6016
rect 523312 5956 523316 6012
rect 523316 5956 523372 6012
rect 523372 5956 523376 6012
rect 523312 5952 523376 5956
rect 558832 6012 558896 6016
rect 558832 5956 558836 6012
rect 558836 5956 558892 6012
rect 558892 5956 558896 6012
rect 558832 5952 558896 5956
rect 558912 6012 558976 6016
rect 558912 5956 558916 6012
rect 558916 5956 558972 6012
rect 558972 5956 558976 6012
rect 558912 5952 558976 5956
rect 558992 6012 559056 6016
rect 558992 5956 558996 6012
rect 558996 5956 559052 6012
rect 559052 5956 559056 6012
rect 558992 5952 559056 5956
rect 559072 6012 559136 6016
rect 559072 5956 559076 6012
rect 559076 5956 559132 6012
rect 559132 5956 559136 6012
rect 559072 5952 559136 5956
rect 559152 6012 559216 6016
rect 559152 5956 559156 6012
rect 559156 5956 559212 6012
rect 559212 5956 559216 6012
rect 559152 5952 559216 5956
rect 559232 6012 559296 6016
rect 559232 5956 559236 6012
rect 559236 5956 559292 6012
rect 559292 5956 559296 6012
rect 559232 5952 559296 5956
rect 559312 6012 559376 6016
rect 559312 5956 559316 6012
rect 559316 5956 559372 6012
rect 559372 5956 559376 6012
rect 559312 5952 559376 5956
rect 36832 5468 36896 5472
rect 36832 5412 36836 5468
rect 36836 5412 36892 5468
rect 36892 5412 36896 5468
rect 36832 5408 36896 5412
rect 36912 5468 36976 5472
rect 36912 5412 36916 5468
rect 36916 5412 36972 5468
rect 36972 5412 36976 5468
rect 36912 5408 36976 5412
rect 36992 5468 37056 5472
rect 36992 5412 36996 5468
rect 36996 5412 37052 5468
rect 37052 5412 37056 5468
rect 36992 5408 37056 5412
rect 37072 5468 37136 5472
rect 37072 5412 37076 5468
rect 37076 5412 37132 5468
rect 37132 5412 37136 5468
rect 37072 5408 37136 5412
rect 37152 5468 37216 5472
rect 37152 5412 37156 5468
rect 37156 5412 37212 5468
rect 37212 5412 37216 5468
rect 37152 5408 37216 5412
rect 37232 5468 37296 5472
rect 37232 5412 37236 5468
rect 37236 5412 37292 5468
rect 37292 5412 37296 5468
rect 37232 5408 37296 5412
rect 37312 5468 37376 5472
rect 37312 5412 37316 5468
rect 37316 5412 37372 5468
rect 37372 5412 37376 5468
rect 37312 5408 37376 5412
rect 72832 5468 72896 5472
rect 72832 5412 72836 5468
rect 72836 5412 72892 5468
rect 72892 5412 72896 5468
rect 72832 5408 72896 5412
rect 72912 5468 72976 5472
rect 72912 5412 72916 5468
rect 72916 5412 72972 5468
rect 72972 5412 72976 5468
rect 72912 5408 72976 5412
rect 72992 5468 73056 5472
rect 72992 5412 72996 5468
rect 72996 5412 73052 5468
rect 73052 5412 73056 5468
rect 72992 5408 73056 5412
rect 73072 5468 73136 5472
rect 73072 5412 73076 5468
rect 73076 5412 73132 5468
rect 73132 5412 73136 5468
rect 73072 5408 73136 5412
rect 73152 5468 73216 5472
rect 73152 5412 73156 5468
rect 73156 5412 73212 5468
rect 73212 5412 73216 5468
rect 73152 5408 73216 5412
rect 73232 5468 73296 5472
rect 73232 5412 73236 5468
rect 73236 5412 73292 5468
rect 73292 5412 73296 5468
rect 73232 5408 73296 5412
rect 73312 5468 73376 5472
rect 73312 5412 73316 5468
rect 73316 5412 73372 5468
rect 73372 5412 73376 5468
rect 73312 5408 73376 5412
rect 108832 5468 108896 5472
rect 108832 5412 108836 5468
rect 108836 5412 108892 5468
rect 108892 5412 108896 5468
rect 108832 5408 108896 5412
rect 108912 5468 108976 5472
rect 108912 5412 108916 5468
rect 108916 5412 108972 5468
rect 108972 5412 108976 5468
rect 108912 5408 108976 5412
rect 108992 5468 109056 5472
rect 108992 5412 108996 5468
rect 108996 5412 109052 5468
rect 109052 5412 109056 5468
rect 108992 5408 109056 5412
rect 109072 5468 109136 5472
rect 109072 5412 109076 5468
rect 109076 5412 109132 5468
rect 109132 5412 109136 5468
rect 109072 5408 109136 5412
rect 109152 5468 109216 5472
rect 109152 5412 109156 5468
rect 109156 5412 109212 5468
rect 109212 5412 109216 5468
rect 109152 5408 109216 5412
rect 109232 5468 109296 5472
rect 109232 5412 109236 5468
rect 109236 5412 109292 5468
rect 109292 5412 109296 5468
rect 109232 5408 109296 5412
rect 109312 5468 109376 5472
rect 109312 5412 109316 5468
rect 109316 5412 109372 5468
rect 109372 5412 109376 5468
rect 109312 5408 109376 5412
rect 144832 5468 144896 5472
rect 144832 5412 144836 5468
rect 144836 5412 144892 5468
rect 144892 5412 144896 5468
rect 144832 5408 144896 5412
rect 144912 5468 144976 5472
rect 144912 5412 144916 5468
rect 144916 5412 144972 5468
rect 144972 5412 144976 5468
rect 144912 5408 144976 5412
rect 144992 5468 145056 5472
rect 144992 5412 144996 5468
rect 144996 5412 145052 5468
rect 145052 5412 145056 5468
rect 144992 5408 145056 5412
rect 145072 5468 145136 5472
rect 145072 5412 145076 5468
rect 145076 5412 145132 5468
rect 145132 5412 145136 5468
rect 145072 5408 145136 5412
rect 145152 5468 145216 5472
rect 145152 5412 145156 5468
rect 145156 5412 145212 5468
rect 145212 5412 145216 5468
rect 145152 5408 145216 5412
rect 145232 5468 145296 5472
rect 145232 5412 145236 5468
rect 145236 5412 145292 5468
rect 145292 5412 145296 5468
rect 145232 5408 145296 5412
rect 145312 5468 145376 5472
rect 145312 5412 145316 5468
rect 145316 5412 145372 5468
rect 145372 5412 145376 5468
rect 145312 5408 145376 5412
rect 180832 5468 180896 5472
rect 180832 5412 180836 5468
rect 180836 5412 180892 5468
rect 180892 5412 180896 5468
rect 180832 5408 180896 5412
rect 180912 5468 180976 5472
rect 180912 5412 180916 5468
rect 180916 5412 180972 5468
rect 180972 5412 180976 5468
rect 180912 5408 180976 5412
rect 180992 5468 181056 5472
rect 180992 5412 180996 5468
rect 180996 5412 181052 5468
rect 181052 5412 181056 5468
rect 180992 5408 181056 5412
rect 181072 5468 181136 5472
rect 181072 5412 181076 5468
rect 181076 5412 181132 5468
rect 181132 5412 181136 5468
rect 181072 5408 181136 5412
rect 181152 5468 181216 5472
rect 181152 5412 181156 5468
rect 181156 5412 181212 5468
rect 181212 5412 181216 5468
rect 181152 5408 181216 5412
rect 181232 5468 181296 5472
rect 181232 5412 181236 5468
rect 181236 5412 181292 5468
rect 181292 5412 181296 5468
rect 181232 5408 181296 5412
rect 181312 5468 181376 5472
rect 181312 5412 181316 5468
rect 181316 5412 181372 5468
rect 181372 5412 181376 5468
rect 181312 5408 181376 5412
rect 216832 5468 216896 5472
rect 216832 5412 216836 5468
rect 216836 5412 216892 5468
rect 216892 5412 216896 5468
rect 216832 5408 216896 5412
rect 216912 5468 216976 5472
rect 216912 5412 216916 5468
rect 216916 5412 216972 5468
rect 216972 5412 216976 5468
rect 216912 5408 216976 5412
rect 216992 5468 217056 5472
rect 216992 5412 216996 5468
rect 216996 5412 217052 5468
rect 217052 5412 217056 5468
rect 216992 5408 217056 5412
rect 217072 5468 217136 5472
rect 217072 5412 217076 5468
rect 217076 5412 217132 5468
rect 217132 5412 217136 5468
rect 217072 5408 217136 5412
rect 217152 5468 217216 5472
rect 217152 5412 217156 5468
rect 217156 5412 217212 5468
rect 217212 5412 217216 5468
rect 217152 5408 217216 5412
rect 217232 5468 217296 5472
rect 217232 5412 217236 5468
rect 217236 5412 217292 5468
rect 217292 5412 217296 5468
rect 217232 5408 217296 5412
rect 217312 5468 217376 5472
rect 217312 5412 217316 5468
rect 217316 5412 217372 5468
rect 217372 5412 217376 5468
rect 217312 5408 217376 5412
rect 252832 5468 252896 5472
rect 252832 5412 252836 5468
rect 252836 5412 252892 5468
rect 252892 5412 252896 5468
rect 252832 5408 252896 5412
rect 252912 5468 252976 5472
rect 252912 5412 252916 5468
rect 252916 5412 252972 5468
rect 252972 5412 252976 5468
rect 252912 5408 252976 5412
rect 252992 5468 253056 5472
rect 252992 5412 252996 5468
rect 252996 5412 253052 5468
rect 253052 5412 253056 5468
rect 252992 5408 253056 5412
rect 253072 5468 253136 5472
rect 253072 5412 253076 5468
rect 253076 5412 253132 5468
rect 253132 5412 253136 5468
rect 253072 5408 253136 5412
rect 253152 5468 253216 5472
rect 253152 5412 253156 5468
rect 253156 5412 253212 5468
rect 253212 5412 253216 5468
rect 253152 5408 253216 5412
rect 253232 5468 253296 5472
rect 253232 5412 253236 5468
rect 253236 5412 253292 5468
rect 253292 5412 253296 5468
rect 253232 5408 253296 5412
rect 253312 5468 253376 5472
rect 253312 5412 253316 5468
rect 253316 5412 253372 5468
rect 253372 5412 253376 5468
rect 253312 5408 253376 5412
rect 288832 5468 288896 5472
rect 288832 5412 288836 5468
rect 288836 5412 288892 5468
rect 288892 5412 288896 5468
rect 288832 5408 288896 5412
rect 288912 5468 288976 5472
rect 288912 5412 288916 5468
rect 288916 5412 288972 5468
rect 288972 5412 288976 5468
rect 288912 5408 288976 5412
rect 288992 5468 289056 5472
rect 288992 5412 288996 5468
rect 288996 5412 289052 5468
rect 289052 5412 289056 5468
rect 288992 5408 289056 5412
rect 289072 5468 289136 5472
rect 289072 5412 289076 5468
rect 289076 5412 289132 5468
rect 289132 5412 289136 5468
rect 289072 5408 289136 5412
rect 289152 5468 289216 5472
rect 289152 5412 289156 5468
rect 289156 5412 289212 5468
rect 289212 5412 289216 5468
rect 289152 5408 289216 5412
rect 289232 5468 289296 5472
rect 289232 5412 289236 5468
rect 289236 5412 289292 5468
rect 289292 5412 289296 5468
rect 289232 5408 289296 5412
rect 289312 5468 289376 5472
rect 289312 5412 289316 5468
rect 289316 5412 289372 5468
rect 289372 5412 289376 5468
rect 289312 5408 289376 5412
rect 324832 5468 324896 5472
rect 324832 5412 324836 5468
rect 324836 5412 324892 5468
rect 324892 5412 324896 5468
rect 324832 5408 324896 5412
rect 324912 5468 324976 5472
rect 324912 5412 324916 5468
rect 324916 5412 324972 5468
rect 324972 5412 324976 5468
rect 324912 5408 324976 5412
rect 324992 5468 325056 5472
rect 324992 5412 324996 5468
rect 324996 5412 325052 5468
rect 325052 5412 325056 5468
rect 324992 5408 325056 5412
rect 325072 5468 325136 5472
rect 325072 5412 325076 5468
rect 325076 5412 325132 5468
rect 325132 5412 325136 5468
rect 325072 5408 325136 5412
rect 325152 5468 325216 5472
rect 325152 5412 325156 5468
rect 325156 5412 325212 5468
rect 325212 5412 325216 5468
rect 325152 5408 325216 5412
rect 325232 5468 325296 5472
rect 325232 5412 325236 5468
rect 325236 5412 325292 5468
rect 325292 5412 325296 5468
rect 325232 5408 325296 5412
rect 325312 5468 325376 5472
rect 325312 5412 325316 5468
rect 325316 5412 325372 5468
rect 325372 5412 325376 5468
rect 325312 5408 325376 5412
rect 360832 5468 360896 5472
rect 360832 5412 360836 5468
rect 360836 5412 360892 5468
rect 360892 5412 360896 5468
rect 360832 5408 360896 5412
rect 360912 5468 360976 5472
rect 360912 5412 360916 5468
rect 360916 5412 360972 5468
rect 360972 5412 360976 5468
rect 360912 5408 360976 5412
rect 360992 5468 361056 5472
rect 360992 5412 360996 5468
rect 360996 5412 361052 5468
rect 361052 5412 361056 5468
rect 360992 5408 361056 5412
rect 361072 5468 361136 5472
rect 361072 5412 361076 5468
rect 361076 5412 361132 5468
rect 361132 5412 361136 5468
rect 361072 5408 361136 5412
rect 361152 5468 361216 5472
rect 361152 5412 361156 5468
rect 361156 5412 361212 5468
rect 361212 5412 361216 5468
rect 361152 5408 361216 5412
rect 361232 5468 361296 5472
rect 361232 5412 361236 5468
rect 361236 5412 361292 5468
rect 361292 5412 361296 5468
rect 361232 5408 361296 5412
rect 361312 5468 361376 5472
rect 361312 5412 361316 5468
rect 361316 5412 361372 5468
rect 361372 5412 361376 5468
rect 361312 5408 361376 5412
rect 396832 5468 396896 5472
rect 396832 5412 396836 5468
rect 396836 5412 396892 5468
rect 396892 5412 396896 5468
rect 396832 5408 396896 5412
rect 396912 5468 396976 5472
rect 396912 5412 396916 5468
rect 396916 5412 396972 5468
rect 396972 5412 396976 5468
rect 396912 5408 396976 5412
rect 396992 5468 397056 5472
rect 396992 5412 396996 5468
rect 396996 5412 397052 5468
rect 397052 5412 397056 5468
rect 396992 5408 397056 5412
rect 397072 5468 397136 5472
rect 397072 5412 397076 5468
rect 397076 5412 397132 5468
rect 397132 5412 397136 5468
rect 397072 5408 397136 5412
rect 397152 5468 397216 5472
rect 397152 5412 397156 5468
rect 397156 5412 397212 5468
rect 397212 5412 397216 5468
rect 397152 5408 397216 5412
rect 397232 5468 397296 5472
rect 397232 5412 397236 5468
rect 397236 5412 397292 5468
rect 397292 5412 397296 5468
rect 397232 5408 397296 5412
rect 397312 5468 397376 5472
rect 397312 5412 397316 5468
rect 397316 5412 397372 5468
rect 397372 5412 397376 5468
rect 397312 5408 397376 5412
rect 432832 5468 432896 5472
rect 432832 5412 432836 5468
rect 432836 5412 432892 5468
rect 432892 5412 432896 5468
rect 432832 5408 432896 5412
rect 432912 5468 432976 5472
rect 432912 5412 432916 5468
rect 432916 5412 432972 5468
rect 432972 5412 432976 5468
rect 432912 5408 432976 5412
rect 432992 5468 433056 5472
rect 432992 5412 432996 5468
rect 432996 5412 433052 5468
rect 433052 5412 433056 5468
rect 432992 5408 433056 5412
rect 433072 5468 433136 5472
rect 433072 5412 433076 5468
rect 433076 5412 433132 5468
rect 433132 5412 433136 5468
rect 433072 5408 433136 5412
rect 433152 5468 433216 5472
rect 433152 5412 433156 5468
rect 433156 5412 433212 5468
rect 433212 5412 433216 5468
rect 433152 5408 433216 5412
rect 433232 5468 433296 5472
rect 433232 5412 433236 5468
rect 433236 5412 433292 5468
rect 433292 5412 433296 5468
rect 433232 5408 433296 5412
rect 433312 5468 433376 5472
rect 433312 5412 433316 5468
rect 433316 5412 433372 5468
rect 433372 5412 433376 5468
rect 433312 5408 433376 5412
rect 468832 5468 468896 5472
rect 468832 5412 468836 5468
rect 468836 5412 468892 5468
rect 468892 5412 468896 5468
rect 468832 5408 468896 5412
rect 468912 5468 468976 5472
rect 468912 5412 468916 5468
rect 468916 5412 468972 5468
rect 468972 5412 468976 5468
rect 468912 5408 468976 5412
rect 468992 5468 469056 5472
rect 468992 5412 468996 5468
rect 468996 5412 469052 5468
rect 469052 5412 469056 5468
rect 468992 5408 469056 5412
rect 469072 5468 469136 5472
rect 469072 5412 469076 5468
rect 469076 5412 469132 5468
rect 469132 5412 469136 5468
rect 469072 5408 469136 5412
rect 469152 5468 469216 5472
rect 469152 5412 469156 5468
rect 469156 5412 469212 5468
rect 469212 5412 469216 5468
rect 469152 5408 469216 5412
rect 469232 5468 469296 5472
rect 469232 5412 469236 5468
rect 469236 5412 469292 5468
rect 469292 5412 469296 5468
rect 469232 5408 469296 5412
rect 469312 5468 469376 5472
rect 469312 5412 469316 5468
rect 469316 5412 469372 5468
rect 469372 5412 469376 5468
rect 469312 5408 469376 5412
rect 504832 5468 504896 5472
rect 504832 5412 504836 5468
rect 504836 5412 504892 5468
rect 504892 5412 504896 5468
rect 504832 5408 504896 5412
rect 504912 5468 504976 5472
rect 504912 5412 504916 5468
rect 504916 5412 504972 5468
rect 504972 5412 504976 5468
rect 504912 5408 504976 5412
rect 504992 5468 505056 5472
rect 504992 5412 504996 5468
rect 504996 5412 505052 5468
rect 505052 5412 505056 5468
rect 504992 5408 505056 5412
rect 505072 5468 505136 5472
rect 505072 5412 505076 5468
rect 505076 5412 505132 5468
rect 505132 5412 505136 5468
rect 505072 5408 505136 5412
rect 505152 5468 505216 5472
rect 505152 5412 505156 5468
rect 505156 5412 505212 5468
rect 505212 5412 505216 5468
rect 505152 5408 505216 5412
rect 505232 5468 505296 5472
rect 505232 5412 505236 5468
rect 505236 5412 505292 5468
rect 505292 5412 505296 5468
rect 505232 5408 505296 5412
rect 505312 5468 505376 5472
rect 505312 5412 505316 5468
rect 505316 5412 505372 5468
rect 505372 5412 505376 5468
rect 505312 5408 505376 5412
rect 540832 5468 540896 5472
rect 540832 5412 540836 5468
rect 540836 5412 540892 5468
rect 540892 5412 540896 5468
rect 540832 5408 540896 5412
rect 540912 5468 540976 5472
rect 540912 5412 540916 5468
rect 540916 5412 540972 5468
rect 540972 5412 540976 5468
rect 540912 5408 540976 5412
rect 540992 5468 541056 5472
rect 540992 5412 540996 5468
rect 540996 5412 541052 5468
rect 541052 5412 541056 5468
rect 540992 5408 541056 5412
rect 541072 5468 541136 5472
rect 541072 5412 541076 5468
rect 541076 5412 541132 5468
rect 541132 5412 541136 5468
rect 541072 5408 541136 5412
rect 541152 5468 541216 5472
rect 541152 5412 541156 5468
rect 541156 5412 541212 5468
rect 541212 5412 541216 5468
rect 541152 5408 541216 5412
rect 541232 5468 541296 5472
rect 541232 5412 541236 5468
rect 541236 5412 541292 5468
rect 541292 5412 541296 5468
rect 541232 5408 541296 5412
rect 541312 5468 541376 5472
rect 541312 5412 541316 5468
rect 541316 5412 541372 5468
rect 541372 5412 541376 5468
rect 541312 5408 541376 5412
rect 576832 5468 576896 5472
rect 576832 5412 576836 5468
rect 576836 5412 576892 5468
rect 576892 5412 576896 5468
rect 576832 5408 576896 5412
rect 576912 5468 576976 5472
rect 576912 5412 576916 5468
rect 576916 5412 576972 5468
rect 576972 5412 576976 5468
rect 576912 5408 576976 5412
rect 576992 5468 577056 5472
rect 576992 5412 576996 5468
rect 576996 5412 577052 5468
rect 577052 5412 577056 5468
rect 576992 5408 577056 5412
rect 577072 5468 577136 5472
rect 577072 5412 577076 5468
rect 577076 5412 577132 5468
rect 577132 5412 577136 5468
rect 577072 5408 577136 5412
rect 577152 5468 577216 5472
rect 577152 5412 577156 5468
rect 577156 5412 577212 5468
rect 577212 5412 577216 5468
rect 577152 5408 577216 5412
rect 577232 5468 577296 5472
rect 577232 5412 577236 5468
rect 577236 5412 577292 5468
rect 577292 5412 577296 5468
rect 577232 5408 577296 5412
rect 577312 5468 577376 5472
rect 577312 5412 577316 5468
rect 577316 5412 577372 5468
rect 577372 5412 577376 5468
rect 577312 5408 577376 5412
rect 18832 4924 18896 4928
rect 18832 4868 18836 4924
rect 18836 4868 18892 4924
rect 18892 4868 18896 4924
rect 18832 4864 18896 4868
rect 18912 4924 18976 4928
rect 18912 4868 18916 4924
rect 18916 4868 18972 4924
rect 18972 4868 18976 4924
rect 18912 4864 18976 4868
rect 18992 4924 19056 4928
rect 18992 4868 18996 4924
rect 18996 4868 19052 4924
rect 19052 4868 19056 4924
rect 18992 4864 19056 4868
rect 19072 4924 19136 4928
rect 19072 4868 19076 4924
rect 19076 4868 19132 4924
rect 19132 4868 19136 4924
rect 19072 4864 19136 4868
rect 19152 4924 19216 4928
rect 19152 4868 19156 4924
rect 19156 4868 19212 4924
rect 19212 4868 19216 4924
rect 19152 4864 19216 4868
rect 19232 4924 19296 4928
rect 19232 4868 19236 4924
rect 19236 4868 19292 4924
rect 19292 4868 19296 4924
rect 19232 4864 19296 4868
rect 19312 4924 19376 4928
rect 19312 4868 19316 4924
rect 19316 4868 19372 4924
rect 19372 4868 19376 4924
rect 19312 4864 19376 4868
rect 54832 4924 54896 4928
rect 54832 4868 54836 4924
rect 54836 4868 54892 4924
rect 54892 4868 54896 4924
rect 54832 4864 54896 4868
rect 54912 4924 54976 4928
rect 54912 4868 54916 4924
rect 54916 4868 54972 4924
rect 54972 4868 54976 4924
rect 54912 4864 54976 4868
rect 54992 4924 55056 4928
rect 54992 4868 54996 4924
rect 54996 4868 55052 4924
rect 55052 4868 55056 4924
rect 54992 4864 55056 4868
rect 55072 4924 55136 4928
rect 55072 4868 55076 4924
rect 55076 4868 55132 4924
rect 55132 4868 55136 4924
rect 55072 4864 55136 4868
rect 55152 4924 55216 4928
rect 55152 4868 55156 4924
rect 55156 4868 55212 4924
rect 55212 4868 55216 4924
rect 55152 4864 55216 4868
rect 55232 4924 55296 4928
rect 55232 4868 55236 4924
rect 55236 4868 55292 4924
rect 55292 4868 55296 4924
rect 55232 4864 55296 4868
rect 55312 4924 55376 4928
rect 55312 4868 55316 4924
rect 55316 4868 55372 4924
rect 55372 4868 55376 4924
rect 55312 4864 55376 4868
rect 90832 4924 90896 4928
rect 90832 4868 90836 4924
rect 90836 4868 90892 4924
rect 90892 4868 90896 4924
rect 90832 4864 90896 4868
rect 90912 4924 90976 4928
rect 90912 4868 90916 4924
rect 90916 4868 90972 4924
rect 90972 4868 90976 4924
rect 90912 4864 90976 4868
rect 90992 4924 91056 4928
rect 90992 4868 90996 4924
rect 90996 4868 91052 4924
rect 91052 4868 91056 4924
rect 90992 4864 91056 4868
rect 91072 4924 91136 4928
rect 91072 4868 91076 4924
rect 91076 4868 91132 4924
rect 91132 4868 91136 4924
rect 91072 4864 91136 4868
rect 91152 4924 91216 4928
rect 91152 4868 91156 4924
rect 91156 4868 91212 4924
rect 91212 4868 91216 4924
rect 91152 4864 91216 4868
rect 91232 4924 91296 4928
rect 91232 4868 91236 4924
rect 91236 4868 91292 4924
rect 91292 4868 91296 4924
rect 91232 4864 91296 4868
rect 91312 4924 91376 4928
rect 91312 4868 91316 4924
rect 91316 4868 91372 4924
rect 91372 4868 91376 4924
rect 91312 4864 91376 4868
rect 126832 4924 126896 4928
rect 126832 4868 126836 4924
rect 126836 4868 126892 4924
rect 126892 4868 126896 4924
rect 126832 4864 126896 4868
rect 126912 4924 126976 4928
rect 126912 4868 126916 4924
rect 126916 4868 126972 4924
rect 126972 4868 126976 4924
rect 126912 4864 126976 4868
rect 126992 4924 127056 4928
rect 126992 4868 126996 4924
rect 126996 4868 127052 4924
rect 127052 4868 127056 4924
rect 126992 4864 127056 4868
rect 127072 4924 127136 4928
rect 127072 4868 127076 4924
rect 127076 4868 127132 4924
rect 127132 4868 127136 4924
rect 127072 4864 127136 4868
rect 127152 4924 127216 4928
rect 127152 4868 127156 4924
rect 127156 4868 127212 4924
rect 127212 4868 127216 4924
rect 127152 4864 127216 4868
rect 127232 4924 127296 4928
rect 127232 4868 127236 4924
rect 127236 4868 127292 4924
rect 127292 4868 127296 4924
rect 127232 4864 127296 4868
rect 127312 4924 127376 4928
rect 127312 4868 127316 4924
rect 127316 4868 127372 4924
rect 127372 4868 127376 4924
rect 127312 4864 127376 4868
rect 162832 4924 162896 4928
rect 162832 4868 162836 4924
rect 162836 4868 162892 4924
rect 162892 4868 162896 4924
rect 162832 4864 162896 4868
rect 162912 4924 162976 4928
rect 162912 4868 162916 4924
rect 162916 4868 162972 4924
rect 162972 4868 162976 4924
rect 162912 4864 162976 4868
rect 162992 4924 163056 4928
rect 162992 4868 162996 4924
rect 162996 4868 163052 4924
rect 163052 4868 163056 4924
rect 162992 4864 163056 4868
rect 163072 4924 163136 4928
rect 163072 4868 163076 4924
rect 163076 4868 163132 4924
rect 163132 4868 163136 4924
rect 163072 4864 163136 4868
rect 163152 4924 163216 4928
rect 163152 4868 163156 4924
rect 163156 4868 163212 4924
rect 163212 4868 163216 4924
rect 163152 4864 163216 4868
rect 163232 4924 163296 4928
rect 163232 4868 163236 4924
rect 163236 4868 163292 4924
rect 163292 4868 163296 4924
rect 163232 4864 163296 4868
rect 163312 4924 163376 4928
rect 163312 4868 163316 4924
rect 163316 4868 163372 4924
rect 163372 4868 163376 4924
rect 163312 4864 163376 4868
rect 198832 4924 198896 4928
rect 198832 4868 198836 4924
rect 198836 4868 198892 4924
rect 198892 4868 198896 4924
rect 198832 4864 198896 4868
rect 198912 4924 198976 4928
rect 198912 4868 198916 4924
rect 198916 4868 198972 4924
rect 198972 4868 198976 4924
rect 198912 4864 198976 4868
rect 198992 4924 199056 4928
rect 198992 4868 198996 4924
rect 198996 4868 199052 4924
rect 199052 4868 199056 4924
rect 198992 4864 199056 4868
rect 199072 4924 199136 4928
rect 199072 4868 199076 4924
rect 199076 4868 199132 4924
rect 199132 4868 199136 4924
rect 199072 4864 199136 4868
rect 199152 4924 199216 4928
rect 199152 4868 199156 4924
rect 199156 4868 199212 4924
rect 199212 4868 199216 4924
rect 199152 4864 199216 4868
rect 199232 4924 199296 4928
rect 199232 4868 199236 4924
rect 199236 4868 199292 4924
rect 199292 4868 199296 4924
rect 199232 4864 199296 4868
rect 199312 4924 199376 4928
rect 199312 4868 199316 4924
rect 199316 4868 199372 4924
rect 199372 4868 199376 4924
rect 199312 4864 199376 4868
rect 234832 4924 234896 4928
rect 234832 4868 234836 4924
rect 234836 4868 234892 4924
rect 234892 4868 234896 4924
rect 234832 4864 234896 4868
rect 234912 4924 234976 4928
rect 234912 4868 234916 4924
rect 234916 4868 234972 4924
rect 234972 4868 234976 4924
rect 234912 4864 234976 4868
rect 234992 4924 235056 4928
rect 234992 4868 234996 4924
rect 234996 4868 235052 4924
rect 235052 4868 235056 4924
rect 234992 4864 235056 4868
rect 235072 4924 235136 4928
rect 235072 4868 235076 4924
rect 235076 4868 235132 4924
rect 235132 4868 235136 4924
rect 235072 4864 235136 4868
rect 235152 4924 235216 4928
rect 235152 4868 235156 4924
rect 235156 4868 235212 4924
rect 235212 4868 235216 4924
rect 235152 4864 235216 4868
rect 235232 4924 235296 4928
rect 235232 4868 235236 4924
rect 235236 4868 235292 4924
rect 235292 4868 235296 4924
rect 235232 4864 235296 4868
rect 235312 4924 235376 4928
rect 235312 4868 235316 4924
rect 235316 4868 235372 4924
rect 235372 4868 235376 4924
rect 235312 4864 235376 4868
rect 270832 4924 270896 4928
rect 270832 4868 270836 4924
rect 270836 4868 270892 4924
rect 270892 4868 270896 4924
rect 270832 4864 270896 4868
rect 270912 4924 270976 4928
rect 270912 4868 270916 4924
rect 270916 4868 270972 4924
rect 270972 4868 270976 4924
rect 270912 4864 270976 4868
rect 270992 4924 271056 4928
rect 270992 4868 270996 4924
rect 270996 4868 271052 4924
rect 271052 4868 271056 4924
rect 270992 4864 271056 4868
rect 271072 4924 271136 4928
rect 271072 4868 271076 4924
rect 271076 4868 271132 4924
rect 271132 4868 271136 4924
rect 271072 4864 271136 4868
rect 271152 4924 271216 4928
rect 271152 4868 271156 4924
rect 271156 4868 271212 4924
rect 271212 4868 271216 4924
rect 271152 4864 271216 4868
rect 271232 4924 271296 4928
rect 271232 4868 271236 4924
rect 271236 4868 271292 4924
rect 271292 4868 271296 4924
rect 271232 4864 271296 4868
rect 271312 4924 271376 4928
rect 271312 4868 271316 4924
rect 271316 4868 271372 4924
rect 271372 4868 271376 4924
rect 271312 4864 271376 4868
rect 306832 4924 306896 4928
rect 306832 4868 306836 4924
rect 306836 4868 306892 4924
rect 306892 4868 306896 4924
rect 306832 4864 306896 4868
rect 306912 4924 306976 4928
rect 306912 4868 306916 4924
rect 306916 4868 306972 4924
rect 306972 4868 306976 4924
rect 306912 4864 306976 4868
rect 306992 4924 307056 4928
rect 306992 4868 306996 4924
rect 306996 4868 307052 4924
rect 307052 4868 307056 4924
rect 306992 4864 307056 4868
rect 307072 4924 307136 4928
rect 307072 4868 307076 4924
rect 307076 4868 307132 4924
rect 307132 4868 307136 4924
rect 307072 4864 307136 4868
rect 307152 4924 307216 4928
rect 307152 4868 307156 4924
rect 307156 4868 307212 4924
rect 307212 4868 307216 4924
rect 307152 4864 307216 4868
rect 307232 4924 307296 4928
rect 307232 4868 307236 4924
rect 307236 4868 307292 4924
rect 307292 4868 307296 4924
rect 307232 4864 307296 4868
rect 307312 4924 307376 4928
rect 307312 4868 307316 4924
rect 307316 4868 307372 4924
rect 307372 4868 307376 4924
rect 307312 4864 307376 4868
rect 342832 4924 342896 4928
rect 342832 4868 342836 4924
rect 342836 4868 342892 4924
rect 342892 4868 342896 4924
rect 342832 4864 342896 4868
rect 342912 4924 342976 4928
rect 342912 4868 342916 4924
rect 342916 4868 342972 4924
rect 342972 4868 342976 4924
rect 342912 4864 342976 4868
rect 342992 4924 343056 4928
rect 342992 4868 342996 4924
rect 342996 4868 343052 4924
rect 343052 4868 343056 4924
rect 342992 4864 343056 4868
rect 343072 4924 343136 4928
rect 343072 4868 343076 4924
rect 343076 4868 343132 4924
rect 343132 4868 343136 4924
rect 343072 4864 343136 4868
rect 343152 4924 343216 4928
rect 343152 4868 343156 4924
rect 343156 4868 343212 4924
rect 343212 4868 343216 4924
rect 343152 4864 343216 4868
rect 343232 4924 343296 4928
rect 343232 4868 343236 4924
rect 343236 4868 343292 4924
rect 343292 4868 343296 4924
rect 343232 4864 343296 4868
rect 343312 4924 343376 4928
rect 343312 4868 343316 4924
rect 343316 4868 343372 4924
rect 343372 4868 343376 4924
rect 343312 4864 343376 4868
rect 378832 4924 378896 4928
rect 378832 4868 378836 4924
rect 378836 4868 378892 4924
rect 378892 4868 378896 4924
rect 378832 4864 378896 4868
rect 378912 4924 378976 4928
rect 378912 4868 378916 4924
rect 378916 4868 378972 4924
rect 378972 4868 378976 4924
rect 378912 4864 378976 4868
rect 378992 4924 379056 4928
rect 378992 4868 378996 4924
rect 378996 4868 379052 4924
rect 379052 4868 379056 4924
rect 378992 4864 379056 4868
rect 379072 4924 379136 4928
rect 379072 4868 379076 4924
rect 379076 4868 379132 4924
rect 379132 4868 379136 4924
rect 379072 4864 379136 4868
rect 379152 4924 379216 4928
rect 379152 4868 379156 4924
rect 379156 4868 379212 4924
rect 379212 4868 379216 4924
rect 379152 4864 379216 4868
rect 379232 4924 379296 4928
rect 379232 4868 379236 4924
rect 379236 4868 379292 4924
rect 379292 4868 379296 4924
rect 379232 4864 379296 4868
rect 379312 4924 379376 4928
rect 379312 4868 379316 4924
rect 379316 4868 379372 4924
rect 379372 4868 379376 4924
rect 379312 4864 379376 4868
rect 414832 4924 414896 4928
rect 414832 4868 414836 4924
rect 414836 4868 414892 4924
rect 414892 4868 414896 4924
rect 414832 4864 414896 4868
rect 414912 4924 414976 4928
rect 414912 4868 414916 4924
rect 414916 4868 414972 4924
rect 414972 4868 414976 4924
rect 414912 4864 414976 4868
rect 414992 4924 415056 4928
rect 414992 4868 414996 4924
rect 414996 4868 415052 4924
rect 415052 4868 415056 4924
rect 414992 4864 415056 4868
rect 415072 4924 415136 4928
rect 415072 4868 415076 4924
rect 415076 4868 415132 4924
rect 415132 4868 415136 4924
rect 415072 4864 415136 4868
rect 415152 4924 415216 4928
rect 415152 4868 415156 4924
rect 415156 4868 415212 4924
rect 415212 4868 415216 4924
rect 415152 4864 415216 4868
rect 415232 4924 415296 4928
rect 415232 4868 415236 4924
rect 415236 4868 415292 4924
rect 415292 4868 415296 4924
rect 415232 4864 415296 4868
rect 415312 4924 415376 4928
rect 415312 4868 415316 4924
rect 415316 4868 415372 4924
rect 415372 4868 415376 4924
rect 415312 4864 415376 4868
rect 450832 4924 450896 4928
rect 450832 4868 450836 4924
rect 450836 4868 450892 4924
rect 450892 4868 450896 4924
rect 450832 4864 450896 4868
rect 450912 4924 450976 4928
rect 450912 4868 450916 4924
rect 450916 4868 450972 4924
rect 450972 4868 450976 4924
rect 450912 4864 450976 4868
rect 450992 4924 451056 4928
rect 450992 4868 450996 4924
rect 450996 4868 451052 4924
rect 451052 4868 451056 4924
rect 450992 4864 451056 4868
rect 451072 4924 451136 4928
rect 451072 4868 451076 4924
rect 451076 4868 451132 4924
rect 451132 4868 451136 4924
rect 451072 4864 451136 4868
rect 451152 4924 451216 4928
rect 451152 4868 451156 4924
rect 451156 4868 451212 4924
rect 451212 4868 451216 4924
rect 451152 4864 451216 4868
rect 451232 4924 451296 4928
rect 451232 4868 451236 4924
rect 451236 4868 451292 4924
rect 451292 4868 451296 4924
rect 451232 4864 451296 4868
rect 451312 4924 451376 4928
rect 451312 4868 451316 4924
rect 451316 4868 451372 4924
rect 451372 4868 451376 4924
rect 451312 4864 451376 4868
rect 486832 4924 486896 4928
rect 486832 4868 486836 4924
rect 486836 4868 486892 4924
rect 486892 4868 486896 4924
rect 486832 4864 486896 4868
rect 486912 4924 486976 4928
rect 486912 4868 486916 4924
rect 486916 4868 486972 4924
rect 486972 4868 486976 4924
rect 486912 4864 486976 4868
rect 486992 4924 487056 4928
rect 486992 4868 486996 4924
rect 486996 4868 487052 4924
rect 487052 4868 487056 4924
rect 486992 4864 487056 4868
rect 487072 4924 487136 4928
rect 487072 4868 487076 4924
rect 487076 4868 487132 4924
rect 487132 4868 487136 4924
rect 487072 4864 487136 4868
rect 487152 4924 487216 4928
rect 487152 4868 487156 4924
rect 487156 4868 487212 4924
rect 487212 4868 487216 4924
rect 487152 4864 487216 4868
rect 487232 4924 487296 4928
rect 487232 4868 487236 4924
rect 487236 4868 487292 4924
rect 487292 4868 487296 4924
rect 487232 4864 487296 4868
rect 487312 4924 487376 4928
rect 487312 4868 487316 4924
rect 487316 4868 487372 4924
rect 487372 4868 487376 4924
rect 487312 4864 487376 4868
rect 522832 4924 522896 4928
rect 522832 4868 522836 4924
rect 522836 4868 522892 4924
rect 522892 4868 522896 4924
rect 522832 4864 522896 4868
rect 522912 4924 522976 4928
rect 522912 4868 522916 4924
rect 522916 4868 522972 4924
rect 522972 4868 522976 4924
rect 522912 4864 522976 4868
rect 522992 4924 523056 4928
rect 522992 4868 522996 4924
rect 522996 4868 523052 4924
rect 523052 4868 523056 4924
rect 522992 4864 523056 4868
rect 523072 4924 523136 4928
rect 523072 4868 523076 4924
rect 523076 4868 523132 4924
rect 523132 4868 523136 4924
rect 523072 4864 523136 4868
rect 523152 4924 523216 4928
rect 523152 4868 523156 4924
rect 523156 4868 523212 4924
rect 523212 4868 523216 4924
rect 523152 4864 523216 4868
rect 523232 4924 523296 4928
rect 523232 4868 523236 4924
rect 523236 4868 523292 4924
rect 523292 4868 523296 4924
rect 523232 4864 523296 4868
rect 523312 4924 523376 4928
rect 523312 4868 523316 4924
rect 523316 4868 523372 4924
rect 523372 4868 523376 4924
rect 523312 4864 523376 4868
rect 558832 4924 558896 4928
rect 558832 4868 558836 4924
rect 558836 4868 558892 4924
rect 558892 4868 558896 4924
rect 558832 4864 558896 4868
rect 558912 4924 558976 4928
rect 558912 4868 558916 4924
rect 558916 4868 558972 4924
rect 558972 4868 558976 4924
rect 558912 4864 558976 4868
rect 558992 4924 559056 4928
rect 558992 4868 558996 4924
rect 558996 4868 559052 4924
rect 559052 4868 559056 4924
rect 558992 4864 559056 4868
rect 559072 4924 559136 4928
rect 559072 4868 559076 4924
rect 559076 4868 559132 4924
rect 559132 4868 559136 4924
rect 559072 4864 559136 4868
rect 559152 4924 559216 4928
rect 559152 4868 559156 4924
rect 559156 4868 559212 4924
rect 559212 4868 559216 4924
rect 559152 4864 559216 4868
rect 559232 4924 559296 4928
rect 559232 4868 559236 4924
rect 559236 4868 559292 4924
rect 559292 4868 559296 4924
rect 559232 4864 559296 4868
rect 559312 4924 559376 4928
rect 559312 4868 559316 4924
rect 559316 4868 559372 4924
rect 559372 4868 559376 4924
rect 559312 4864 559376 4868
rect 36832 4380 36896 4384
rect 36832 4324 36836 4380
rect 36836 4324 36892 4380
rect 36892 4324 36896 4380
rect 36832 4320 36896 4324
rect 36912 4380 36976 4384
rect 36912 4324 36916 4380
rect 36916 4324 36972 4380
rect 36972 4324 36976 4380
rect 36912 4320 36976 4324
rect 36992 4380 37056 4384
rect 36992 4324 36996 4380
rect 36996 4324 37052 4380
rect 37052 4324 37056 4380
rect 36992 4320 37056 4324
rect 37072 4380 37136 4384
rect 37072 4324 37076 4380
rect 37076 4324 37132 4380
rect 37132 4324 37136 4380
rect 37072 4320 37136 4324
rect 37152 4380 37216 4384
rect 37152 4324 37156 4380
rect 37156 4324 37212 4380
rect 37212 4324 37216 4380
rect 37152 4320 37216 4324
rect 37232 4380 37296 4384
rect 37232 4324 37236 4380
rect 37236 4324 37292 4380
rect 37292 4324 37296 4380
rect 37232 4320 37296 4324
rect 37312 4380 37376 4384
rect 37312 4324 37316 4380
rect 37316 4324 37372 4380
rect 37372 4324 37376 4380
rect 37312 4320 37376 4324
rect 72832 4380 72896 4384
rect 72832 4324 72836 4380
rect 72836 4324 72892 4380
rect 72892 4324 72896 4380
rect 72832 4320 72896 4324
rect 72912 4380 72976 4384
rect 72912 4324 72916 4380
rect 72916 4324 72972 4380
rect 72972 4324 72976 4380
rect 72912 4320 72976 4324
rect 72992 4380 73056 4384
rect 72992 4324 72996 4380
rect 72996 4324 73052 4380
rect 73052 4324 73056 4380
rect 72992 4320 73056 4324
rect 73072 4380 73136 4384
rect 73072 4324 73076 4380
rect 73076 4324 73132 4380
rect 73132 4324 73136 4380
rect 73072 4320 73136 4324
rect 73152 4380 73216 4384
rect 73152 4324 73156 4380
rect 73156 4324 73212 4380
rect 73212 4324 73216 4380
rect 73152 4320 73216 4324
rect 73232 4380 73296 4384
rect 73232 4324 73236 4380
rect 73236 4324 73292 4380
rect 73292 4324 73296 4380
rect 73232 4320 73296 4324
rect 73312 4380 73376 4384
rect 73312 4324 73316 4380
rect 73316 4324 73372 4380
rect 73372 4324 73376 4380
rect 73312 4320 73376 4324
rect 108832 4380 108896 4384
rect 108832 4324 108836 4380
rect 108836 4324 108892 4380
rect 108892 4324 108896 4380
rect 108832 4320 108896 4324
rect 108912 4380 108976 4384
rect 108912 4324 108916 4380
rect 108916 4324 108972 4380
rect 108972 4324 108976 4380
rect 108912 4320 108976 4324
rect 108992 4380 109056 4384
rect 108992 4324 108996 4380
rect 108996 4324 109052 4380
rect 109052 4324 109056 4380
rect 108992 4320 109056 4324
rect 109072 4380 109136 4384
rect 109072 4324 109076 4380
rect 109076 4324 109132 4380
rect 109132 4324 109136 4380
rect 109072 4320 109136 4324
rect 109152 4380 109216 4384
rect 109152 4324 109156 4380
rect 109156 4324 109212 4380
rect 109212 4324 109216 4380
rect 109152 4320 109216 4324
rect 109232 4380 109296 4384
rect 109232 4324 109236 4380
rect 109236 4324 109292 4380
rect 109292 4324 109296 4380
rect 109232 4320 109296 4324
rect 109312 4380 109376 4384
rect 109312 4324 109316 4380
rect 109316 4324 109372 4380
rect 109372 4324 109376 4380
rect 109312 4320 109376 4324
rect 144832 4380 144896 4384
rect 144832 4324 144836 4380
rect 144836 4324 144892 4380
rect 144892 4324 144896 4380
rect 144832 4320 144896 4324
rect 144912 4380 144976 4384
rect 144912 4324 144916 4380
rect 144916 4324 144972 4380
rect 144972 4324 144976 4380
rect 144912 4320 144976 4324
rect 144992 4380 145056 4384
rect 144992 4324 144996 4380
rect 144996 4324 145052 4380
rect 145052 4324 145056 4380
rect 144992 4320 145056 4324
rect 145072 4380 145136 4384
rect 145072 4324 145076 4380
rect 145076 4324 145132 4380
rect 145132 4324 145136 4380
rect 145072 4320 145136 4324
rect 145152 4380 145216 4384
rect 145152 4324 145156 4380
rect 145156 4324 145212 4380
rect 145212 4324 145216 4380
rect 145152 4320 145216 4324
rect 145232 4380 145296 4384
rect 145232 4324 145236 4380
rect 145236 4324 145292 4380
rect 145292 4324 145296 4380
rect 145232 4320 145296 4324
rect 145312 4380 145376 4384
rect 145312 4324 145316 4380
rect 145316 4324 145372 4380
rect 145372 4324 145376 4380
rect 145312 4320 145376 4324
rect 180832 4380 180896 4384
rect 180832 4324 180836 4380
rect 180836 4324 180892 4380
rect 180892 4324 180896 4380
rect 180832 4320 180896 4324
rect 180912 4380 180976 4384
rect 180912 4324 180916 4380
rect 180916 4324 180972 4380
rect 180972 4324 180976 4380
rect 180912 4320 180976 4324
rect 180992 4380 181056 4384
rect 180992 4324 180996 4380
rect 180996 4324 181052 4380
rect 181052 4324 181056 4380
rect 180992 4320 181056 4324
rect 181072 4380 181136 4384
rect 181072 4324 181076 4380
rect 181076 4324 181132 4380
rect 181132 4324 181136 4380
rect 181072 4320 181136 4324
rect 181152 4380 181216 4384
rect 181152 4324 181156 4380
rect 181156 4324 181212 4380
rect 181212 4324 181216 4380
rect 181152 4320 181216 4324
rect 181232 4380 181296 4384
rect 181232 4324 181236 4380
rect 181236 4324 181292 4380
rect 181292 4324 181296 4380
rect 181232 4320 181296 4324
rect 181312 4380 181376 4384
rect 181312 4324 181316 4380
rect 181316 4324 181372 4380
rect 181372 4324 181376 4380
rect 181312 4320 181376 4324
rect 216832 4380 216896 4384
rect 216832 4324 216836 4380
rect 216836 4324 216892 4380
rect 216892 4324 216896 4380
rect 216832 4320 216896 4324
rect 216912 4380 216976 4384
rect 216912 4324 216916 4380
rect 216916 4324 216972 4380
rect 216972 4324 216976 4380
rect 216912 4320 216976 4324
rect 216992 4380 217056 4384
rect 216992 4324 216996 4380
rect 216996 4324 217052 4380
rect 217052 4324 217056 4380
rect 216992 4320 217056 4324
rect 217072 4380 217136 4384
rect 217072 4324 217076 4380
rect 217076 4324 217132 4380
rect 217132 4324 217136 4380
rect 217072 4320 217136 4324
rect 217152 4380 217216 4384
rect 217152 4324 217156 4380
rect 217156 4324 217212 4380
rect 217212 4324 217216 4380
rect 217152 4320 217216 4324
rect 217232 4380 217296 4384
rect 217232 4324 217236 4380
rect 217236 4324 217292 4380
rect 217292 4324 217296 4380
rect 217232 4320 217296 4324
rect 217312 4380 217376 4384
rect 217312 4324 217316 4380
rect 217316 4324 217372 4380
rect 217372 4324 217376 4380
rect 217312 4320 217376 4324
rect 252832 4380 252896 4384
rect 252832 4324 252836 4380
rect 252836 4324 252892 4380
rect 252892 4324 252896 4380
rect 252832 4320 252896 4324
rect 252912 4380 252976 4384
rect 252912 4324 252916 4380
rect 252916 4324 252972 4380
rect 252972 4324 252976 4380
rect 252912 4320 252976 4324
rect 252992 4380 253056 4384
rect 252992 4324 252996 4380
rect 252996 4324 253052 4380
rect 253052 4324 253056 4380
rect 252992 4320 253056 4324
rect 253072 4380 253136 4384
rect 253072 4324 253076 4380
rect 253076 4324 253132 4380
rect 253132 4324 253136 4380
rect 253072 4320 253136 4324
rect 253152 4380 253216 4384
rect 253152 4324 253156 4380
rect 253156 4324 253212 4380
rect 253212 4324 253216 4380
rect 253152 4320 253216 4324
rect 253232 4380 253296 4384
rect 253232 4324 253236 4380
rect 253236 4324 253292 4380
rect 253292 4324 253296 4380
rect 253232 4320 253296 4324
rect 253312 4380 253376 4384
rect 253312 4324 253316 4380
rect 253316 4324 253372 4380
rect 253372 4324 253376 4380
rect 253312 4320 253376 4324
rect 288832 4380 288896 4384
rect 288832 4324 288836 4380
rect 288836 4324 288892 4380
rect 288892 4324 288896 4380
rect 288832 4320 288896 4324
rect 288912 4380 288976 4384
rect 288912 4324 288916 4380
rect 288916 4324 288972 4380
rect 288972 4324 288976 4380
rect 288912 4320 288976 4324
rect 288992 4380 289056 4384
rect 288992 4324 288996 4380
rect 288996 4324 289052 4380
rect 289052 4324 289056 4380
rect 288992 4320 289056 4324
rect 289072 4380 289136 4384
rect 289072 4324 289076 4380
rect 289076 4324 289132 4380
rect 289132 4324 289136 4380
rect 289072 4320 289136 4324
rect 289152 4380 289216 4384
rect 289152 4324 289156 4380
rect 289156 4324 289212 4380
rect 289212 4324 289216 4380
rect 289152 4320 289216 4324
rect 289232 4380 289296 4384
rect 289232 4324 289236 4380
rect 289236 4324 289292 4380
rect 289292 4324 289296 4380
rect 289232 4320 289296 4324
rect 289312 4380 289376 4384
rect 289312 4324 289316 4380
rect 289316 4324 289372 4380
rect 289372 4324 289376 4380
rect 289312 4320 289376 4324
rect 324832 4380 324896 4384
rect 324832 4324 324836 4380
rect 324836 4324 324892 4380
rect 324892 4324 324896 4380
rect 324832 4320 324896 4324
rect 324912 4380 324976 4384
rect 324912 4324 324916 4380
rect 324916 4324 324972 4380
rect 324972 4324 324976 4380
rect 324912 4320 324976 4324
rect 324992 4380 325056 4384
rect 324992 4324 324996 4380
rect 324996 4324 325052 4380
rect 325052 4324 325056 4380
rect 324992 4320 325056 4324
rect 325072 4380 325136 4384
rect 325072 4324 325076 4380
rect 325076 4324 325132 4380
rect 325132 4324 325136 4380
rect 325072 4320 325136 4324
rect 325152 4380 325216 4384
rect 325152 4324 325156 4380
rect 325156 4324 325212 4380
rect 325212 4324 325216 4380
rect 325152 4320 325216 4324
rect 325232 4380 325296 4384
rect 325232 4324 325236 4380
rect 325236 4324 325292 4380
rect 325292 4324 325296 4380
rect 325232 4320 325296 4324
rect 325312 4380 325376 4384
rect 325312 4324 325316 4380
rect 325316 4324 325372 4380
rect 325372 4324 325376 4380
rect 325312 4320 325376 4324
rect 360832 4380 360896 4384
rect 360832 4324 360836 4380
rect 360836 4324 360892 4380
rect 360892 4324 360896 4380
rect 360832 4320 360896 4324
rect 360912 4380 360976 4384
rect 360912 4324 360916 4380
rect 360916 4324 360972 4380
rect 360972 4324 360976 4380
rect 360912 4320 360976 4324
rect 360992 4380 361056 4384
rect 360992 4324 360996 4380
rect 360996 4324 361052 4380
rect 361052 4324 361056 4380
rect 360992 4320 361056 4324
rect 361072 4380 361136 4384
rect 361072 4324 361076 4380
rect 361076 4324 361132 4380
rect 361132 4324 361136 4380
rect 361072 4320 361136 4324
rect 361152 4380 361216 4384
rect 361152 4324 361156 4380
rect 361156 4324 361212 4380
rect 361212 4324 361216 4380
rect 361152 4320 361216 4324
rect 361232 4380 361296 4384
rect 361232 4324 361236 4380
rect 361236 4324 361292 4380
rect 361292 4324 361296 4380
rect 361232 4320 361296 4324
rect 361312 4380 361376 4384
rect 361312 4324 361316 4380
rect 361316 4324 361372 4380
rect 361372 4324 361376 4380
rect 361312 4320 361376 4324
rect 396832 4380 396896 4384
rect 396832 4324 396836 4380
rect 396836 4324 396892 4380
rect 396892 4324 396896 4380
rect 396832 4320 396896 4324
rect 396912 4380 396976 4384
rect 396912 4324 396916 4380
rect 396916 4324 396972 4380
rect 396972 4324 396976 4380
rect 396912 4320 396976 4324
rect 396992 4380 397056 4384
rect 396992 4324 396996 4380
rect 396996 4324 397052 4380
rect 397052 4324 397056 4380
rect 396992 4320 397056 4324
rect 397072 4380 397136 4384
rect 397072 4324 397076 4380
rect 397076 4324 397132 4380
rect 397132 4324 397136 4380
rect 397072 4320 397136 4324
rect 397152 4380 397216 4384
rect 397152 4324 397156 4380
rect 397156 4324 397212 4380
rect 397212 4324 397216 4380
rect 397152 4320 397216 4324
rect 397232 4380 397296 4384
rect 397232 4324 397236 4380
rect 397236 4324 397292 4380
rect 397292 4324 397296 4380
rect 397232 4320 397296 4324
rect 397312 4380 397376 4384
rect 397312 4324 397316 4380
rect 397316 4324 397372 4380
rect 397372 4324 397376 4380
rect 397312 4320 397376 4324
rect 432832 4380 432896 4384
rect 432832 4324 432836 4380
rect 432836 4324 432892 4380
rect 432892 4324 432896 4380
rect 432832 4320 432896 4324
rect 432912 4380 432976 4384
rect 432912 4324 432916 4380
rect 432916 4324 432972 4380
rect 432972 4324 432976 4380
rect 432912 4320 432976 4324
rect 432992 4380 433056 4384
rect 432992 4324 432996 4380
rect 432996 4324 433052 4380
rect 433052 4324 433056 4380
rect 432992 4320 433056 4324
rect 433072 4380 433136 4384
rect 433072 4324 433076 4380
rect 433076 4324 433132 4380
rect 433132 4324 433136 4380
rect 433072 4320 433136 4324
rect 433152 4380 433216 4384
rect 433152 4324 433156 4380
rect 433156 4324 433212 4380
rect 433212 4324 433216 4380
rect 433152 4320 433216 4324
rect 433232 4380 433296 4384
rect 433232 4324 433236 4380
rect 433236 4324 433292 4380
rect 433292 4324 433296 4380
rect 433232 4320 433296 4324
rect 433312 4380 433376 4384
rect 433312 4324 433316 4380
rect 433316 4324 433372 4380
rect 433372 4324 433376 4380
rect 433312 4320 433376 4324
rect 468832 4380 468896 4384
rect 468832 4324 468836 4380
rect 468836 4324 468892 4380
rect 468892 4324 468896 4380
rect 468832 4320 468896 4324
rect 468912 4380 468976 4384
rect 468912 4324 468916 4380
rect 468916 4324 468972 4380
rect 468972 4324 468976 4380
rect 468912 4320 468976 4324
rect 468992 4380 469056 4384
rect 468992 4324 468996 4380
rect 468996 4324 469052 4380
rect 469052 4324 469056 4380
rect 468992 4320 469056 4324
rect 469072 4380 469136 4384
rect 469072 4324 469076 4380
rect 469076 4324 469132 4380
rect 469132 4324 469136 4380
rect 469072 4320 469136 4324
rect 469152 4380 469216 4384
rect 469152 4324 469156 4380
rect 469156 4324 469212 4380
rect 469212 4324 469216 4380
rect 469152 4320 469216 4324
rect 469232 4380 469296 4384
rect 469232 4324 469236 4380
rect 469236 4324 469292 4380
rect 469292 4324 469296 4380
rect 469232 4320 469296 4324
rect 469312 4380 469376 4384
rect 469312 4324 469316 4380
rect 469316 4324 469372 4380
rect 469372 4324 469376 4380
rect 469312 4320 469376 4324
rect 504832 4380 504896 4384
rect 504832 4324 504836 4380
rect 504836 4324 504892 4380
rect 504892 4324 504896 4380
rect 504832 4320 504896 4324
rect 504912 4380 504976 4384
rect 504912 4324 504916 4380
rect 504916 4324 504972 4380
rect 504972 4324 504976 4380
rect 504912 4320 504976 4324
rect 504992 4380 505056 4384
rect 504992 4324 504996 4380
rect 504996 4324 505052 4380
rect 505052 4324 505056 4380
rect 504992 4320 505056 4324
rect 505072 4380 505136 4384
rect 505072 4324 505076 4380
rect 505076 4324 505132 4380
rect 505132 4324 505136 4380
rect 505072 4320 505136 4324
rect 505152 4380 505216 4384
rect 505152 4324 505156 4380
rect 505156 4324 505212 4380
rect 505212 4324 505216 4380
rect 505152 4320 505216 4324
rect 505232 4380 505296 4384
rect 505232 4324 505236 4380
rect 505236 4324 505292 4380
rect 505292 4324 505296 4380
rect 505232 4320 505296 4324
rect 505312 4380 505376 4384
rect 505312 4324 505316 4380
rect 505316 4324 505372 4380
rect 505372 4324 505376 4380
rect 505312 4320 505376 4324
rect 540832 4380 540896 4384
rect 540832 4324 540836 4380
rect 540836 4324 540892 4380
rect 540892 4324 540896 4380
rect 540832 4320 540896 4324
rect 540912 4380 540976 4384
rect 540912 4324 540916 4380
rect 540916 4324 540972 4380
rect 540972 4324 540976 4380
rect 540912 4320 540976 4324
rect 540992 4380 541056 4384
rect 540992 4324 540996 4380
rect 540996 4324 541052 4380
rect 541052 4324 541056 4380
rect 540992 4320 541056 4324
rect 541072 4380 541136 4384
rect 541072 4324 541076 4380
rect 541076 4324 541132 4380
rect 541132 4324 541136 4380
rect 541072 4320 541136 4324
rect 541152 4380 541216 4384
rect 541152 4324 541156 4380
rect 541156 4324 541212 4380
rect 541212 4324 541216 4380
rect 541152 4320 541216 4324
rect 541232 4380 541296 4384
rect 541232 4324 541236 4380
rect 541236 4324 541292 4380
rect 541292 4324 541296 4380
rect 541232 4320 541296 4324
rect 541312 4380 541376 4384
rect 541312 4324 541316 4380
rect 541316 4324 541372 4380
rect 541372 4324 541376 4380
rect 541312 4320 541376 4324
rect 576832 4380 576896 4384
rect 576832 4324 576836 4380
rect 576836 4324 576892 4380
rect 576892 4324 576896 4380
rect 576832 4320 576896 4324
rect 576912 4380 576976 4384
rect 576912 4324 576916 4380
rect 576916 4324 576972 4380
rect 576972 4324 576976 4380
rect 576912 4320 576976 4324
rect 576992 4380 577056 4384
rect 576992 4324 576996 4380
rect 576996 4324 577052 4380
rect 577052 4324 577056 4380
rect 576992 4320 577056 4324
rect 577072 4380 577136 4384
rect 577072 4324 577076 4380
rect 577076 4324 577132 4380
rect 577132 4324 577136 4380
rect 577072 4320 577136 4324
rect 577152 4380 577216 4384
rect 577152 4324 577156 4380
rect 577156 4324 577212 4380
rect 577212 4324 577216 4380
rect 577152 4320 577216 4324
rect 577232 4380 577296 4384
rect 577232 4324 577236 4380
rect 577236 4324 577292 4380
rect 577292 4324 577296 4380
rect 577232 4320 577296 4324
rect 577312 4380 577376 4384
rect 577312 4324 577316 4380
rect 577316 4324 577372 4380
rect 577372 4324 577376 4380
rect 577312 4320 577376 4324
rect 18832 3836 18896 3840
rect 18832 3780 18836 3836
rect 18836 3780 18892 3836
rect 18892 3780 18896 3836
rect 18832 3776 18896 3780
rect 18912 3836 18976 3840
rect 18912 3780 18916 3836
rect 18916 3780 18972 3836
rect 18972 3780 18976 3836
rect 18912 3776 18976 3780
rect 18992 3836 19056 3840
rect 18992 3780 18996 3836
rect 18996 3780 19052 3836
rect 19052 3780 19056 3836
rect 18992 3776 19056 3780
rect 19072 3836 19136 3840
rect 19072 3780 19076 3836
rect 19076 3780 19132 3836
rect 19132 3780 19136 3836
rect 19072 3776 19136 3780
rect 19152 3836 19216 3840
rect 19152 3780 19156 3836
rect 19156 3780 19212 3836
rect 19212 3780 19216 3836
rect 19152 3776 19216 3780
rect 19232 3836 19296 3840
rect 19232 3780 19236 3836
rect 19236 3780 19292 3836
rect 19292 3780 19296 3836
rect 19232 3776 19296 3780
rect 19312 3836 19376 3840
rect 19312 3780 19316 3836
rect 19316 3780 19372 3836
rect 19372 3780 19376 3836
rect 19312 3776 19376 3780
rect 54832 3836 54896 3840
rect 54832 3780 54836 3836
rect 54836 3780 54892 3836
rect 54892 3780 54896 3836
rect 54832 3776 54896 3780
rect 54912 3836 54976 3840
rect 54912 3780 54916 3836
rect 54916 3780 54972 3836
rect 54972 3780 54976 3836
rect 54912 3776 54976 3780
rect 54992 3836 55056 3840
rect 54992 3780 54996 3836
rect 54996 3780 55052 3836
rect 55052 3780 55056 3836
rect 54992 3776 55056 3780
rect 55072 3836 55136 3840
rect 55072 3780 55076 3836
rect 55076 3780 55132 3836
rect 55132 3780 55136 3836
rect 55072 3776 55136 3780
rect 55152 3836 55216 3840
rect 55152 3780 55156 3836
rect 55156 3780 55212 3836
rect 55212 3780 55216 3836
rect 55152 3776 55216 3780
rect 55232 3836 55296 3840
rect 55232 3780 55236 3836
rect 55236 3780 55292 3836
rect 55292 3780 55296 3836
rect 55232 3776 55296 3780
rect 55312 3836 55376 3840
rect 55312 3780 55316 3836
rect 55316 3780 55372 3836
rect 55372 3780 55376 3836
rect 55312 3776 55376 3780
rect 90832 3836 90896 3840
rect 90832 3780 90836 3836
rect 90836 3780 90892 3836
rect 90892 3780 90896 3836
rect 90832 3776 90896 3780
rect 90912 3836 90976 3840
rect 90912 3780 90916 3836
rect 90916 3780 90972 3836
rect 90972 3780 90976 3836
rect 90912 3776 90976 3780
rect 90992 3836 91056 3840
rect 90992 3780 90996 3836
rect 90996 3780 91052 3836
rect 91052 3780 91056 3836
rect 90992 3776 91056 3780
rect 91072 3836 91136 3840
rect 91072 3780 91076 3836
rect 91076 3780 91132 3836
rect 91132 3780 91136 3836
rect 91072 3776 91136 3780
rect 91152 3836 91216 3840
rect 91152 3780 91156 3836
rect 91156 3780 91212 3836
rect 91212 3780 91216 3836
rect 91152 3776 91216 3780
rect 91232 3836 91296 3840
rect 91232 3780 91236 3836
rect 91236 3780 91292 3836
rect 91292 3780 91296 3836
rect 91232 3776 91296 3780
rect 91312 3836 91376 3840
rect 91312 3780 91316 3836
rect 91316 3780 91372 3836
rect 91372 3780 91376 3836
rect 91312 3776 91376 3780
rect 126832 3836 126896 3840
rect 126832 3780 126836 3836
rect 126836 3780 126892 3836
rect 126892 3780 126896 3836
rect 126832 3776 126896 3780
rect 126912 3836 126976 3840
rect 126912 3780 126916 3836
rect 126916 3780 126972 3836
rect 126972 3780 126976 3836
rect 126912 3776 126976 3780
rect 126992 3836 127056 3840
rect 126992 3780 126996 3836
rect 126996 3780 127052 3836
rect 127052 3780 127056 3836
rect 126992 3776 127056 3780
rect 127072 3836 127136 3840
rect 127072 3780 127076 3836
rect 127076 3780 127132 3836
rect 127132 3780 127136 3836
rect 127072 3776 127136 3780
rect 127152 3836 127216 3840
rect 127152 3780 127156 3836
rect 127156 3780 127212 3836
rect 127212 3780 127216 3836
rect 127152 3776 127216 3780
rect 127232 3836 127296 3840
rect 127232 3780 127236 3836
rect 127236 3780 127292 3836
rect 127292 3780 127296 3836
rect 127232 3776 127296 3780
rect 127312 3836 127376 3840
rect 127312 3780 127316 3836
rect 127316 3780 127372 3836
rect 127372 3780 127376 3836
rect 127312 3776 127376 3780
rect 162832 3836 162896 3840
rect 162832 3780 162836 3836
rect 162836 3780 162892 3836
rect 162892 3780 162896 3836
rect 162832 3776 162896 3780
rect 162912 3836 162976 3840
rect 162912 3780 162916 3836
rect 162916 3780 162972 3836
rect 162972 3780 162976 3836
rect 162912 3776 162976 3780
rect 162992 3836 163056 3840
rect 162992 3780 162996 3836
rect 162996 3780 163052 3836
rect 163052 3780 163056 3836
rect 162992 3776 163056 3780
rect 163072 3836 163136 3840
rect 163072 3780 163076 3836
rect 163076 3780 163132 3836
rect 163132 3780 163136 3836
rect 163072 3776 163136 3780
rect 163152 3836 163216 3840
rect 163152 3780 163156 3836
rect 163156 3780 163212 3836
rect 163212 3780 163216 3836
rect 163152 3776 163216 3780
rect 163232 3836 163296 3840
rect 163232 3780 163236 3836
rect 163236 3780 163292 3836
rect 163292 3780 163296 3836
rect 163232 3776 163296 3780
rect 163312 3836 163376 3840
rect 163312 3780 163316 3836
rect 163316 3780 163372 3836
rect 163372 3780 163376 3836
rect 163312 3776 163376 3780
rect 198832 3836 198896 3840
rect 198832 3780 198836 3836
rect 198836 3780 198892 3836
rect 198892 3780 198896 3836
rect 198832 3776 198896 3780
rect 198912 3836 198976 3840
rect 198912 3780 198916 3836
rect 198916 3780 198972 3836
rect 198972 3780 198976 3836
rect 198912 3776 198976 3780
rect 198992 3836 199056 3840
rect 198992 3780 198996 3836
rect 198996 3780 199052 3836
rect 199052 3780 199056 3836
rect 198992 3776 199056 3780
rect 199072 3836 199136 3840
rect 199072 3780 199076 3836
rect 199076 3780 199132 3836
rect 199132 3780 199136 3836
rect 199072 3776 199136 3780
rect 199152 3836 199216 3840
rect 199152 3780 199156 3836
rect 199156 3780 199212 3836
rect 199212 3780 199216 3836
rect 199152 3776 199216 3780
rect 199232 3836 199296 3840
rect 199232 3780 199236 3836
rect 199236 3780 199292 3836
rect 199292 3780 199296 3836
rect 199232 3776 199296 3780
rect 199312 3836 199376 3840
rect 199312 3780 199316 3836
rect 199316 3780 199372 3836
rect 199372 3780 199376 3836
rect 199312 3776 199376 3780
rect 234832 3836 234896 3840
rect 234832 3780 234836 3836
rect 234836 3780 234892 3836
rect 234892 3780 234896 3836
rect 234832 3776 234896 3780
rect 234912 3836 234976 3840
rect 234912 3780 234916 3836
rect 234916 3780 234972 3836
rect 234972 3780 234976 3836
rect 234912 3776 234976 3780
rect 234992 3836 235056 3840
rect 234992 3780 234996 3836
rect 234996 3780 235052 3836
rect 235052 3780 235056 3836
rect 234992 3776 235056 3780
rect 235072 3836 235136 3840
rect 235072 3780 235076 3836
rect 235076 3780 235132 3836
rect 235132 3780 235136 3836
rect 235072 3776 235136 3780
rect 235152 3836 235216 3840
rect 235152 3780 235156 3836
rect 235156 3780 235212 3836
rect 235212 3780 235216 3836
rect 235152 3776 235216 3780
rect 235232 3836 235296 3840
rect 235232 3780 235236 3836
rect 235236 3780 235292 3836
rect 235292 3780 235296 3836
rect 235232 3776 235296 3780
rect 235312 3836 235376 3840
rect 235312 3780 235316 3836
rect 235316 3780 235372 3836
rect 235372 3780 235376 3836
rect 235312 3776 235376 3780
rect 270832 3836 270896 3840
rect 270832 3780 270836 3836
rect 270836 3780 270892 3836
rect 270892 3780 270896 3836
rect 270832 3776 270896 3780
rect 270912 3836 270976 3840
rect 270912 3780 270916 3836
rect 270916 3780 270972 3836
rect 270972 3780 270976 3836
rect 270912 3776 270976 3780
rect 270992 3836 271056 3840
rect 270992 3780 270996 3836
rect 270996 3780 271052 3836
rect 271052 3780 271056 3836
rect 270992 3776 271056 3780
rect 271072 3836 271136 3840
rect 271072 3780 271076 3836
rect 271076 3780 271132 3836
rect 271132 3780 271136 3836
rect 271072 3776 271136 3780
rect 271152 3836 271216 3840
rect 271152 3780 271156 3836
rect 271156 3780 271212 3836
rect 271212 3780 271216 3836
rect 271152 3776 271216 3780
rect 271232 3836 271296 3840
rect 271232 3780 271236 3836
rect 271236 3780 271292 3836
rect 271292 3780 271296 3836
rect 271232 3776 271296 3780
rect 271312 3836 271376 3840
rect 271312 3780 271316 3836
rect 271316 3780 271372 3836
rect 271372 3780 271376 3836
rect 271312 3776 271376 3780
rect 306832 3836 306896 3840
rect 306832 3780 306836 3836
rect 306836 3780 306892 3836
rect 306892 3780 306896 3836
rect 306832 3776 306896 3780
rect 306912 3836 306976 3840
rect 306912 3780 306916 3836
rect 306916 3780 306972 3836
rect 306972 3780 306976 3836
rect 306912 3776 306976 3780
rect 306992 3836 307056 3840
rect 306992 3780 306996 3836
rect 306996 3780 307052 3836
rect 307052 3780 307056 3836
rect 306992 3776 307056 3780
rect 307072 3836 307136 3840
rect 307072 3780 307076 3836
rect 307076 3780 307132 3836
rect 307132 3780 307136 3836
rect 307072 3776 307136 3780
rect 307152 3836 307216 3840
rect 307152 3780 307156 3836
rect 307156 3780 307212 3836
rect 307212 3780 307216 3836
rect 307152 3776 307216 3780
rect 307232 3836 307296 3840
rect 307232 3780 307236 3836
rect 307236 3780 307292 3836
rect 307292 3780 307296 3836
rect 307232 3776 307296 3780
rect 307312 3836 307376 3840
rect 307312 3780 307316 3836
rect 307316 3780 307372 3836
rect 307372 3780 307376 3836
rect 307312 3776 307376 3780
rect 342832 3836 342896 3840
rect 342832 3780 342836 3836
rect 342836 3780 342892 3836
rect 342892 3780 342896 3836
rect 342832 3776 342896 3780
rect 342912 3836 342976 3840
rect 342912 3780 342916 3836
rect 342916 3780 342972 3836
rect 342972 3780 342976 3836
rect 342912 3776 342976 3780
rect 342992 3836 343056 3840
rect 342992 3780 342996 3836
rect 342996 3780 343052 3836
rect 343052 3780 343056 3836
rect 342992 3776 343056 3780
rect 343072 3836 343136 3840
rect 343072 3780 343076 3836
rect 343076 3780 343132 3836
rect 343132 3780 343136 3836
rect 343072 3776 343136 3780
rect 343152 3836 343216 3840
rect 343152 3780 343156 3836
rect 343156 3780 343212 3836
rect 343212 3780 343216 3836
rect 343152 3776 343216 3780
rect 343232 3836 343296 3840
rect 343232 3780 343236 3836
rect 343236 3780 343292 3836
rect 343292 3780 343296 3836
rect 343232 3776 343296 3780
rect 343312 3836 343376 3840
rect 343312 3780 343316 3836
rect 343316 3780 343372 3836
rect 343372 3780 343376 3836
rect 343312 3776 343376 3780
rect 378832 3836 378896 3840
rect 378832 3780 378836 3836
rect 378836 3780 378892 3836
rect 378892 3780 378896 3836
rect 378832 3776 378896 3780
rect 378912 3836 378976 3840
rect 378912 3780 378916 3836
rect 378916 3780 378972 3836
rect 378972 3780 378976 3836
rect 378912 3776 378976 3780
rect 378992 3836 379056 3840
rect 378992 3780 378996 3836
rect 378996 3780 379052 3836
rect 379052 3780 379056 3836
rect 378992 3776 379056 3780
rect 379072 3836 379136 3840
rect 379072 3780 379076 3836
rect 379076 3780 379132 3836
rect 379132 3780 379136 3836
rect 379072 3776 379136 3780
rect 379152 3836 379216 3840
rect 379152 3780 379156 3836
rect 379156 3780 379212 3836
rect 379212 3780 379216 3836
rect 379152 3776 379216 3780
rect 379232 3836 379296 3840
rect 379232 3780 379236 3836
rect 379236 3780 379292 3836
rect 379292 3780 379296 3836
rect 379232 3776 379296 3780
rect 379312 3836 379376 3840
rect 379312 3780 379316 3836
rect 379316 3780 379372 3836
rect 379372 3780 379376 3836
rect 379312 3776 379376 3780
rect 414832 3836 414896 3840
rect 414832 3780 414836 3836
rect 414836 3780 414892 3836
rect 414892 3780 414896 3836
rect 414832 3776 414896 3780
rect 414912 3836 414976 3840
rect 414912 3780 414916 3836
rect 414916 3780 414972 3836
rect 414972 3780 414976 3836
rect 414912 3776 414976 3780
rect 414992 3836 415056 3840
rect 414992 3780 414996 3836
rect 414996 3780 415052 3836
rect 415052 3780 415056 3836
rect 414992 3776 415056 3780
rect 415072 3836 415136 3840
rect 415072 3780 415076 3836
rect 415076 3780 415132 3836
rect 415132 3780 415136 3836
rect 415072 3776 415136 3780
rect 415152 3836 415216 3840
rect 415152 3780 415156 3836
rect 415156 3780 415212 3836
rect 415212 3780 415216 3836
rect 415152 3776 415216 3780
rect 415232 3836 415296 3840
rect 415232 3780 415236 3836
rect 415236 3780 415292 3836
rect 415292 3780 415296 3836
rect 415232 3776 415296 3780
rect 415312 3836 415376 3840
rect 415312 3780 415316 3836
rect 415316 3780 415372 3836
rect 415372 3780 415376 3836
rect 415312 3776 415376 3780
rect 450832 3836 450896 3840
rect 450832 3780 450836 3836
rect 450836 3780 450892 3836
rect 450892 3780 450896 3836
rect 450832 3776 450896 3780
rect 450912 3836 450976 3840
rect 450912 3780 450916 3836
rect 450916 3780 450972 3836
rect 450972 3780 450976 3836
rect 450912 3776 450976 3780
rect 450992 3836 451056 3840
rect 450992 3780 450996 3836
rect 450996 3780 451052 3836
rect 451052 3780 451056 3836
rect 450992 3776 451056 3780
rect 451072 3836 451136 3840
rect 451072 3780 451076 3836
rect 451076 3780 451132 3836
rect 451132 3780 451136 3836
rect 451072 3776 451136 3780
rect 451152 3836 451216 3840
rect 451152 3780 451156 3836
rect 451156 3780 451212 3836
rect 451212 3780 451216 3836
rect 451152 3776 451216 3780
rect 451232 3836 451296 3840
rect 451232 3780 451236 3836
rect 451236 3780 451292 3836
rect 451292 3780 451296 3836
rect 451232 3776 451296 3780
rect 451312 3836 451376 3840
rect 451312 3780 451316 3836
rect 451316 3780 451372 3836
rect 451372 3780 451376 3836
rect 451312 3776 451376 3780
rect 486832 3836 486896 3840
rect 486832 3780 486836 3836
rect 486836 3780 486892 3836
rect 486892 3780 486896 3836
rect 486832 3776 486896 3780
rect 486912 3836 486976 3840
rect 486912 3780 486916 3836
rect 486916 3780 486972 3836
rect 486972 3780 486976 3836
rect 486912 3776 486976 3780
rect 486992 3836 487056 3840
rect 486992 3780 486996 3836
rect 486996 3780 487052 3836
rect 487052 3780 487056 3836
rect 486992 3776 487056 3780
rect 487072 3836 487136 3840
rect 487072 3780 487076 3836
rect 487076 3780 487132 3836
rect 487132 3780 487136 3836
rect 487072 3776 487136 3780
rect 487152 3836 487216 3840
rect 487152 3780 487156 3836
rect 487156 3780 487212 3836
rect 487212 3780 487216 3836
rect 487152 3776 487216 3780
rect 487232 3836 487296 3840
rect 487232 3780 487236 3836
rect 487236 3780 487292 3836
rect 487292 3780 487296 3836
rect 487232 3776 487296 3780
rect 487312 3836 487376 3840
rect 487312 3780 487316 3836
rect 487316 3780 487372 3836
rect 487372 3780 487376 3836
rect 487312 3776 487376 3780
rect 522832 3836 522896 3840
rect 522832 3780 522836 3836
rect 522836 3780 522892 3836
rect 522892 3780 522896 3836
rect 522832 3776 522896 3780
rect 522912 3836 522976 3840
rect 522912 3780 522916 3836
rect 522916 3780 522972 3836
rect 522972 3780 522976 3836
rect 522912 3776 522976 3780
rect 522992 3836 523056 3840
rect 522992 3780 522996 3836
rect 522996 3780 523052 3836
rect 523052 3780 523056 3836
rect 522992 3776 523056 3780
rect 523072 3836 523136 3840
rect 523072 3780 523076 3836
rect 523076 3780 523132 3836
rect 523132 3780 523136 3836
rect 523072 3776 523136 3780
rect 523152 3836 523216 3840
rect 523152 3780 523156 3836
rect 523156 3780 523212 3836
rect 523212 3780 523216 3836
rect 523152 3776 523216 3780
rect 523232 3836 523296 3840
rect 523232 3780 523236 3836
rect 523236 3780 523292 3836
rect 523292 3780 523296 3836
rect 523232 3776 523296 3780
rect 523312 3836 523376 3840
rect 523312 3780 523316 3836
rect 523316 3780 523372 3836
rect 523372 3780 523376 3836
rect 523312 3776 523376 3780
rect 558832 3836 558896 3840
rect 558832 3780 558836 3836
rect 558836 3780 558892 3836
rect 558892 3780 558896 3836
rect 558832 3776 558896 3780
rect 558912 3836 558976 3840
rect 558912 3780 558916 3836
rect 558916 3780 558972 3836
rect 558972 3780 558976 3836
rect 558912 3776 558976 3780
rect 558992 3836 559056 3840
rect 558992 3780 558996 3836
rect 558996 3780 559052 3836
rect 559052 3780 559056 3836
rect 558992 3776 559056 3780
rect 559072 3836 559136 3840
rect 559072 3780 559076 3836
rect 559076 3780 559132 3836
rect 559132 3780 559136 3836
rect 559072 3776 559136 3780
rect 559152 3836 559216 3840
rect 559152 3780 559156 3836
rect 559156 3780 559212 3836
rect 559212 3780 559216 3836
rect 559152 3776 559216 3780
rect 559232 3836 559296 3840
rect 559232 3780 559236 3836
rect 559236 3780 559292 3836
rect 559292 3780 559296 3836
rect 559232 3776 559296 3780
rect 559312 3836 559376 3840
rect 559312 3780 559316 3836
rect 559316 3780 559372 3836
rect 559372 3780 559376 3836
rect 559312 3776 559376 3780
rect 36832 3292 36896 3296
rect 36832 3236 36836 3292
rect 36836 3236 36892 3292
rect 36892 3236 36896 3292
rect 36832 3232 36896 3236
rect 36912 3292 36976 3296
rect 36912 3236 36916 3292
rect 36916 3236 36972 3292
rect 36972 3236 36976 3292
rect 36912 3232 36976 3236
rect 36992 3292 37056 3296
rect 36992 3236 36996 3292
rect 36996 3236 37052 3292
rect 37052 3236 37056 3292
rect 36992 3232 37056 3236
rect 37072 3292 37136 3296
rect 37072 3236 37076 3292
rect 37076 3236 37132 3292
rect 37132 3236 37136 3292
rect 37072 3232 37136 3236
rect 37152 3292 37216 3296
rect 37152 3236 37156 3292
rect 37156 3236 37212 3292
rect 37212 3236 37216 3292
rect 37152 3232 37216 3236
rect 37232 3292 37296 3296
rect 37232 3236 37236 3292
rect 37236 3236 37292 3292
rect 37292 3236 37296 3292
rect 37232 3232 37296 3236
rect 37312 3292 37376 3296
rect 37312 3236 37316 3292
rect 37316 3236 37372 3292
rect 37372 3236 37376 3292
rect 37312 3232 37376 3236
rect 72832 3292 72896 3296
rect 72832 3236 72836 3292
rect 72836 3236 72892 3292
rect 72892 3236 72896 3292
rect 72832 3232 72896 3236
rect 72912 3292 72976 3296
rect 72912 3236 72916 3292
rect 72916 3236 72972 3292
rect 72972 3236 72976 3292
rect 72912 3232 72976 3236
rect 72992 3292 73056 3296
rect 72992 3236 72996 3292
rect 72996 3236 73052 3292
rect 73052 3236 73056 3292
rect 72992 3232 73056 3236
rect 73072 3292 73136 3296
rect 73072 3236 73076 3292
rect 73076 3236 73132 3292
rect 73132 3236 73136 3292
rect 73072 3232 73136 3236
rect 73152 3292 73216 3296
rect 73152 3236 73156 3292
rect 73156 3236 73212 3292
rect 73212 3236 73216 3292
rect 73152 3232 73216 3236
rect 73232 3292 73296 3296
rect 73232 3236 73236 3292
rect 73236 3236 73292 3292
rect 73292 3236 73296 3292
rect 73232 3232 73296 3236
rect 73312 3292 73376 3296
rect 73312 3236 73316 3292
rect 73316 3236 73372 3292
rect 73372 3236 73376 3292
rect 73312 3232 73376 3236
rect 108832 3292 108896 3296
rect 108832 3236 108836 3292
rect 108836 3236 108892 3292
rect 108892 3236 108896 3292
rect 108832 3232 108896 3236
rect 108912 3292 108976 3296
rect 108912 3236 108916 3292
rect 108916 3236 108972 3292
rect 108972 3236 108976 3292
rect 108912 3232 108976 3236
rect 108992 3292 109056 3296
rect 108992 3236 108996 3292
rect 108996 3236 109052 3292
rect 109052 3236 109056 3292
rect 108992 3232 109056 3236
rect 109072 3292 109136 3296
rect 109072 3236 109076 3292
rect 109076 3236 109132 3292
rect 109132 3236 109136 3292
rect 109072 3232 109136 3236
rect 109152 3292 109216 3296
rect 109152 3236 109156 3292
rect 109156 3236 109212 3292
rect 109212 3236 109216 3292
rect 109152 3232 109216 3236
rect 109232 3292 109296 3296
rect 109232 3236 109236 3292
rect 109236 3236 109292 3292
rect 109292 3236 109296 3292
rect 109232 3232 109296 3236
rect 109312 3292 109376 3296
rect 109312 3236 109316 3292
rect 109316 3236 109372 3292
rect 109372 3236 109376 3292
rect 109312 3232 109376 3236
rect 144832 3292 144896 3296
rect 144832 3236 144836 3292
rect 144836 3236 144892 3292
rect 144892 3236 144896 3292
rect 144832 3232 144896 3236
rect 144912 3292 144976 3296
rect 144912 3236 144916 3292
rect 144916 3236 144972 3292
rect 144972 3236 144976 3292
rect 144912 3232 144976 3236
rect 144992 3292 145056 3296
rect 144992 3236 144996 3292
rect 144996 3236 145052 3292
rect 145052 3236 145056 3292
rect 144992 3232 145056 3236
rect 145072 3292 145136 3296
rect 145072 3236 145076 3292
rect 145076 3236 145132 3292
rect 145132 3236 145136 3292
rect 145072 3232 145136 3236
rect 145152 3292 145216 3296
rect 145152 3236 145156 3292
rect 145156 3236 145212 3292
rect 145212 3236 145216 3292
rect 145152 3232 145216 3236
rect 145232 3292 145296 3296
rect 145232 3236 145236 3292
rect 145236 3236 145292 3292
rect 145292 3236 145296 3292
rect 145232 3232 145296 3236
rect 145312 3292 145376 3296
rect 145312 3236 145316 3292
rect 145316 3236 145372 3292
rect 145372 3236 145376 3292
rect 145312 3232 145376 3236
rect 180832 3292 180896 3296
rect 180832 3236 180836 3292
rect 180836 3236 180892 3292
rect 180892 3236 180896 3292
rect 180832 3232 180896 3236
rect 180912 3292 180976 3296
rect 180912 3236 180916 3292
rect 180916 3236 180972 3292
rect 180972 3236 180976 3292
rect 180912 3232 180976 3236
rect 180992 3292 181056 3296
rect 180992 3236 180996 3292
rect 180996 3236 181052 3292
rect 181052 3236 181056 3292
rect 180992 3232 181056 3236
rect 181072 3292 181136 3296
rect 181072 3236 181076 3292
rect 181076 3236 181132 3292
rect 181132 3236 181136 3292
rect 181072 3232 181136 3236
rect 181152 3292 181216 3296
rect 181152 3236 181156 3292
rect 181156 3236 181212 3292
rect 181212 3236 181216 3292
rect 181152 3232 181216 3236
rect 181232 3292 181296 3296
rect 181232 3236 181236 3292
rect 181236 3236 181292 3292
rect 181292 3236 181296 3292
rect 181232 3232 181296 3236
rect 181312 3292 181376 3296
rect 181312 3236 181316 3292
rect 181316 3236 181372 3292
rect 181372 3236 181376 3292
rect 181312 3232 181376 3236
rect 216832 3292 216896 3296
rect 216832 3236 216836 3292
rect 216836 3236 216892 3292
rect 216892 3236 216896 3292
rect 216832 3232 216896 3236
rect 216912 3292 216976 3296
rect 216912 3236 216916 3292
rect 216916 3236 216972 3292
rect 216972 3236 216976 3292
rect 216912 3232 216976 3236
rect 216992 3292 217056 3296
rect 216992 3236 216996 3292
rect 216996 3236 217052 3292
rect 217052 3236 217056 3292
rect 216992 3232 217056 3236
rect 217072 3292 217136 3296
rect 217072 3236 217076 3292
rect 217076 3236 217132 3292
rect 217132 3236 217136 3292
rect 217072 3232 217136 3236
rect 217152 3292 217216 3296
rect 217152 3236 217156 3292
rect 217156 3236 217212 3292
rect 217212 3236 217216 3292
rect 217152 3232 217216 3236
rect 217232 3292 217296 3296
rect 217232 3236 217236 3292
rect 217236 3236 217292 3292
rect 217292 3236 217296 3292
rect 217232 3232 217296 3236
rect 217312 3292 217376 3296
rect 217312 3236 217316 3292
rect 217316 3236 217372 3292
rect 217372 3236 217376 3292
rect 217312 3232 217376 3236
rect 252832 3292 252896 3296
rect 252832 3236 252836 3292
rect 252836 3236 252892 3292
rect 252892 3236 252896 3292
rect 252832 3232 252896 3236
rect 252912 3292 252976 3296
rect 252912 3236 252916 3292
rect 252916 3236 252972 3292
rect 252972 3236 252976 3292
rect 252912 3232 252976 3236
rect 252992 3292 253056 3296
rect 252992 3236 252996 3292
rect 252996 3236 253052 3292
rect 253052 3236 253056 3292
rect 252992 3232 253056 3236
rect 253072 3292 253136 3296
rect 253072 3236 253076 3292
rect 253076 3236 253132 3292
rect 253132 3236 253136 3292
rect 253072 3232 253136 3236
rect 253152 3292 253216 3296
rect 253152 3236 253156 3292
rect 253156 3236 253212 3292
rect 253212 3236 253216 3292
rect 253152 3232 253216 3236
rect 253232 3292 253296 3296
rect 253232 3236 253236 3292
rect 253236 3236 253292 3292
rect 253292 3236 253296 3292
rect 253232 3232 253296 3236
rect 253312 3292 253376 3296
rect 253312 3236 253316 3292
rect 253316 3236 253372 3292
rect 253372 3236 253376 3292
rect 253312 3232 253376 3236
rect 288832 3292 288896 3296
rect 288832 3236 288836 3292
rect 288836 3236 288892 3292
rect 288892 3236 288896 3292
rect 288832 3232 288896 3236
rect 288912 3292 288976 3296
rect 288912 3236 288916 3292
rect 288916 3236 288972 3292
rect 288972 3236 288976 3292
rect 288912 3232 288976 3236
rect 288992 3292 289056 3296
rect 288992 3236 288996 3292
rect 288996 3236 289052 3292
rect 289052 3236 289056 3292
rect 288992 3232 289056 3236
rect 289072 3292 289136 3296
rect 289072 3236 289076 3292
rect 289076 3236 289132 3292
rect 289132 3236 289136 3292
rect 289072 3232 289136 3236
rect 289152 3292 289216 3296
rect 289152 3236 289156 3292
rect 289156 3236 289212 3292
rect 289212 3236 289216 3292
rect 289152 3232 289216 3236
rect 289232 3292 289296 3296
rect 289232 3236 289236 3292
rect 289236 3236 289292 3292
rect 289292 3236 289296 3292
rect 289232 3232 289296 3236
rect 289312 3292 289376 3296
rect 289312 3236 289316 3292
rect 289316 3236 289372 3292
rect 289372 3236 289376 3292
rect 289312 3232 289376 3236
rect 324832 3292 324896 3296
rect 324832 3236 324836 3292
rect 324836 3236 324892 3292
rect 324892 3236 324896 3292
rect 324832 3232 324896 3236
rect 324912 3292 324976 3296
rect 324912 3236 324916 3292
rect 324916 3236 324972 3292
rect 324972 3236 324976 3292
rect 324912 3232 324976 3236
rect 324992 3292 325056 3296
rect 324992 3236 324996 3292
rect 324996 3236 325052 3292
rect 325052 3236 325056 3292
rect 324992 3232 325056 3236
rect 325072 3292 325136 3296
rect 325072 3236 325076 3292
rect 325076 3236 325132 3292
rect 325132 3236 325136 3292
rect 325072 3232 325136 3236
rect 325152 3292 325216 3296
rect 325152 3236 325156 3292
rect 325156 3236 325212 3292
rect 325212 3236 325216 3292
rect 325152 3232 325216 3236
rect 325232 3292 325296 3296
rect 325232 3236 325236 3292
rect 325236 3236 325292 3292
rect 325292 3236 325296 3292
rect 325232 3232 325296 3236
rect 325312 3292 325376 3296
rect 325312 3236 325316 3292
rect 325316 3236 325372 3292
rect 325372 3236 325376 3292
rect 325312 3232 325376 3236
rect 360832 3292 360896 3296
rect 360832 3236 360836 3292
rect 360836 3236 360892 3292
rect 360892 3236 360896 3292
rect 360832 3232 360896 3236
rect 360912 3292 360976 3296
rect 360912 3236 360916 3292
rect 360916 3236 360972 3292
rect 360972 3236 360976 3292
rect 360912 3232 360976 3236
rect 360992 3292 361056 3296
rect 360992 3236 360996 3292
rect 360996 3236 361052 3292
rect 361052 3236 361056 3292
rect 360992 3232 361056 3236
rect 361072 3292 361136 3296
rect 361072 3236 361076 3292
rect 361076 3236 361132 3292
rect 361132 3236 361136 3292
rect 361072 3232 361136 3236
rect 361152 3292 361216 3296
rect 361152 3236 361156 3292
rect 361156 3236 361212 3292
rect 361212 3236 361216 3292
rect 361152 3232 361216 3236
rect 361232 3292 361296 3296
rect 361232 3236 361236 3292
rect 361236 3236 361292 3292
rect 361292 3236 361296 3292
rect 361232 3232 361296 3236
rect 361312 3292 361376 3296
rect 361312 3236 361316 3292
rect 361316 3236 361372 3292
rect 361372 3236 361376 3292
rect 361312 3232 361376 3236
rect 396832 3292 396896 3296
rect 396832 3236 396836 3292
rect 396836 3236 396892 3292
rect 396892 3236 396896 3292
rect 396832 3232 396896 3236
rect 396912 3292 396976 3296
rect 396912 3236 396916 3292
rect 396916 3236 396972 3292
rect 396972 3236 396976 3292
rect 396912 3232 396976 3236
rect 396992 3292 397056 3296
rect 396992 3236 396996 3292
rect 396996 3236 397052 3292
rect 397052 3236 397056 3292
rect 396992 3232 397056 3236
rect 397072 3292 397136 3296
rect 397072 3236 397076 3292
rect 397076 3236 397132 3292
rect 397132 3236 397136 3292
rect 397072 3232 397136 3236
rect 397152 3292 397216 3296
rect 397152 3236 397156 3292
rect 397156 3236 397212 3292
rect 397212 3236 397216 3292
rect 397152 3232 397216 3236
rect 397232 3292 397296 3296
rect 397232 3236 397236 3292
rect 397236 3236 397292 3292
rect 397292 3236 397296 3292
rect 397232 3232 397296 3236
rect 397312 3292 397376 3296
rect 397312 3236 397316 3292
rect 397316 3236 397372 3292
rect 397372 3236 397376 3292
rect 397312 3232 397376 3236
rect 432832 3292 432896 3296
rect 432832 3236 432836 3292
rect 432836 3236 432892 3292
rect 432892 3236 432896 3292
rect 432832 3232 432896 3236
rect 432912 3292 432976 3296
rect 432912 3236 432916 3292
rect 432916 3236 432972 3292
rect 432972 3236 432976 3292
rect 432912 3232 432976 3236
rect 432992 3292 433056 3296
rect 432992 3236 432996 3292
rect 432996 3236 433052 3292
rect 433052 3236 433056 3292
rect 432992 3232 433056 3236
rect 433072 3292 433136 3296
rect 433072 3236 433076 3292
rect 433076 3236 433132 3292
rect 433132 3236 433136 3292
rect 433072 3232 433136 3236
rect 433152 3292 433216 3296
rect 433152 3236 433156 3292
rect 433156 3236 433212 3292
rect 433212 3236 433216 3292
rect 433152 3232 433216 3236
rect 433232 3292 433296 3296
rect 433232 3236 433236 3292
rect 433236 3236 433292 3292
rect 433292 3236 433296 3292
rect 433232 3232 433296 3236
rect 433312 3292 433376 3296
rect 433312 3236 433316 3292
rect 433316 3236 433372 3292
rect 433372 3236 433376 3292
rect 433312 3232 433376 3236
rect 468832 3292 468896 3296
rect 468832 3236 468836 3292
rect 468836 3236 468892 3292
rect 468892 3236 468896 3292
rect 468832 3232 468896 3236
rect 468912 3292 468976 3296
rect 468912 3236 468916 3292
rect 468916 3236 468972 3292
rect 468972 3236 468976 3292
rect 468912 3232 468976 3236
rect 468992 3292 469056 3296
rect 468992 3236 468996 3292
rect 468996 3236 469052 3292
rect 469052 3236 469056 3292
rect 468992 3232 469056 3236
rect 469072 3292 469136 3296
rect 469072 3236 469076 3292
rect 469076 3236 469132 3292
rect 469132 3236 469136 3292
rect 469072 3232 469136 3236
rect 469152 3292 469216 3296
rect 469152 3236 469156 3292
rect 469156 3236 469212 3292
rect 469212 3236 469216 3292
rect 469152 3232 469216 3236
rect 469232 3292 469296 3296
rect 469232 3236 469236 3292
rect 469236 3236 469292 3292
rect 469292 3236 469296 3292
rect 469232 3232 469296 3236
rect 469312 3292 469376 3296
rect 469312 3236 469316 3292
rect 469316 3236 469372 3292
rect 469372 3236 469376 3292
rect 469312 3232 469376 3236
rect 504832 3292 504896 3296
rect 504832 3236 504836 3292
rect 504836 3236 504892 3292
rect 504892 3236 504896 3292
rect 504832 3232 504896 3236
rect 504912 3292 504976 3296
rect 504912 3236 504916 3292
rect 504916 3236 504972 3292
rect 504972 3236 504976 3292
rect 504912 3232 504976 3236
rect 504992 3292 505056 3296
rect 504992 3236 504996 3292
rect 504996 3236 505052 3292
rect 505052 3236 505056 3292
rect 504992 3232 505056 3236
rect 505072 3292 505136 3296
rect 505072 3236 505076 3292
rect 505076 3236 505132 3292
rect 505132 3236 505136 3292
rect 505072 3232 505136 3236
rect 505152 3292 505216 3296
rect 505152 3236 505156 3292
rect 505156 3236 505212 3292
rect 505212 3236 505216 3292
rect 505152 3232 505216 3236
rect 505232 3292 505296 3296
rect 505232 3236 505236 3292
rect 505236 3236 505292 3292
rect 505292 3236 505296 3292
rect 505232 3232 505296 3236
rect 505312 3292 505376 3296
rect 505312 3236 505316 3292
rect 505316 3236 505372 3292
rect 505372 3236 505376 3292
rect 505312 3232 505376 3236
rect 540832 3292 540896 3296
rect 540832 3236 540836 3292
rect 540836 3236 540892 3292
rect 540892 3236 540896 3292
rect 540832 3232 540896 3236
rect 540912 3292 540976 3296
rect 540912 3236 540916 3292
rect 540916 3236 540972 3292
rect 540972 3236 540976 3292
rect 540912 3232 540976 3236
rect 540992 3292 541056 3296
rect 540992 3236 540996 3292
rect 540996 3236 541052 3292
rect 541052 3236 541056 3292
rect 540992 3232 541056 3236
rect 541072 3292 541136 3296
rect 541072 3236 541076 3292
rect 541076 3236 541132 3292
rect 541132 3236 541136 3292
rect 541072 3232 541136 3236
rect 541152 3292 541216 3296
rect 541152 3236 541156 3292
rect 541156 3236 541212 3292
rect 541212 3236 541216 3292
rect 541152 3232 541216 3236
rect 541232 3292 541296 3296
rect 541232 3236 541236 3292
rect 541236 3236 541292 3292
rect 541292 3236 541296 3292
rect 541232 3232 541296 3236
rect 541312 3292 541376 3296
rect 541312 3236 541316 3292
rect 541316 3236 541372 3292
rect 541372 3236 541376 3292
rect 541312 3232 541376 3236
rect 576832 3292 576896 3296
rect 576832 3236 576836 3292
rect 576836 3236 576892 3292
rect 576892 3236 576896 3292
rect 576832 3232 576896 3236
rect 576912 3292 576976 3296
rect 576912 3236 576916 3292
rect 576916 3236 576972 3292
rect 576972 3236 576976 3292
rect 576912 3232 576976 3236
rect 576992 3292 577056 3296
rect 576992 3236 576996 3292
rect 576996 3236 577052 3292
rect 577052 3236 577056 3292
rect 576992 3232 577056 3236
rect 577072 3292 577136 3296
rect 577072 3236 577076 3292
rect 577076 3236 577132 3292
rect 577132 3236 577136 3292
rect 577072 3232 577136 3236
rect 577152 3292 577216 3296
rect 577152 3236 577156 3292
rect 577156 3236 577212 3292
rect 577212 3236 577216 3292
rect 577152 3232 577216 3236
rect 577232 3292 577296 3296
rect 577232 3236 577236 3292
rect 577236 3236 577292 3292
rect 577292 3236 577296 3292
rect 577232 3232 577296 3236
rect 577312 3292 577376 3296
rect 577312 3236 577316 3292
rect 577316 3236 577372 3292
rect 577372 3236 577376 3292
rect 577312 3232 577376 3236
rect 18832 2748 18896 2752
rect 18832 2692 18836 2748
rect 18836 2692 18892 2748
rect 18892 2692 18896 2748
rect 18832 2688 18896 2692
rect 18912 2748 18976 2752
rect 18912 2692 18916 2748
rect 18916 2692 18972 2748
rect 18972 2692 18976 2748
rect 18912 2688 18976 2692
rect 18992 2748 19056 2752
rect 18992 2692 18996 2748
rect 18996 2692 19052 2748
rect 19052 2692 19056 2748
rect 18992 2688 19056 2692
rect 19072 2748 19136 2752
rect 19072 2692 19076 2748
rect 19076 2692 19132 2748
rect 19132 2692 19136 2748
rect 19072 2688 19136 2692
rect 19152 2748 19216 2752
rect 19152 2692 19156 2748
rect 19156 2692 19212 2748
rect 19212 2692 19216 2748
rect 19152 2688 19216 2692
rect 19232 2748 19296 2752
rect 19232 2692 19236 2748
rect 19236 2692 19292 2748
rect 19292 2692 19296 2748
rect 19232 2688 19296 2692
rect 19312 2748 19376 2752
rect 19312 2692 19316 2748
rect 19316 2692 19372 2748
rect 19372 2692 19376 2748
rect 19312 2688 19376 2692
rect 54832 2748 54896 2752
rect 54832 2692 54836 2748
rect 54836 2692 54892 2748
rect 54892 2692 54896 2748
rect 54832 2688 54896 2692
rect 54912 2748 54976 2752
rect 54912 2692 54916 2748
rect 54916 2692 54972 2748
rect 54972 2692 54976 2748
rect 54912 2688 54976 2692
rect 54992 2748 55056 2752
rect 54992 2692 54996 2748
rect 54996 2692 55052 2748
rect 55052 2692 55056 2748
rect 54992 2688 55056 2692
rect 55072 2748 55136 2752
rect 55072 2692 55076 2748
rect 55076 2692 55132 2748
rect 55132 2692 55136 2748
rect 55072 2688 55136 2692
rect 55152 2748 55216 2752
rect 55152 2692 55156 2748
rect 55156 2692 55212 2748
rect 55212 2692 55216 2748
rect 55152 2688 55216 2692
rect 55232 2748 55296 2752
rect 55232 2692 55236 2748
rect 55236 2692 55292 2748
rect 55292 2692 55296 2748
rect 55232 2688 55296 2692
rect 55312 2748 55376 2752
rect 55312 2692 55316 2748
rect 55316 2692 55372 2748
rect 55372 2692 55376 2748
rect 55312 2688 55376 2692
rect 90832 2748 90896 2752
rect 90832 2692 90836 2748
rect 90836 2692 90892 2748
rect 90892 2692 90896 2748
rect 90832 2688 90896 2692
rect 90912 2748 90976 2752
rect 90912 2692 90916 2748
rect 90916 2692 90972 2748
rect 90972 2692 90976 2748
rect 90912 2688 90976 2692
rect 90992 2748 91056 2752
rect 90992 2692 90996 2748
rect 90996 2692 91052 2748
rect 91052 2692 91056 2748
rect 90992 2688 91056 2692
rect 91072 2748 91136 2752
rect 91072 2692 91076 2748
rect 91076 2692 91132 2748
rect 91132 2692 91136 2748
rect 91072 2688 91136 2692
rect 91152 2748 91216 2752
rect 91152 2692 91156 2748
rect 91156 2692 91212 2748
rect 91212 2692 91216 2748
rect 91152 2688 91216 2692
rect 91232 2748 91296 2752
rect 91232 2692 91236 2748
rect 91236 2692 91292 2748
rect 91292 2692 91296 2748
rect 91232 2688 91296 2692
rect 91312 2748 91376 2752
rect 91312 2692 91316 2748
rect 91316 2692 91372 2748
rect 91372 2692 91376 2748
rect 91312 2688 91376 2692
rect 126832 2748 126896 2752
rect 126832 2692 126836 2748
rect 126836 2692 126892 2748
rect 126892 2692 126896 2748
rect 126832 2688 126896 2692
rect 126912 2748 126976 2752
rect 126912 2692 126916 2748
rect 126916 2692 126972 2748
rect 126972 2692 126976 2748
rect 126912 2688 126976 2692
rect 126992 2748 127056 2752
rect 126992 2692 126996 2748
rect 126996 2692 127052 2748
rect 127052 2692 127056 2748
rect 126992 2688 127056 2692
rect 127072 2748 127136 2752
rect 127072 2692 127076 2748
rect 127076 2692 127132 2748
rect 127132 2692 127136 2748
rect 127072 2688 127136 2692
rect 127152 2748 127216 2752
rect 127152 2692 127156 2748
rect 127156 2692 127212 2748
rect 127212 2692 127216 2748
rect 127152 2688 127216 2692
rect 127232 2748 127296 2752
rect 127232 2692 127236 2748
rect 127236 2692 127292 2748
rect 127292 2692 127296 2748
rect 127232 2688 127296 2692
rect 127312 2748 127376 2752
rect 127312 2692 127316 2748
rect 127316 2692 127372 2748
rect 127372 2692 127376 2748
rect 127312 2688 127376 2692
rect 162832 2748 162896 2752
rect 162832 2692 162836 2748
rect 162836 2692 162892 2748
rect 162892 2692 162896 2748
rect 162832 2688 162896 2692
rect 162912 2748 162976 2752
rect 162912 2692 162916 2748
rect 162916 2692 162972 2748
rect 162972 2692 162976 2748
rect 162912 2688 162976 2692
rect 162992 2748 163056 2752
rect 162992 2692 162996 2748
rect 162996 2692 163052 2748
rect 163052 2692 163056 2748
rect 162992 2688 163056 2692
rect 163072 2748 163136 2752
rect 163072 2692 163076 2748
rect 163076 2692 163132 2748
rect 163132 2692 163136 2748
rect 163072 2688 163136 2692
rect 163152 2748 163216 2752
rect 163152 2692 163156 2748
rect 163156 2692 163212 2748
rect 163212 2692 163216 2748
rect 163152 2688 163216 2692
rect 163232 2748 163296 2752
rect 163232 2692 163236 2748
rect 163236 2692 163292 2748
rect 163292 2692 163296 2748
rect 163232 2688 163296 2692
rect 163312 2748 163376 2752
rect 163312 2692 163316 2748
rect 163316 2692 163372 2748
rect 163372 2692 163376 2748
rect 163312 2688 163376 2692
rect 198832 2748 198896 2752
rect 198832 2692 198836 2748
rect 198836 2692 198892 2748
rect 198892 2692 198896 2748
rect 198832 2688 198896 2692
rect 198912 2748 198976 2752
rect 198912 2692 198916 2748
rect 198916 2692 198972 2748
rect 198972 2692 198976 2748
rect 198912 2688 198976 2692
rect 198992 2748 199056 2752
rect 198992 2692 198996 2748
rect 198996 2692 199052 2748
rect 199052 2692 199056 2748
rect 198992 2688 199056 2692
rect 199072 2748 199136 2752
rect 199072 2692 199076 2748
rect 199076 2692 199132 2748
rect 199132 2692 199136 2748
rect 199072 2688 199136 2692
rect 199152 2748 199216 2752
rect 199152 2692 199156 2748
rect 199156 2692 199212 2748
rect 199212 2692 199216 2748
rect 199152 2688 199216 2692
rect 199232 2748 199296 2752
rect 199232 2692 199236 2748
rect 199236 2692 199292 2748
rect 199292 2692 199296 2748
rect 199232 2688 199296 2692
rect 199312 2748 199376 2752
rect 199312 2692 199316 2748
rect 199316 2692 199372 2748
rect 199372 2692 199376 2748
rect 199312 2688 199376 2692
rect 234832 2748 234896 2752
rect 234832 2692 234836 2748
rect 234836 2692 234892 2748
rect 234892 2692 234896 2748
rect 234832 2688 234896 2692
rect 234912 2748 234976 2752
rect 234912 2692 234916 2748
rect 234916 2692 234972 2748
rect 234972 2692 234976 2748
rect 234912 2688 234976 2692
rect 234992 2748 235056 2752
rect 234992 2692 234996 2748
rect 234996 2692 235052 2748
rect 235052 2692 235056 2748
rect 234992 2688 235056 2692
rect 235072 2748 235136 2752
rect 235072 2692 235076 2748
rect 235076 2692 235132 2748
rect 235132 2692 235136 2748
rect 235072 2688 235136 2692
rect 235152 2748 235216 2752
rect 235152 2692 235156 2748
rect 235156 2692 235212 2748
rect 235212 2692 235216 2748
rect 235152 2688 235216 2692
rect 235232 2748 235296 2752
rect 235232 2692 235236 2748
rect 235236 2692 235292 2748
rect 235292 2692 235296 2748
rect 235232 2688 235296 2692
rect 235312 2748 235376 2752
rect 235312 2692 235316 2748
rect 235316 2692 235372 2748
rect 235372 2692 235376 2748
rect 235312 2688 235376 2692
rect 270832 2748 270896 2752
rect 270832 2692 270836 2748
rect 270836 2692 270892 2748
rect 270892 2692 270896 2748
rect 270832 2688 270896 2692
rect 270912 2748 270976 2752
rect 270912 2692 270916 2748
rect 270916 2692 270972 2748
rect 270972 2692 270976 2748
rect 270912 2688 270976 2692
rect 270992 2748 271056 2752
rect 270992 2692 270996 2748
rect 270996 2692 271052 2748
rect 271052 2692 271056 2748
rect 270992 2688 271056 2692
rect 271072 2748 271136 2752
rect 271072 2692 271076 2748
rect 271076 2692 271132 2748
rect 271132 2692 271136 2748
rect 271072 2688 271136 2692
rect 271152 2748 271216 2752
rect 271152 2692 271156 2748
rect 271156 2692 271212 2748
rect 271212 2692 271216 2748
rect 271152 2688 271216 2692
rect 271232 2748 271296 2752
rect 271232 2692 271236 2748
rect 271236 2692 271292 2748
rect 271292 2692 271296 2748
rect 271232 2688 271296 2692
rect 271312 2748 271376 2752
rect 271312 2692 271316 2748
rect 271316 2692 271372 2748
rect 271372 2692 271376 2748
rect 271312 2688 271376 2692
rect 306832 2748 306896 2752
rect 306832 2692 306836 2748
rect 306836 2692 306892 2748
rect 306892 2692 306896 2748
rect 306832 2688 306896 2692
rect 306912 2748 306976 2752
rect 306912 2692 306916 2748
rect 306916 2692 306972 2748
rect 306972 2692 306976 2748
rect 306912 2688 306976 2692
rect 306992 2748 307056 2752
rect 306992 2692 306996 2748
rect 306996 2692 307052 2748
rect 307052 2692 307056 2748
rect 306992 2688 307056 2692
rect 307072 2748 307136 2752
rect 307072 2692 307076 2748
rect 307076 2692 307132 2748
rect 307132 2692 307136 2748
rect 307072 2688 307136 2692
rect 307152 2748 307216 2752
rect 307152 2692 307156 2748
rect 307156 2692 307212 2748
rect 307212 2692 307216 2748
rect 307152 2688 307216 2692
rect 307232 2748 307296 2752
rect 307232 2692 307236 2748
rect 307236 2692 307292 2748
rect 307292 2692 307296 2748
rect 307232 2688 307296 2692
rect 307312 2748 307376 2752
rect 307312 2692 307316 2748
rect 307316 2692 307372 2748
rect 307372 2692 307376 2748
rect 307312 2688 307376 2692
rect 342832 2748 342896 2752
rect 342832 2692 342836 2748
rect 342836 2692 342892 2748
rect 342892 2692 342896 2748
rect 342832 2688 342896 2692
rect 342912 2748 342976 2752
rect 342912 2692 342916 2748
rect 342916 2692 342972 2748
rect 342972 2692 342976 2748
rect 342912 2688 342976 2692
rect 342992 2748 343056 2752
rect 342992 2692 342996 2748
rect 342996 2692 343052 2748
rect 343052 2692 343056 2748
rect 342992 2688 343056 2692
rect 343072 2748 343136 2752
rect 343072 2692 343076 2748
rect 343076 2692 343132 2748
rect 343132 2692 343136 2748
rect 343072 2688 343136 2692
rect 343152 2748 343216 2752
rect 343152 2692 343156 2748
rect 343156 2692 343212 2748
rect 343212 2692 343216 2748
rect 343152 2688 343216 2692
rect 343232 2748 343296 2752
rect 343232 2692 343236 2748
rect 343236 2692 343292 2748
rect 343292 2692 343296 2748
rect 343232 2688 343296 2692
rect 343312 2748 343376 2752
rect 343312 2692 343316 2748
rect 343316 2692 343372 2748
rect 343372 2692 343376 2748
rect 343312 2688 343376 2692
rect 378832 2748 378896 2752
rect 378832 2692 378836 2748
rect 378836 2692 378892 2748
rect 378892 2692 378896 2748
rect 378832 2688 378896 2692
rect 378912 2748 378976 2752
rect 378912 2692 378916 2748
rect 378916 2692 378972 2748
rect 378972 2692 378976 2748
rect 378912 2688 378976 2692
rect 378992 2748 379056 2752
rect 378992 2692 378996 2748
rect 378996 2692 379052 2748
rect 379052 2692 379056 2748
rect 378992 2688 379056 2692
rect 379072 2748 379136 2752
rect 379072 2692 379076 2748
rect 379076 2692 379132 2748
rect 379132 2692 379136 2748
rect 379072 2688 379136 2692
rect 379152 2748 379216 2752
rect 379152 2692 379156 2748
rect 379156 2692 379212 2748
rect 379212 2692 379216 2748
rect 379152 2688 379216 2692
rect 379232 2748 379296 2752
rect 379232 2692 379236 2748
rect 379236 2692 379292 2748
rect 379292 2692 379296 2748
rect 379232 2688 379296 2692
rect 379312 2748 379376 2752
rect 379312 2692 379316 2748
rect 379316 2692 379372 2748
rect 379372 2692 379376 2748
rect 379312 2688 379376 2692
rect 414832 2748 414896 2752
rect 414832 2692 414836 2748
rect 414836 2692 414892 2748
rect 414892 2692 414896 2748
rect 414832 2688 414896 2692
rect 414912 2748 414976 2752
rect 414912 2692 414916 2748
rect 414916 2692 414972 2748
rect 414972 2692 414976 2748
rect 414912 2688 414976 2692
rect 414992 2748 415056 2752
rect 414992 2692 414996 2748
rect 414996 2692 415052 2748
rect 415052 2692 415056 2748
rect 414992 2688 415056 2692
rect 415072 2748 415136 2752
rect 415072 2692 415076 2748
rect 415076 2692 415132 2748
rect 415132 2692 415136 2748
rect 415072 2688 415136 2692
rect 415152 2748 415216 2752
rect 415152 2692 415156 2748
rect 415156 2692 415212 2748
rect 415212 2692 415216 2748
rect 415152 2688 415216 2692
rect 415232 2748 415296 2752
rect 415232 2692 415236 2748
rect 415236 2692 415292 2748
rect 415292 2692 415296 2748
rect 415232 2688 415296 2692
rect 415312 2748 415376 2752
rect 415312 2692 415316 2748
rect 415316 2692 415372 2748
rect 415372 2692 415376 2748
rect 415312 2688 415376 2692
rect 450832 2748 450896 2752
rect 450832 2692 450836 2748
rect 450836 2692 450892 2748
rect 450892 2692 450896 2748
rect 450832 2688 450896 2692
rect 450912 2748 450976 2752
rect 450912 2692 450916 2748
rect 450916 2692 450972 2748
rect 450972 2692 450976 2748
rect 450912 2688 450976 2692
rect 450992 2748 451056 2752
rect 450992 2692 450996 2748
rect 450996 2692 451052 2748
rect 451052 2692 451056 2748
rect 450992 2688 451056 2692
rect 451072 2748 451136 2752
rect 451072 2692 451076 2748
rect 451076 2692 451132 2748
rect 451132 2692 451136 2748
rect 451072 2688 451136 2692
rect 451152 2748 451216 2752
rect 451152 2692 451156 2748
rect 451156 2692 451212 2748
rect 451212 2692 451216 2748
rect 451152 2688 451216 2692
rect 451232 2748 451296 2752
rect 451232 2692 451236 2748
rect 451236 2692 451292 2748
rect 451292 2692 451296 2748
rect 451232 2688 451296 2692
rect 451312 2748 451376 2752
rect 451312 2692 451316 2748
rect 451316 2692 451372 2748
rect 451372 2692 451376 2748
rect 451312 2688 451376 2692
rect 486832 2748 486896 2752
rect 486832 2692 486836 2748
rect 486836 2692 486892 2748
rect 486892 2692 486896 2748
rect 486832 2688 486896 2692
rect 486912 2748 486976 2752
rect 486912 2692 486916 2748
rect 486916 2692 486972 2748
rect 486972 2692 486976 2748
rect 486912 2688 486976 2692
rect 486992 2748 487056 2752
rect 486992 2692 486996 2748
rect 486996 2692 487052 2748
rect 487052 2692 487056 2748
rect 486992 2688 487056 2692
rect 487072 2748 487136 2752
rect 487072 2692 487076 2748
rect 487076 2692 487132 2748
rect 487132 2692 487136 2748
rect 487072 2688 487136 2692
rect 487152 2748 487216 2752
rect 487152 2692 487156 2748
rect 487156 2692 487212 2748
rect 487212 2692 487216 2748
rect 487152 2688 487216 2692
rect 487232 2748 487296 2752
rect 487232 2692 487236 2748
rect 487236 2692 487292 2748
rect 487292 2692 487296 2748
rect 487232 2688 487296 2692
rect 487312 2748 487376 2752
rect 487312 2692 487316 2748
rect 487316 2692 487372 2748
rect 487372 2692 487376 2748
rect 487312 2688 487376 2692
rect 522832 2748 522896 2752
rect 522832 2692 522836 2748
rect 522836 2692 522892 2748
rect 522892 2692 522896 2748
rect 522832 2688 522896 2692
rect 522912 2748 522976 2752
rect 522912 2692 522916 2748
rect 522916 2692 522972 2748
rect 522972 2692 522976 2748
rect 522912 2688 522976 2692
rect 522992 2748 523056 2752
rect 522992 2692 522996 2748
rect 522996 2692 523052 2748
rect 523052 2692 523056 2748
rect 522992 2688 523056 2692
rect 523072 2748 523136 2752
rect 523072 2692 523076 2748
rect 523076 2692 523132 2748
rect 523132 2692 523136 2748
rect 523072 2688 523136 2692
rect 523152 2748 523216 2752
rect 523152 2692 523156 2748
rect 523156 2692 523212 2748
rect 523212 2692 523216 2748
rect 523152 2688 523216 2692
rect 523232 2748 523296 2752
rect 523232 2692 523236 2748
rect 523236 2692 523292 2748
rect 523292 2692 523296 2748
rect 523232 2688 523296 2692
rect 523312 2748 523376 2752
rect 523312 2692 523316 2748
rect 523316 2692 523372 2748
rect 523372 2692 523376 2748
rect 523312 2688 523376 2692
rect 558832 2748 558896 2752
rect 558832 2692 558836 2748
rect 558836 2692 558892 2748
rect 558892 2692 558896 2748
rect 558832 2688 558896 2692
rect 558912 2748 558976 2752
rect 558912 2692 558916 2748
rect 558916 2692 558972 2748
rect 558972 2692 558976 2748
rect 558912 2688 558976 2692
rect 558992 2748 559056 2752
rect 558992 2692 558996 2748
rect 558996 2692 559052 2748
rect 559052 2692 559056 2748
rect 558992 2688 559056 2692
rect 559072 2748 559136 2752
rect 559072 2692 559076 2748
rect 559076 2692 559132 2748
rect 559132 2692 559136 2748
rect 559072 2688 559136 2692
rect 559152 2748 559216 2752
rect 559152 2692 559156 2748
rect 559156 2692 559212 2748
rect 559212 2692 559216 2748
rect 559152 2688 559216 2692
rect 559232 2748 559296 2752
rect 559232 2692 559236 2748
rect 559236 2692 559292 2748
rect 559292 2692 559296 2748
rect 559232 2688 559296 2692
rect 559312 2748 559376 2752
rect 559312 2692 559316 2748
rect 559316 2692 559372 2748
rect 559372 2692 559376 2748
rect 559312 2688 559376 2692
rect 36832 2204 36896 2208
rect 36832 2148 36836 2204
rect 36836 2148 36892 2204
rect 36892 2148 36896 2204
rect 36832 2144 36896 2148
rect 36912 2204 36976 2208
rect 36912 2148 36916 2204
rect 36916 2148 36972 2204
rect 36972 2148 36976 2204
rect 36912 2144 36976 2148
rect 36992 2204 37056 2208
rect 36992 2148 36996 2204
rect 36996 2148 37052 2204
rect 37052 2148 37056 2204
rect 36992 2144 37056 2148
rect 37072 2204 37136 2208
rect 37072 2148 37076 2204
rect 37076 2148 37132 2204
rect 37132 2148 37136 2204
rect 37072 2144 37136 2148
rect 37152 2204 37216 2208
rect 37152 2148 37156 2204
rect 37156 2148 37212 2204
rect 37212 2148 37216 2204
rect 37152 2144 37216 2148
rect 37232 2204 37296 2208
rect 37232 2148 37236 2204
rect 37236 2148 37292 2204
rect 37292 2148 37296 2204
rect 37232 2144 37296 2148
rect 37312 2204 37376 2208
rect 37312 2148 37316 2204
rect 37316 2148 37372 2204
rect 37372 2148 37376 2204
rect 37312 2144 37376 2148
rect 72832 2204 72896 2208
rect 72832 2148 72836 2204
rect 72836 2148 72892 2204
rect 72892 2148 72896 2204
rect 72832 2144 72896 2148
rect 72912 2204 72976 2208
rect 72912 2148 72916 2204
rect 72916 2148 72972 2204
rect 72972 2148 72976 2204
rect 72912 2144 72976 2148
rect 72992 2204 73056 2208
rect 72992 2148 72996 2204
rect 72996 2148 73052 2204
rect 73052 2148 73056 2204
rect 72992 2144 73056 2148
rect 73072 2204 73136 2208
rect 73072 2148 73076 2204
rect 73076 2148 73132 2204
rect 73132 2148 73136 2204
rect 73072 2144 73136 2148
rect 73152 2204 73216 2208
rect 73152 2148 73156 2204
rect 73156 2148 73212 2204
rect 73212 2148 73216 2204
rect 73152 2144 73216 2148
rect 73232 2204 73296 2208
rect 73232 2148 73236 2204
rect 73236 2148 73292 2204
rect 73292 2148 73296 2204
rect 73232 2144 73296 2148
rect 73312 2204 73376 2208
rect 73312 2148 73316 2204
rect 73316 2148 73372 2204
rect 73372 2148 73376 2204
rect 73312 2144 73376 2148
rect 108832 2204 108896 2208
rect 108832 2148 108836 2204
rect 108836 2148 108892 2204
rect 108892 2148 108896 2204
rect 108832 2144 108896 2148
rect 108912 2204 108976 2208
rect 108912 2148 108916 2204
rect 108916 2148 108972 2204
rect 108972 2148 108976 2204
rect 108912 2144 108976 2148
rect 108992 2204 109056 2208
rect 108992 2148 108996 2204
rect 108996 2148 109052 2204
rect 109052 2148 109056 2204
rect 108992 2144 109056 2148
rect 109072 2204 109136 2208
rect 109072 2148 109076 2204
rect 109076 2148 109132 2204
rect 109132 2148 109136 2204
rect 109072 2144 109136 2148
rect 109152 2204 109216 2208
rect 109152 2148 109156 2204
rect 109156 2148 109212 2204
rect 109212 2148 109216 2204
rect 109152 2144 109216 2148
rect 109232 2204 109296 2208
rect 109232 2148 109236 2204
rect 109236 2148 109292 2204
rect 109292 2148 109296 2204
rect 109232 2144 109296 2148
rect 109312 2204 109376 2208
rect 109312 2148 109316 2204
rect 109316 2148 109372 2204
rect 109372 2148 109376 2204
rect 109312 2144 109376 2148
rect 144832 2204 144896 2208
rect 144832 2148 144836 2204
rect 144836 2148 144892 2204
rect 144892 2148 144896 2204
rect 144832 2144 144896 2148
rect 144912 2204 144976 2208
rect 144912 2148 144916 2204
rect 144916 2148 144972 2204
rect 144972 2148 144976 2204
rect 144912 2144 144976 2148
rect 144992 2204 145056 2208
rect 144992 2148 144996 2204
rect 144996 2148 145052 2204
rect 145052 2148 145056 2204
rect 144992 2144 145056 2148
rect 145072 2204 145136 2208
rect 145072 2148 145076 2204
rect 145076 2148 145132 2204
rect 145132 2148 145136 2204
rect 145072 2144 145136 2148
rect 145152 2204 145216 2208
rect 145152 2148 145156 2204
rect 145156 2148 145212 2204
rect 145212 2148 145216 2204
rect 145152 2144 145216 2148
rect 145232 2204 145296 2208
rect 145232 2148 145236 2204
rect 145236 2148 145292 2204
rect 145292 2148 145296 2204
rect 145232 2144 145296 2148
rect 145312 2204 145376 2208
rect 145312 2148 145316 2204
rect 145316 2148 145372 2204
rect 145372 2148 145376 2204
rect 145312 2144 145376 2148
rect 180832 2204 180896 2208
rect 180832 2148 180836 2204
rect 180836 2148 180892 2204
rect 180892 2148 180896 2204
rect 180832 2144 180896 2148
rect 180912 2204 180976 2208
rect 180912 2148 180916 2204
rect 180916 2148 180972 2204
rect 180972 2148 180976 2204
rect 180912 2144 180976 2148
rect 180992 2204 181056 2208
rect 180992 2148 180996 2204
rect 180996 2148 181052 2204
rect 181052 2148 181056 2204
rect 180992 2144 181056 2148
rect 181072 2204 181136 2208
rect 181072 2148 181076 2204
rect 181076 2148 181132 2204
rect 181132 2148 181136 2204
rect 181072 2144 181136 2148
rect 181152 2204 181216 2208
rect 181152 2148 181156 2204
rect 181156 2148 181212 2204
rect 181212 2148 181216 2204
rect 181152 2144 181216 2148
rect 181232 2204 181296 2208
rect 181232 2148 181236 2204
rect 181236 2148 181292 2204
rect 181292 2148 181296 2204
rect 181232 2144 181296 2148
rect 181312 2204 181376 2208
rect 181312 2148 181316 2204
rect 181316 2148 181372 2204
rect 181372 2148 181376 2204
rect 181312 2144 181376 2148
rect 216832 2204 216896 2208
rect 216832 2148 216836 2204
rect 216836 2148 216892 2204
rect 216892 2148 216896 2204
rect 216832 2144 216896 2148
rect 216912 2204 216976 2208
rect 216912 2148 216916 2204
rect 216916 2148 216972 2204
rect 216972 2148 216976 2204
rect 216912 2144 216976 2148
rect 216992 2204 217056 2208
rect 216992 2148 216996 2204
rect 216996 2148 217052 2204
rect 217052 2148 217056 2204
rect 216992 2144 217056 2148
rect 217072 2204 217136 2208
rect 217072 2148 217076 2204
rect 217076 2148 217132 2204
rect 217132 2148 217136 2204
rect 217072 2144 217136 2148
rect 217152 2204 217216 2208
rect 217152 2148 217156 2204
rect 217156 2148 217212 2204
rect 217212 2148 217216 2204
rect 217152 2144 217216 2148
rect 217232 2204 217296 2208
rect 217232 2148 217236 2204
rect 217236 2148 217292 2204
rect 217292 2148 217296 2204
rect 217232 2144 217296 2148
rect 217312 2204 217376 2208
rect 217312 2148 217316 2204
rect 217316 2148 217372 2204
rect 217372 2148 217376 2204
rect 217312 2144 217376 2148
rect 252832 2204 252896 2208
rect 252832 2148 252836 2204
rect 252836 2148 252892 2204
rect 252892 2148 252896 2204
rect 252832 2144 252896 2148
rect 252912 2204 252976 2208
rect 252912 2148 252916 2204
rect 252916 2148 252972 2204
rect 252972 2148 252976 2204
rect 252912 2144 252976 2148
rect 252992 2204 253056 2208
rect 252992 2148 252996 2204
rect 252996 2148 253052 2204
rect 253052 2148 253056 2204
rect 252992 2144 253056 2148
rect 253072 2204 253136 2208
rect 253072 2148 253076 2204
rect 253076 2148 253132 2204
rect 253132 2148 253136 2204
rect 253072 2144 253136 2148
rect 253152 2204 253216 2208
rect 253152 2148 253156 2204
rect 253156 2148 253212 2204
rect 253212 2148 253216 2204
rect 253152 2144 253216 2148
rect 253232 2204 253296 2208
rect 253232 2148 253236 2204
rect 253236 2148 253292 2204
rect 253292 2148 253296 2204
rect 253232 2144 253296 2148
rect 253312 2204 253376 2208
rect 253312 2148 253316 2204
rect 253316 2148 253372 2204
rect 253372 2148 253376 2204
rect 253312 2144 253376 2148
rect 288832 2204 288896 2208
rect 288832 2148 288836 2204
rect 288836 2148 288892 2204
rect 288892 2148 288896 2204
rect 288832 2144 288896 2148
rect 288912 2204 288976 2208
rect 288912 2148 288916 2204
rect 288916 2148 288972 2204
rect 288972 2148 288976 2204
rect 288912 2144 288976 2148
rect 288992 2204 289056 2208
rect 288992 2148 288996 2204
rect 288996 2148 289052 2204
rect 289052 2148 289056 2204
rect 288992 2144 289056 2148
rect 289072 2204 289136 2208
rect 289072 2148 289076 2204
rect 289076 2148 289132 2204
rect 289132 2148 289136 2204
rect 289072 2144 289136 2148
rect 289152 2204 289216 2208
rect 289152 2148 289156 2204
rect 289156 2148 289212 2204
rect 289212 2148 289216 2204
rect 289152 2144 289216 2148
rect 289232 2204 289296 2208
rect 289232 2148 289236 2204
rect 289236 2148 289292 2204
rect 289292 2148 289296 2204
rect 289232 2144 289296 2148
rect 289312 2204 289376 2208
rect 289312 2148 289316 2204
rect 289316 2148 289372 2204
rect 289372 2148 289376 2204
rect 289312 2144 289376 2148
rect 324832 2204 324896 2208
rect 324832 2148 324836 2204
rect 324836 2148 324892 2204
rect 324892 2148 324896 2204
rect 324832 2144 324896 2148
rect 324912 2204 324976 2208
rect 324912 2148 324916 2204
rect 324916 2148 324972 2204
rect 324972 2148 324976 2204
rect 324912 2144 324976 2148
rect 324992 2204 325056 2208
rect 324992 2148 324996 2204
rect 324996 2148 325052 2204
rect 325052 2148 325056 2204
rect 324992 2144 325056 2148
rect 325072 2204 325136 2208
rect 325072 2148 325076 2204
rect 325076 2148 325132 2204
rect 325132 2148 325136 2204
rect 325072 2144 325136 2148
rect 325152 2204 325216 2208
rect 325152 2148 325156 2204
rect 325156 2148 325212 2204
rect 325212 2148 325216 2204
rect 325152 2144 325216 2148
rect 325232 2204 325296 2208
rect 325232 2148 325236 2204
rect 325236 2148 325292 2204
rect 325292 2148 325296 2204
rect 325232 2144 325296 2148
rect 325312 2204 325376 2208
rect 325312 2148 325316 2204
rect 325316 2148 325372 2204
rect 325372 2148 325376 2204
rect 325312 2144 325376 2148
rect 360832 2204 360896 2208
rect 360832 2148 360836 2204
rect 360836 2148 360892 2204
rect 360892 2148 360896 2204
rect 360832 2144 360896 2148
rect 360912 2204 360976 2208
rect 360912 2148 360916 2204
rect 360916 2148 360972 2204
rect 360972 2148 360976 2204
rect 360912 2144 360976 2148
rect 360992 2204 361056 2208
rect 360992 2148 360996 2204
rect 360996 2148 361052 2204
rect 361052 2148 361056 2204
rect 360992 2144 361056 2148
rect 361072 2204 361136 2208
rect 361072 2148 361076 2204
rect 361076 2148 361132 2204
rect 361132 2148 361136 2204
rect 361072 2144 361136 2148
rect 361152 2204 361216 2208
rect 361152 2148 361156 2204
rect 361156 2148 361212 2204
rect 361212 2148 361216 2204
rect 361152 2144 361216 2148
rect 361232 2204 361296 2208
rect 361232 2148 361236 2204
rect 361236 2148 361292 2204
rect 361292 2148 361296 2204
rect 361232 2144 361296 2148
rect 361312 2204 361376 2208
rect 361312 2148 361316 2204
rect 361316 2148 361372 2204
rect 361372 2148 361376 2204
rect 361312 2144 361376 2148
rect 396832 2204 396896 2208
rect 396832 2148 396836 2204
rect 396836 2148 396892 2204
rect 396892 2148 396896 2204
rect 396832 2144 396896 2148
rect 396912 2204 396976 2208
rect 396912 2148 396916 2204
rect 396916 2148 396972 2204
rect 396972 2148 396976 2204
rect 396912 2144 396976 2148
rect 396992 2204 397056 2208
rect 396992 2148 396996 2204
rect 396996 2148 397052 2204
rect 397052 2148 397056 2204
rect 396992 2144 397056 2148
rect 397072 2204 397136 2208
rect 397072 2148 397076 2204
rect 397076 2148 397132 2204
rect 397132 2148 397136 2204
rect 397072 2144 397136 2148
rect 397152 2204 397216 2208
rect 397152 2148 397156 2204
rect 397156 2148 397212 2204
rect 397212 2148 397216 2204
rect 397152 2144 397216 2148
rect 397232 2204 397296 2208
rect 397232 2148 397236 2204
rect 397236 2148 397292 2204
rect 397292 2148 397296 2204
rect 397232 2144 397296 2148
rect 397312 2204 397376 2208
rect 397312 2148 397316 2204
rect 397316 2148 397372 2204
rect 397372 2148 397376 2204
rect 397312 2144 397376 2148
rect 432832 2204 432896 2208
rect 432832 2148 432836 2204
rect 432836 2148 432892 2204
rect 432892 2148 432896 2204
rect 432832 2144 432896 2148
rect 432912 2204 432976 2208
rect 432912 2148 432916 2204
rect 432916 2148 432972 2204
rect 432972 2148 432976 2204
rect 432912 2144 432976 2148
rect 432992 2204 433056 2208
rect 432992 2148 432996 2204
rect 432996 2148 433052 2204
rect 433052 2148 433056 2204
rect 432992 2144 433056 2148
rect 433072 2204 433136 2208
rect 433072 2148 433076 2204
rect 433076 2148 433132 2204
rect 433132 2148 433136 2204
rect 433072 2144 433136 2148
rect 433152 2204 433216 2208
rect 433152 2148 433156 2204
rect 433156 2148 433212 2204
rect 433212 2148 433216 2204
rect 433152 2144 433216 2148
rect 433232 2204 433296 2208
rect 433232 2148 433236 2204
rect 433236 2148 433292 2204
rect 433292 2148 433296 2204
rect 433232 2144 433296 2148
rect 433312 2204 433376 2208
rect 433312 2148 433316 2204
rect 433316 2148 433372 2204
rect 433372 2148 433376 2204
rect 433312 2144 433376 2148
rect 468832 2204 468896 2208
rect 468832 2148 468836 2204
rect 468836 2148 468892 2204
rect 468892 2148 468896 2204
rect 468832 2144 468896 2148
rect 468912 2204 468976 2208
rect 468912 2148 468916 2204
rect 468916 2148 468972 2204
rect 468972 2148 468976 2204
rect 468912 2144 468976 2148
rect 468992 2204 469056 2208
rect 468992 2148 468996 2204
rect 468996 2148 469052 2204
rect 469052 2148 469056 2204
rect 468992 2144 469056 2148
rect 469072 2204 469136 2208
rect 469072 2148 469076 2204
rect 469076 2148 469132 2204
rect 469132 2148 469136 2204
rect 469072 2144 469136 2148
rect 469152 2204 469216 2208
rect 469152 2148 469156 2204
rect 469156 2148 469212 2204
rect 469212 2148 469216 2204
rect 469152 2144 469216 2148
rect 469232 2204 469296 2208
rect 469232 2148 469236 2204
rect 469236 2148 469292 2204
rect 469292 2148 469296 2204
rect 469232 2144 469296 2148
rect 469312 2204 469376 2208
rect 469312 2148 469316 2204
rect 469316 2148 469372 2204
rect 469372 2148 469376 2204
rect 469312 2144 469376 2148
rect 504832 2204 504896 2208
rect 504832 2148 504836 2204
rect 504836 2148 504892 2204
rect 504892 2148 504896 2204
rect 504832 2144 504896 2148
rect 504912 2204 504976 2208
rect 504912 2148 504916 2204
rect 504916 2148 504972 2204
rect 504972 2148 504976 2204
rect 504912 2144 504976 2148
rect 504992 2204 505056 2208
rect 504992 2148 504996 2204
rect 504996 2148 505052 2204
rect 505052 2148 505056 2204
rect 504992 2144 505056 2148
rect 505072 2204 505136 2208
rect 505072 2148 505076 2204
rect 505076 2148 505132 2204
rect 505132 2148 505136 2204
rect 505072 2144 505136 2148
rect 505152 2204 505216 2208
rect 505152 2148 505156 2204
rect 505156 2148 505212 2204
rect 505212 2148 505216 2204
rect 505152 2144 505216 2148
rect 505232 2204 505296 2208
rect 505232 2148 505236 2204
rect 505236 2148 505292 2204
rect 505292 2148 505296 2204
rect 505232 2144 505296 2148
rect 505312 2204 505376 2208
rect 505312 2148 505316 2204
rect 505316 2148 505372 2204
rect 505372 2148 505376 2204
rect 505312 2144 505376 2148
rect 540832 2204 540896 2208
rect 540832 2148 540836 2204
rect 540836 2148 540892 2204
rect 540892 2148 540896 2204
rect 540832 2144 540896 2148
rect 540912 2204 540976 2208
rect 540912 2148 540916 2204
rect 540916 2148 540972 2204
rect 540972 2148 540976 2204
rect 540912 2144 540976 2148
rect 540992 2204 541056 2208
rect 540992 2148 540996 2204
rect 540996 2148 541052 2204
rect 541052 2148 541056 2204
rect 540992 2144 541056 2148
rect 541072 2204 541136 2208
rect 541072 2148 541076 2204
rect 541076 2148 541132 2204
rect 541132 2148 541136 2204
rect 541072 2144 541136 2148
rect 541152 2204 541216 2208
rect 541152 2148 541156 2204
rect 541156 2148 541212 2204
rect 541212 2148 541216 2204
rect 541152 2144 541216 2148
rect 541232 2204 541296 2208
rect 541232 2148 541236 2204
rect 541236 2148 541292 2204
rect 541292 2148 541296 2204
rect 541232 2144 541296 2148
rect 541312 2204 541376 2208
rect 541312 2148 541316 2204
rect 541316 2148 541372 2204
rect 541372 2148 541376 2204
rect 541312 2144 541376 2148
rect 576832 2204 576896 2208
rect 576832 2148 576836 2204
rect 576836 2148 576892 2204
rect 576892 2148 576896 2204
rect 576832 2144 576896 2148
rect 576912 2204 576976 2208
rect 576912 2148 576916 2204
rect 576916 2148 576972 2204
rect 576972 2148 576976 2204
rect 576912 2144 576976 2148
rect 576992 2204 577056 2208
rect 576992 2148 576996 2204
rect 576996 2148 577052 2204
rect 577052 2148 577056 2204
rect 576992 2144 577056 2148
rect 577072 2204 577136 2208
rect 577072 2148 577076 2204
rect 577076 2148 577132 2204
rect 577132 2148 577136 2204
rect 577072 2144 577136 2148
rect 577152 2204 577216 2208
rect 577152 2148 577156 2204
rect 577156 2148 577212 2204
rect 577212 2148 577216 2204
rect 577152 2144 577216 2148
rect 577232 2204 577296 2208
rect 577232 2148 577236 2204
rect 577236 2148 577292 2204
rect 577292 2148 577296 2204
rect 577232 2144 577296 2148
rect 577312 2204 577376 2208
rect 577312 2148 577316 2204
rect 577316 2148 577372 2204
rect 577372 2148 577376 2204
rect 577312 2144 577376 2148
<< metal4 >>
rect -8576 711418 -7976 711440
rect -8576 711182 -8394 711418
rect -8158 711182 -7976 711418
rect -8576 711098 -7976 711182
rect -8576 710862 -8394 711098
rect -8158 710862 -7976 711098
rect -8576 679254 -7976 710862
rect -8576 679018 -8394 679254
rect -8158 679018 -7976 679254
rect -8576 678934 -7976 679018
rect -8576 678698 -8394 678934
rect -8158 678698 -7976 678934
rect -8576 643254 -7976 678698
rect -8576 643018 -8394 643254
rect -8158 643018 -7976 643254
rect -8576 642934 -7976 643018
rect -8576 642698 -8394 642934
rect -8158 642698 -7976 642934
rect -8576 607254 -7976 642698
rect -8576 607018 -8394 607254
rect -8158 607018 -7976 607254
rect -8576 606934 -7976 607018
rect -8576 606698 -8394 606934
rect -8158 606698 -7976 606934
rect -8576 571254 -7976 606698
rect -8576 571018 -8394 571254
rect -8158 571018 -7976 571254
rect -8576 570934 -7976 571018
rect -8576 570698 -8394 570934
rect -8158 570698 -7976 570934
rect -8576 535254 -7976 570698
rect -8576 535018 -8394 535254
rect -8158 535018 -7976 535254
rect -8576 534934 -7976 535018
rect -8576 534698 -8394 534934
rect -8158 534698 -7976 534934
rect -8576 499254 -7976 534698
rect -8576 499018 -8394 499254
rect -8158 499018 -7976 499254
rect -8576 498934 -7976 499018
rect -8576 498698 -8394 498934
rect -8158 498698 -7976 498934
rect -8576 463254 -7976 498698
rect -8576 463018 -8394 463254
rect -8158 463018 -7976 463254
rect -8576 462934 -7976 463018
rect -8576 462698 -8394 462934
rect -8158 462698 -7976 462934
rect -8576 427254 -7976 462698
rect -8576 427018 -8394 427254
rect -8158 427018 -7976 427254
rect -8576 426934 -7976 427018
rect -8576 426698 -8394 426934
rect -8158 426698 -7976 426934
rect -8576 391254 -7976 426698
rect -8576 391018 -8394 391254
rect -8158 391018 -7976 391254
rect -8576 390934 -7976 391018
rect -8576 390698 -8394 390934
rect -8158 390698 -7976 390934
rect -8576 355254 -7976 390698
rect -8576 355018 -8394 355254
rect -8158 355018 -7976 355254
rect -8576 354934 -7976 355018
rect -8576 354698 -8394 354934
rect -8158 354698 -7976 354934
rect -8576 319254 -7976 354698
rect -8576 319018 -8394 319254
rect -8158 319018 -7976 319254
rect -8576 318934 -7976 319018
rect -8576 318698 -8394 318934
rect -8158 318698 -7976 318934
rect -8576 283254 -7976 318698
rect -8576 283018 -8394 283254
rect -8158 283018 -7976 283254
rect -8576 282934 -7976 283018
rect -8576 282698 -8394 282934
rect -8158 282698 -7976 282934
rect -8576 247254 -7976 282698
rect -8576 247018 -8394 247254
rect -8158 247018 -7976 247254
rect -8576 246934 -7976 247018
rect -8576 246698 -8394 246934
rect -8158 246698 -7976 246934
rect -8576 211254 -7976 246698
rect -8576 211018 -8394 211254
rect -8158 211018 -7976 211254
rect -8576 210934 -7976 211018
rect -8576 210698 -8394 210934
rect -8158 210698 -7976 210934
rect -8576 175254 -7976 210698
rect -8576 175018 -8394 175254
rect -8158 175018 -7976 175254
rect -8576 174934 -7976 175018
rect -8576 174698 -8394 174934
rect -8158 174698 -7976 174934
rect -8576 139254 -7976 174698
rect -8576 139018 -8394 139254
rect -8158 139018 -7976 139254
rect -8576 138934 -7976 139018
rect -8576 138698 -8394 138934
rect -8158 138698 -7976 138934
rect -8576 103254 -7976 138698
rect -8576 103018 -8394 103254
rect -8158 103018 -7976 103254
rect -8576 102934 -7976 103018
rect -8576 102698 -8394 102934
rect -8158 102698 -7976 102934
rect -8576 67254 -7976 102698
rect -8576 67018 -8394 67254
rect -8158 67018 -7976 67254
rect -8576 66934 -7976 67018
rect -8576 66698 -8394 66934
rect -8158 66698 -7976 66934
rect -8576 31254 -7976 66698
rect -8576 31018 -8394 31254
rect -8158 31018 -7976 31254
rect -8576 30934 -7976 31018
rect -8576 30698 -8394 30934
rect -8158 30698 -7976 30934
rect -8576 -6926 -7976 30698
rect -7636 710478 -7036 710500
rect -7636 710242 -7454 710478
rect -7218 710242 -7036 710478
rect -7636 710158 -7036 710242
rect -7636 709922 -7454 710158
rect -7218 709922 -7036 710158
rect -7636 697254 -7036 709922
rect 11604 710478 12204 711440
rect 11604 710242 11786 710478
rect 12022 710242 12204 710478
rect 11604 710158 12204 710242
rect 11604 709922 11786 710158
rect 12022 709922 12204 710158
rect -7636 697018 -7454 697254
rect -7218 697018 -7036 697254
rect -7636 696934 -7036 697018
rect -7636 696698 -7454 696934
rect -7218 696698 -7036 696934
rect -7636 661254 -7036 696698
rect -7636 661018 -7454 661254
rect -7218 661018 -7036 661254
rect -7636 660934 -7036 661018
rect -7636 660698 -7454 660934
rect -7218 660698 -7036 660934
rect -7636 625254 -7036 660698
rect -7636 625018 -7454 625254
rect -7218 625018 -7036 625254
rect -7636 624934 -7036 625018
rect -7636 624698 -7454 624934
rect -7218 624698 -7036 624934
rect -7636 589254 -7036 624698
rect -7636 589018 -7454 589254
rect -7218 589018 -7036 589254
rect -7636 588934 -7036 589018
rect -7636 588698 -7454 588934
rect -7218 588698 -7036 588934
rect -7636 553254 -7036 588698
rect -7636 553018 -7454 553254
rect -7218 553018 -7036 553254
rect -7636 552934 -7036 553018
rect -7636 552698 -7454 552934
rect -7218 552698 -7036 552934
rect -7636 517254 -7036 552698
rect -7636 517018 -7454 517254
rect -7218 517018 -7036 517254
rect -7636 516934 -7036 517018
rect -7636 516698 -7454 516934
rect -7218 516698 -7036 516934
rect -7636 481254 -7036 516698
rect -7636 481018 -7454 481254
rect -7218 481018 -7036 481254
rect -7636 480934 -7036 481018
rect -7636 480698 -7454 480934
rect -7218 480698 -7036 480934
rect -7636 445254 -7036 480698
rect -7636 445018 -7454 445254
rect -7218 445018 -7036 445254
rect -7636 444934 -7036 445018
rect -7636 444698 -7454 444934
rect -7218 444698 -7036 444934
rect -7636 409254 -7036 444698
rect -7636 409018 -7454 409254
rect -7218 409018 -7036 409254
rect -7636 408934 -7036 409018
rect -7636 408698 -7454 408934
rect -7218 408698 -7036 408934
rect -7636 373254 -7036 408698
rect -7636 373018 -7454 373254
rect -7218 373018 -7036 373254
rect -7636 372934 -7036 373018
rect -7636 372698 -7454 372934
rect -7218 372698 -7036 372934
rect -7636 337254 -7036 372698
rect -7636 337018 -7454 337254
rect -7218 337018 -7036 337254
rect -7636 336934 -7036 337018
rect -7636 336698 -7454 336934
rect -7218 336698 -7036 336934
rect -7636 301254 -7036 336698
rect -7636 301018 -7454 301254
rect -7218 301018 -7036 301254
rect -7636 300934 -7036 301018
rect -7636 300698 -7454 300934
rect -7218 300698 -7036 300934
rect -7636 265254 -7036 300698
rect -7636 265018 -7454 265254
rect -7218 265018 -7036 265254
rect -7636 264934 -7036 265018
rect -7636 264698 -7454 264934
rect -7218 264698 -7036 264934
rect -7636 229254 -7036 264698
rect -7636 229018 -7454 229254
rect -7218 229018 -7036 229254
rect -7636 228934 -7036 229018
rect -7636 228698 -7454 228934
rect -7218 228698 -7036 228934
rect -7636 193254 -7036 228698
rect -7636 193018 -7454 193254
rect -7218 193018 -7036 193254
rect -7636 192934 -7036 193018
rect -7636 192698 -7454 192934
rect -7218 192698 -7036 192934
rect -7636 157254 -7036 192698
rect -7636 157018 -7454 157254
rect -7218 157018 -7036 157254
rect -7636 156934 -7036 157018
rect -7636 156698 -7454 156934
rect -7218 156698 -7036 156934
rect -7636 121254 -7036 156698
rect -7636 121018 -7454 121254
rect -7218 121018 -7036 121254
rect -7636 120934 -7036 121018
rect -7636 120698 -7454 120934
rect -7218 120698 -7036 120934
rect -7636 85254 -7036 120698
rect -7636 85018 -7454 85254
rect -7218 85018 -7036 85254
rect -7636 84934 -7036 85018
rect -7636 84698 -7454 84934
rect -7218 84698 -7036 84934
rect -7636 49254 -7036 84698
rect -7636 49018 -7454 49254
rect -7218 49018 -7036 49254
rect -7636 48934 -7036 49018
rect -7636 48698 -7454 48934
rect -7218 48698 -7036 48934
rect -7636 13254 -7036 48698
rect -7636 13018 -7454 13254
rect -7218 13018 -7036 13254
rect -7636 12934 -7036 13018
rect -7636 12698 -7454 12934
rect -7218 12698 -7036 12934
rect -7636 -5986 -7036 12698
rect -6696 709538 -6096 709560
rect -6696 709302 -6514 709538
rect -6278 709302 -6096 709538
rect -6696 709218 -6096 709302
rect -6696 708982 -6514 709218
rect -6278 708982 -6096 709218
rect -6696 675654 -6096 708982
rect -6696 675418 -6514 675654
rect -6278 675418 -6096 675654
rect -6696 675334 -6096 675418
rect -6696 675098 -6514 675334
rect -6278 675098 -6096 675334
rect -6696 639654 -6096 675098
rect -6696 639418 -6514 639654
rect -6278 639418 -6096 639654
rect -6696 639334 -6096 639418
rect -6696 639098 -6514 639334
rect -6278 639098 -6096 639334
rect -6696 603654 -6096 639098
rect -6696 603418 -6514 603654
rect -6278 603418 -6096 603654
rect -6696 603334 -6096 603418
rect -6696 603098 -6514 603334
rect -6278 603098 -6096 603334
rect -6696 567654 -6096 603098
rect -6696 567418 -6514 567654
rect -6278 567418 -6096 567654
rect -6696 567334 -6096 567418
rect -6696 567098 -6514 567334
rect -6278 567098 -6096 567334
rect -6696 531654 -6096 567098
rect -6696 531418 -6514 531654
rect -6278 531418 -6096 531654
rect -6696 531334 -6096 531418
rect -6696 531098 -6514 531334
rect -6278 531098 -6096 531334
rect -6696 495654 -6096 531098
rect -6696 495418 -6514 495654
rect -6278 495418 -6096 495654
rect -6696 495334 -6096 495418
rect -6696 495098 -6514 495334
rect -6278 495098 -6096 495334
rect -6696 459654 -6096 495098
rect -6696 459418 -6514 459654
rect -6278 459418 -6096 459654
rect -6696 459334 -6096 459418
rect -6696 459098 -6514 459334
rect -6278 459098 -6096 459334
rect -6696 423654 -6096 459098
rect -6696 423418 -6514 423654
rect -6278 423418 -6096 423654
rect -6696 423334 -6096 423418
rect -6696 423098 -6514 423334
rect -6278 423098 -6096 423334
rect -6696 387654 -6096 423098
rect -6696 387418 -6514 387654
rect -6278 387418 -6096 387654
rect -6696 387334 -6096 387418
rect -6696 387098 -6514 387334
rect -6278 387098 -6096 387334
rect -6696 351654 -6096 387098
rect -6696 351418 -6514 351654
rect -6278 351418 -6096 351654
rect -6696 351334 -6096 351418
rect -6696 351098 -6514 351334
rect -6278 351098 -6096 351334
rect -6696 315654 -6096 351098
rect -6696 315418 -6514 315654
rect -6278 315418 -6096 315654
rect -6696 315334 -6096 315418
rect -6696 315098 -6514 315334
rect -6278 315098 -6096 315334
rect -6696 279654 -6096 315098
rect -6696 279418 -6514 279654
rect -6278 279418 -6096 279654
rect -6696 279334 -6096 279418
rect -6696 279098 -6514 279334
rect -6278 279098 -6096 279334
rect -6696 243654 -6096 279098
rect -6696 243418 -6514 243654
rect -6278 243418 -6096 243654
rect -6696 243334 -6096 243418
rect -6696 243098 -6514 243334
rect -6278 243098 -6096 243334
rect -6696 207654 -6096 243098
rect -6696 207418 -6514 207654
rect -6278 207418 -6096 207654
rect -6696 207334 -6096 207418
rect -6696 207098 -6514 207334
rect -6278 207098 -6096 207334
rect -6696 171654 -6096 207098
rect -6696 171418 -6514 171654
rect -6278 171418 -6096 171654
rect -6696 171334 -6096 171418
rect -6696 171098 -6514 171334
rect -6278 171098 -6096 171334
rect -6696 135654 -6096 171098
rect -6696 135418 -6514 135654
rect -6278 135418 -6096 135654
rect -6696 135334 -6096 135418
rect -6696 135098 -6514 135334
rect -6278 135098 -6096 135334
rect -6696 99654 -6096 135098
rect -6696 99418 -6514 99654
rect -6278 99418 -6096 99654
rect -6696 99334 -6096 99418
rect -6696 99098 -6514 99334
rect -6278 99098 -6096 99334
rect -6696 63654 -6096 99098
rect -6696 63418 -6514 63654
rect -6278 63418 -6096 63654
rect -6696 63334 -6096 63418
rect -6696 63098 -6514 63334
rect -6278 63098 -6096 63334
rect -6696 27654 -6096 63098
rect -6696 27418 -6514 27654
rect -6278 27418 -6096 27654
rect -6696 27334 -6096 27418
rect -6696 27098 -6514 27334
rect -6278 27098 -6096 27334
rect -6696 -5046 -6096 27098
rect -5756 708598 -5156 708620
rect -5756 708362 -5574 708598
rect -5338 708362 -5156 708598
rect -5756 708278 -5156 708362
rect -5756 708042 -5574 708278
rect -5338 708042 -5156 708278
rect -5756 693654 -5156 708042
rect 8004 708598 8604 709560
rect 8004 708362 8186 708598
rect 8422 708362 8604 708598
rect 8004 708278 8604 708362
rect 8004 708042 8186 708278
rect 8422 708042 8604 708278
rect -5756 693418 -5574 693654
rect -5338 693418 -5156 693654
rect -5756 693334 -5156 693418
rect -5756 693098 -5574 693334
rect -5338 693098 -5156 693334
rect -5756 657654 -5156 693098
rect -5756 657418 -5574 657654
rect -5338 657418 -5156 657654
rect -5756 657334 -5156 657418
rect -5756 657098 -5574 657334
rect -5338 657098 -5156 657334
rect -5756 621654 -5156 657098
rect -5756 621418 -5574 621654
rect -5338 621418 -5156 621654
rect -5756 621334 -5156 621418
rect -5756 621098 -5574 621334
rect -5338 621098 -5156 621334
rect -5756 585654 -5156 621098
rect -5756 585418 -5574 585654
rect -5338 585418 -5156 585654
rect -5756 585334 -5156 585418
rect -5756 585098 -5574 585334
rect -5338 585098 -5156 585334
rect -5756 549654 -5156 585098
rect -5756 549418 -5574 549654
rect -5338 549418 -5156 549654
rect -5756 549334 -5156 549418
rect -5756 549098 -5574 549334
rect -5338 549098 -5156 549334
rect -5756 513654 -5156 549098
rect -5756 513418 -5574 513654
rect -5338 513418 -5156 513654
rect -5756 513334 -5156 513418
rect -5756 513098 -5574 513334
rect -5338 513098 -5156 513334
rect -5756 477654 -5156 513098
rect -5756 477418 -5574 477654
rect -5338 477418 -5156 477654
rect -5756 477334 -5156 477418
rect -5756 477098 -5574 477334
rect -5338 477098 -5156 477334
rect -5756 441654 -5156 477098
rect -5756 441418 -5574 441654
rect -5338 441418 -5156 441654
rect -5756 441334 -5156 441418
rect -5756 441098 -5574 441334
rect -5338 441098 -5156 441334
rect -5756 405654 -5156 441098
rect -5756 405418 -5574 405654
rect -5338 405418 -5156 405654
rect -5756 405334 -5156 405418
rect -5756 405098 -5574 405334
rect -5338 405098 -5156 405334
rect -5756 369654 -5156 405098
rect -5756 369418 -5574 369654
rect -5338 369418 -5156 369654
rect -5756 369334 -5156 369418
rect -5756 369098 -5574 369334
rect -5338 369098 -5156 369334
rect -5756 333654 -5156 369098
rect -5756 333418 -5574 333654
rect -5338 333418 -5156 333654
rect -5756 333334 -5156 333418
rect -5756 333098 -5574 333334
rect -5338 333098 -5156 333334
rect -5756 297654 -5156 333098
rect -5756 297418 -5574 297654
rect -5338 297418 -5156 297654
rect -5756 297334 -5156 297418
rect -5756 297098 -5574 297334
rect -5338 297098 -5156 297334
rect -5756 261654 -5156 297098
rect -5756 261418 -5574 261654
rect -5338 261418 -5156 261654
rect -5756 261334 -5156 261418
rect -5756 261098 -5574 261334
rect -5338 261098 -5156 261334
rect -5756 225654 -5156 261098
rect -5756 225418 -5574 225654
rect -5338 225418 -5156 225654
rect -5756 225334 -5156 225418
rect -5756 225098 -5574 225334
rect -5338 225098 -5156 225334
rect -5756 189654 -5156 225098
rect -5756 189418 -5574 189654
rect -5338 189418 -5156 189654
rect -5756 189334 -5156 189418
rect -5756 189098 -5574 189334
rect -5338 189098 -5156 189334
rect -5756 153654 -5156 189098
rect -5756 153418 -5574 153654
rect -5338 153418 -5156 153654
rect -5756 153334 -5156 153418
rect -5756 153098 -5574 153334
rect -5338 153098 -5156 153334
rect -5756 117654 -5156 153098
rect -5756 117418 -5574 117654
rect -5338 117418 -5156 117654
rect -5756 117334 -5156 117418
rect -5756 117098 -5574 117334
rect -5338 117098 -5156 117334
rect -5756 81654 -5156 117098
rect -5756 81418 -5574 81654
rect -5338 81418 -5156 81654
rect -5756 81334 -5156 81418
rect -5756 81098 -5574 81334
rect -5338 81098 -5156 81334
rect -5756 45654 -5156 81098
rect -5756 45418 -5574 45654
rect -5338 45418 -5156 45654
rect -5756 45334 -5156 45418
rect -5756 45098 -5574 45334
rect -5338 45098 -5156 45334
rect -5756 9654 -5156 45098
rect -5756 9418 -5574 9654
rect -5338 9418 -5156 9654
rect -5756 9334 -5156 9418
rect -5756 9098 -5574 9334
rect -5338 9098 -5156 9334
rect -5756 -4106 -5156 9098
rect -4816 707658 -4216 707680
rect -4816 707422 -4634 707658
rect -4398 707422 -4216 707658
rect -4816 707338 -4216 707422
rect -4816 707102 -4634 707338
rect -4398 707102 -4216 707338
rect -4816 672054 -4216 707102
rect -4816 671818 -4634 672054
rect -4398 671818 -4216 672054
rect -4816 671734 -4216 671818
rect -4816 671498 -4634 671734
rect -4398 671498 -4216 671734
rect -4816 636054 -4216 671498
rect -4816 635818 -4634 636054
rect -4398 635818 -4216 636054
rect -4816 635734 -4216 635818
rect -4816 635498 -4634 635734
rect -4398 635498 -4216 635734
rect -4816 600054 -4216 635498
rect -4816 599818 -4634 600054
rect -4398 599818 -4216 600054
rect -4816 599734 -4216 599818
rect -4816 599498 -4634 599734
rect -4398 599498 -4216 599734
rect -4816 564054 -4216 599498
rect -4816 563818 -4634 564054
rect -4398 563818 -4216 564054
rect -4816 563734 -4216 563818
rect -4816 563498 -4634 563734
rect -4398 563498 -4216 563734
rect -4816 528054 -4216 563498
rect -4816 527818 -4634 528054
rect -4398 527818 -4216 528054
rect -4816 527734 -4216 527818
rect -4816 527498 -4634 527734
rect -4398 527498 -4216 527734
rect -4816 492054 -4216 527498
rect -4816 491818 -4634 492054
rect -4398 491818 -4216 492054
rect -4816 491734 -4216 491818
rect -4816 491498 -4634 491734
rect -4398 491498 -4216 491734
rect -4816 456054 -4216 491498
rect -4816 455818 -4634 456054
rect -4398 455818 -4216 456054
rect -4816 455734 -4216 455818
rect -4816 455498 -4634 455734
rect -4398 455498 -4216 455734
rect -4816 420054 -4216 455498
rect -4816 419818 -4634 420054
rect -4398 419818 -4216 420054
rect -4816 419734 -4216 419818
rect -4816 419498 -4634 419734
rect -4398 419498 -4216 419734
rect -4816 384054 -4216 419498
rect -4816 383818 -4634 384054
rect -4398 383818 -4216 384054
rect -4816 383734 -4216 383818
rect -4816 383498 -4634 383734
rect -4398 383498 -4216 383734
rect -4816 348054 -4216 383498
rect -4816 347818 -4634 348054
rect -4398 347818 -4216 348054
rect -4816 347734 -4216 347818
rect -4816 347498 -4634 347734
rect -4398 347498 -4216 347734
rect -4816 312054 -4216 347498
rect -4816 311818 -4634 312054
rect -4398 311818 -4216 312054
rect -4816 311734 -4216 311818
rect -4816 311498 -4634 311734
rect -4398 311498 -4216 311734
rect -4816 276054 -4216 311498
rect -4816 275818 -4634 276054
rect -4398 275818 -4216 276054
rect -4816 275734 -4216 275818
rect -4816 275498 -4634 275734
rect -4398 275498 -4216 275734
rect -4816 240054 -4216 275498
rect -4816 239818 -4634 240054
rect -4398 239818 -4216 240054
rect -4816 239734 -4216 239818
rect -4816 239498 -4634 239734
rect -4398 239498 -4216 239734
rect -4816 204054 -4216 239498
rect -4816 203818 -4634 204054
rect -4398 203818 -4216 204054
rect -4816 203734 -4216 203818
rect -4816 203498 -4634 203734
rect -4398 203498 -4216 203734
rect -4816 168054 -4216 203498
rect -4816 167818 -4634 168054
rect -4398 167818 -4216 168054
rect -4816 167734 -4216 167818
rect -4816 167498 -4634 167734
rect -4398 167498 -4216 167734
rect -4816 132054 -4216 167498
rect -4816 131818 -4634 132054
rect -4398 131818 -4216 132054
rect -4816 131734 -4216 131818
rect -4816 131498 -4634 131734
rect -4398 131498 -4216 131734
rect -4816 96054 -4216 131498
rect -4816 95818 -4634 96054
rect -4398 95818 -4216 96054
rect -4816 95734 -4216 95818
rect -4816 95498 -4634 95734
rect -4398 95498 -4216 95734
rect -4816 60054 -4216 95498
rect -4816 59818 -4634 60054
rect -4398 59818 -4216 60054
rect -4816 59734 -4216 59818
rect -4816 59498 -4634 59734
rect -4398 59498 -4216 59734
rect -4816 24054 -4216 59498
rect -4816 23818 -4634 24054
rect -4398 23818 -4216 24054
rect -4816 23734 -4216 23818
rect -4816 23498 -4634 23734
rect -4398 23498 -4216 23734
rect -4816 -3166 -4216 23498
rect -3876 706718 -3276 706740
rect -3876 706482 -3694 706718
rect -3458 706482 -3276 706718
rect -3876 706398 -3276 706482
rect -3876 706162 -3694 706398
rect -3458 706162 -3276 706398
rect -3876 690054 -3276 706162
rect 4404 706718 5004 707680
rect 4404 706482 4586 706718
rect 4822 706482 5004 706718
rect 4404 706398 5004 706482
rect 4404 706162 4586 706398
rect 4822 706162 5004 706398
rect -3876 689818 -3694 690054
rect -3458 689818 -3276 690054
rect -3876 689734 -3276 689818
rect -3876 689498 -3694 689734
rect -3458 689498 -3276 689734
rect -3876 654054 -3276 689498
rect -3876 653818 -3694 654054
rect -3458 653818 -3276 654054
rect -3876 653734 -3276 653818
rect -3876 653498 -3694 653734
rect -3458 653498 -3276 653734
rect -3876 618054 -3276 653498
rect -3876 617818 -3694 618054
rect -3458 617818 -3276 618054
rect -3876 617734 -3276 617818
rect -3876 617498 -3694 617734
rect -3458 617498 -3276 617734
rect -3876 582054 -3276 617498
rect -3876 581818 -3694 582054
rect -3458 581818 -3276 582054
rect -3876 581734 -3276 581818
rect -3876 581498 -3694 581734
rect -3458 581498 -3276 581734
rect -3876 546054 -3276 581498
rect -3876 545818 -3694 546054
rect -3458 545818 -3276 546054
rect -3876 545734 -3276 545818
rect -3876 545498 -3694 545734
rect -3458 545498 -3276 545734
rect -3876 510054 -3276 545498
rect -3876 509818 -3694 510054
rect -3458 509818 -3276 510054
rect -3876 509734 -3276 509818
rect -3876 509498 -3694 509734
rect -3458 509498 -3276 509734
rect -3876 474054 -3276 509498
rect -3876 473818 -3694 474054
rect -3458 473818 -3276 474054
rect -3876 473734 -3276 473818
rect -3876 473498 -3694 473734
rect -3458 473498 -3276 473734
rect -3876 438054 -3276 473498
rect -3876 437818 -3694 438054
rect -3458 437818 -3276 438054
rect -3876 437734 -3276 437818
rect -3876 437498 -3694 437734
rect -3458 437498 -3276 437734
rect -3876 402054 -3276 437498
rect -3876 401818 -3694 402054
rect -3458 401818 -3276 402054
rect -3876 401734 -3276 401818
rect -3876 401498 -3694 401734
rect -3458 401498 -3276 401734
rect -3876 366054 -3276 401498
rect -3876 365818 -3694 366054
rect -3458 365818 -3276 366054
rect -3876 365734 -3276 365818
rect -3876 365498 -3694 365734
rect -3458 365498 -3276 365734
rect -3876 330054 -3276 365498
rect -3876 329818 -3694 330054
rect -3458 329818 -3276 330054
rect -3876 329734 -3276 329818
rect -3876 329498 -3694 329734
rect -3458 329498 -3276 329734
rect -3876 294054 -3276 329498
rect -3876 293818 -3694 294054
rect -3458 293818 -3276 294054
rect -3876 293734 -3276 293818
rect -3876 293498 -3694 293734
rect -3458 293498 -3276 293734
rect -3876 258054 -3276 293498
rect -3876 257818 -3694 258054
rect -3458 257818 -3276 258054
rect -3876 257734 -3276 257818
rect -3876 257498 -3694 257734
rect -3458 257498 -3276 257734
rect -3876 222054 -3276 257498
rect -3876 221818 -3694 222054
rect -3458 221818 -3276 222054
rect -3876 221734 -3276 221818
rect -3876 221498 -3694 221734
rect -3458 221498 -3276 221734
rect -3876 186054 -3276 221498
rect -3876 185818 -3694 186054
rect -3458 185818 -3276 186054
rect -3876 185734 -3276 185818
rect -3876 185498 -3694 185734
rect -3458 185498 -3276 185734
rect -3876 150054 -3276 185498
rect -3876 149818 -3694 150054
rect -3458 149818 -3276 150054
rect -3876 149734 -3276 149818
rect -3876 149498 -3694 149734
rect -3458 149498 -3276 149734
rect -3876 114054 -3276 149498
rect -3876 113818 -3694 114054
rect -3458 113818 -3276 114054
rect -3876 113734 -3276 113818
rect -3876 113498 -3694 113734
rect -3458 113498 -3276 113734
rect -3876 78054 -3276 113498
rect -3876 77818 -3694 78054
rect -3458 77818 -3276 78054
rect -3876 77734 -3276 77818
rect -3876 77498 -3694 77734
rect -3458 77498 -3276 77734
rect -3876 42054 -3276 77498
rect -3876 41818 -3694 42054
rect -3458 41818 -3276 42054
rect -3876 41734 -3276 41818
rect -3876 41498 -3694 41734
rect -3458 41498 -3276 41734
rect -3876 6054 -3276 41498
rect -3876 5818 -3694 6054
rect -3458 5818 -3276 6054
rect -3876 5734 -3276 5818
rect -3876 5498 -3694 5734
rect -3458 5498 -3276 5734
rect -3876 -2226 -3276 5498
rect -2936 705778 -2336 705800
rect -2936 705542 -2754 705778
rect -2518 705542 -2336 705778
rect -2936 705458 -2336 705542
rect -2936 705222 -2754 705458
rect -2518 705222 -2336 705458
rect -2936 668406 -2336 705222
rect -2936 668170 -2754 668406
rect -2518 668170 -2336 668406
rect -2936 668086 -2336 668170
rect -2936 667850 -2754 668086
rect -2518 667850 -2336 668086
rect -2936 632406 -2336 667850
rect -2936 632170 -2754 632406
rect -2518 632170 -2336 632406
rect -2936 632086 -2336 632170
rect -2936 631850 -2754 632086
rect -2518 631850 -2336 632086
rect -2936 596406 -2336 631850
rect -2936 596170 -2754 596406
rect -2518 596170 -2336 596406
rect -2936 596086 -2336 596170
rect -2936 595850 -2754 596086
rect -2518 595850 -2336 596086
rect -2936 560406 -2336 595850
rect -2936 560170 -2754 560406
rect -2518 560170 -2336 560406
rect -2936 560086 -2336 560170
rect -2936 559850 -2754 560086
rect -2518 559850 -2336 560086
rect -2936 524406 -2336 559850
rect -2936 524170 -2754 524406
rect -2518 524170 -2336 524406
rect -2936 524086 -2336 524170
rect -2936 523850 -2754 524086
rect -2518 523850 -2336 524086
rect -2936 488406 -2336 523850
rect -2936 488170 -2754 488406
rect -2518 488170 -2336 488406
rect -2936 488086 -2336 488170
rect -2936 487850 -2754 488086
rect -2518 487850 -2336 488086
rect -2936 452406 -2336 487850
rect -2936 452170 -2754 452406
rect -2518 452170 -2336 452406
rect -2936 452086 -2336 452170
rect -2936 451850 -2754 452086
rect -2518 451850 -2336 452086
rect -2936 416406 -2336 451850
rect -2936 416170 -2754 416406
rect -2518 416170 -2336 416406
rect -2936 416086 -2336 416170
rect -2936 415850 -2754 416086
rect -2518 415850 -2336 416086
rect -2936 380406 -2336 415850
rect -2936 380170 -2754 380406
rect -2518 380170 -2336 380406
rect -2936 380086 -2336 380170
rect -2936 379850 -2754 380086
rect -2518 379850 -2336 380086
rect -2936 344406 -2336 379850
rect -2936 344170 -2754 344406
rect -2518 344170 -2336 344406
rect -2936 344086 -2336 344170
rect -2936 343850 -2754 344086
rect -2518 343850 -2336 344086
rect -2936 308406 -2336 343850
rect -2936 308170 -2754 308406
rect -2518 308170 -2336 308406
rect -2936 308086 -2336 308170
rect -2936 307850 -2754 308086
rect -2518 307850 -2336 308086
rect -2936 272406 -2336 307850
rect -2936 272170 -2754 272406
rect -2518 272170 -2336 272406
rect -2936 272086 -2336 272170
rect -2936 271850 -2754 272086
rect -2518 271850 -2336 272086
rect -2936 236406 -2336 271850
rect -2936 236170 -2754 236406
rect -2518 236170 -2336 236406
rect -2936 236086 -2336 236170
rect -2936 235850 -2754 236086
rect -2518 235850 -2336 236086
rect -2936 200406 -2336 235850
rect -2936 200170 -2754 200406
rect -2518 200170 -2336 200406
rect -2936 200086 -2336 200170
rect -2936 199850 -2754 200086
rect -2518 199850 -2336 200086
rect -2936 164406 -2336 199850
rect -2936 164170 -2754 164406
rect -2518 164170 -2336 164406
rect -2936 164086 -2336 164170
rect -2936 163850 -2754 164086
rect -2518 163850 -2336 164086
rect -2936 128406 -2336 163850
rect -2936 128170 -2754 128406
rect -2518 128170 -2336 128406
rect -2936 128086 -2336 128170
rect -2936 127850 -2754 128086
rect -2518 127850 -2336 128086
rect -2936 92406 -2336 127850
rect -2936 92170 -2754 92406
rect -2518 92170 -2336 92406
rect -2936 92086 -2336 92170
rect -2936 91850 -2754 92086
rect -2518 91850 -2336 92086
rect -2936 56406 -2336 91850
rect -2936 56170 -2754 56406
rect -2518 56170 -2336 56406
rect -2936 56086 -2336 56170
rect -2936 55850 -2754 56086
rect -2518 55850 -2336 56086
rect -2936 20406 -2336 55850
rect -2936 20170 -2754 20406
rect -2518 20170 -2336 20406
rect -2936 20086 -2336 20170
rect -2936 19850 -2754 20086
rect -2518 19850 -2336 20086
rect -2936 -1286 -2336 19850
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686406 -1396 704282
rect -1996 686170 -1814 686406
rect -1578 686170 -1396 686406
rect -1996 686086 -1396 686170
rect -1996 685850 -1814 686086
rect -1578 685850 -1396 686086
rect -1996 650406 -1396 685850
rect -1996 650170 -1814 650406
rect -1578 650170 -1396 650406
rect -1996 650086 -1396 650170
rect -1996 649850 -1814 650086
rect -1578 649850 -1396 650086
rect -1996 614406 -1396 649850
rect -1996 614170 -1814 614406
rect -1578 614170 -1396 614406
rect -1996 614086 -1396 614170
rect -1996 613850 -1814 614086
rect -1578 613850 -1396 614086
rect -1996 578406 -1396 613850
rect -1996 578170 -1814 578406
rect -1578 578170 -1396 578406
rect -1996 578086 -1396 578170
rect -1996 577850 -1814 578086
rect -1578 577850 -1396 578086
rect -1996 542406 -1396 577850
rect -1996 542170 -1814 542406
rect -1578 542170 -1396 542406
rect -1996 542086 -1396 542170
rect -1996 541850 -1814 542086
rect -1578 541850 -1396 542086
rect -1996 506406 -1396 541850
rect -1996 506170 -1814 506406
rect -1578 506170 -1396 506406
rect -1996 506086 -1396 506170
rect -1996 505850 -1814 506086
rect -1578 505850 -1396 506086
rect -1996 470406 -1396 505850
rect -1996 470170 -1814 470406
rect -1578 470170 -1396 470406
rect -1996 470086 -1396 470170
rect -1996 469850 -1814 470086
rect -1578 469850 -1396 470086
rect -1996 434406 -1396 469850
rect -1996 434170 -1814 434406
rect -1578 434170 -1396 434406
rect -1996 434086 -1396 434170
rect -1996 433850 -1814 434086
rect -1578 433850 -1396 434086
rect -1996 398406 -1396 433850
rect -1996 398170 -1814 398406
rect -1578 398170 -1396 398406
rect -1996 398086 -1396 398170
rect -1996 397850 -1814 398086
rect -1578 397850 -1396 398086
rect -1996 362406 -1396 397850
rect -1996 362170 -1814 362406
rect -1578 362170 -1396 362406
rect -1996 362086 -1396 362170
rect -1996 361850 -1814 362086
rect -1578 361850 -1396 362086
rect -1996 326406 -1396 361850
rect -1996 326170 -1814 326406
rect -1578 326170 -1396 326406
rect -1996 326086 -1396 326170
rect -1996 325850 -1814 326086
rect -1578 325850 -1396 326086
rect -1996 290406 -1396 325850
rect -1996 290170 -1814 290406
rect -1578 290170 -1396 290406
rect -1996 290086 -1396 290170
rect -1996 289850 -1814 290086
rect -1578 289850 -1396 290086
rect -1996 254406 -1396 289850
rect -1996 254170 -1814 254406
rect -1578 254170 -1396 254406
rect -1996 254086 -1396 254170
rect -1996 253850 -1814 254086
rect -1578 253850 -1396 254086
rect -1996 218406 -1396 253850
rect -1996 218170 -1814 218406
rect -1578 218170 -1396 218406
rect -1996 218086 -1396 218170
rect -1996 217850 -1814 218086
rect -1578 217850 -1396 218086
rect -1996 182406 -1396 217850
rect -1996 182170 -1814 182406
rect -1578 182170 -1396 182406
rect -1996 182086 -1396 182170
rect -1996 181850 -1814 182086
rect -1578 181850 -1396 182086
rect -1996 146406 -1396 181850
rect -1996 146170 -1814 146406
rect -1578 146170 -1396 146406
rect -1996 146086 -1396 146170
rect -1996 145850 -1814 146086
rect -1578 145850 -1396 146086
rect -1996 110406 -1396 145850
rect -1996 110170 -1814 110406
rect -1578 110170 -1396 110406
rect -1996 110086 -1396 110170
rect -1996 109850 -1814 110086
rect -1578 109850 -1396 110086
rect -1996 74406 -1396 109850
rect -1996 74170 -1814 74406
rect -1578 74170 -1396 74406
rect -1996 74086 -1396 74170
rect -1996 73850 -1814 74086
rect -1578 73850 -1396 74086
rect -1996 38406 -1396 73850
rect -1996 38170 -1814 38406
rect -1578 38170 -1396 38406
rect -1996 38086 -1396 38170
rect -1996 37850 -1814 38086
rect -1578 37850 -1396 38086
rect -1996 2406 -1396 37850
rect -1996 2170 -1814 2406
rect -1578 2170 -1396 2406
rect -1996 2086 -1396 2170
rect -1996 1850 -1814 2086
rect -1578 1850 -1396 2086
rect -1996 -346 -1396 1850
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705800
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686406 1404 704282
rect 804 686170 986 686406
rect 1222 686170 1404 686406
rect 804 686086 1404 686170
rect 804 685850 986 686086
rect 1222 685850 1404 686086
rect 804 650406 1404 685850
rect 804 650170 986 650406
rect 1222 650170 1404 650406
rect 804 650086 1404 650170
rect 804 649850 986 650086
rect 1222 649850 1404 650086
rect 804 614406 1404 649850
rect 804 614170 986 614406
rect 1222 614170 1404 614406
rect 804 614086 1404 614170
rect 804 613850 986 614086
rect 1222 613850 1404 614086
rect 804 578406 1404 613850
rect 804 578170 986 578406
rect 1222 578170 1404 578406
rect 804 578086 1404 578170
rect 804 577850 986 578086
rect 1222 577850 1404 578086
rect 804 542406 1404 577850
rect 804 542170 986 542406
rect 1222 542170 1404 542406
rect 804 542086 1404 542170
rect 804 541850 986 542086
rect 1222 541850 1404 542086
rect 804 506406 1404 541850
rect 804 506170 986 506406
rect 1222 506170 1404 506406
rect 804 506086 1404 506170
rect 804 505850 986 506086
rect 1222 505850 1404 506086
rect 804 470406 1404 505850
rect 804 470170 986 470406
rect 1222 470170 1404 470406
rect 804 470086 1404 470170
rect 804 469850 986 470086
rect 1222 469850 1404 470086
rect 804 434406 1404 469850
rect 804 434170 986 434406
rect 1222 434170 1404 434406
rect 804 434086 1404 434170
rect 804 433850 986 434086
rect 1222 433850 1404 434086
rect 804 398406 1404 433850
rect 804 398170 986 398406
rect 1222 398170 1404 398406
rect 804 398086 1404 398170
rect 804 397850 986 398086
rect 1222 397850 1404 398086
rect 804 362406 1404 397850
rect 804 362170 986 362406
rect 1222 362170 1404 362406
rect 804 362086 1404 362170
rect 804 361850 986 362086
rect 1222 361850 1404 362086
rect 804 326406 1404 361850
rect 804 326170 986 326406
rect 1222 326170 1404 326406
rect 804 326086 1404 326170
rect 804 325850 986 326086
rect 1222 325850 1404 326086
rect 804 290406 1404 325850
rect 804 290170 986 290406
rect 1222 290170 1404 290406
rect 804 290086 1404 290170
rect 804 289850 986 290086
rect 1222 289850 1404 290086
rect 804 254406 1404 289850
rect 804 254170 986 254406
rect 1222 254170 1404 254406
rect 804 254086 1404 254170
rect 804 253850 986 254086
rect 1222 253850 1404 254086
rect 804 218406 1404 253850
rect 804 218170 986 218406
rect 1222 218170 1404 218406
rect 804 218086 1404 218170
rect 804 217850 986 218086
rect 1222 217850 1404 218086
rect 804 182406 1404 217850
rect 804 182170 986 182406
rect 1222 182170 1404 182406
rect 804 182086 1404 182170
rect 804 181850 986 182086
rect 1222 181850 1404 182086
rect 804 146406 1404 181850
rect 804 146170 986 146406
rect 1222 146170 1404 146406
rect 804 146086 1404 146170
rect 804 145850 986 146086
rect 1222 145850 1404 146086
rect 804 110406 1404 145850
rect 804 110170 986 110406
rect 1222 110170 1404 110406
rect 804 110086 1404 110170
rect 804 109850 986 110086
rect 1222 109850 1404 110086
rect 804 74406 1404 109850
rect 804 74170 986 74406
rect 1222 74170 1404 74406
rect 804 74086 1404 74170
rect 804 73850 986 74086
rect 1222 73850 1404 74086
rect 804 38406 1404 73850
rect 804 38170 986 38406
rect 1222 38170 1404 38406
rect 804 38086 1404 38170
rect 804 37850 986 38086
rect 1222 37850 1404 38086
rect 804 2406 1404 37850
rect 804 2170 986 2406
rect 1222 2170 1404 2406
rect 804 2086 1404 2170
rect 804 1850 986 2086
rect 1222 1850 1404 2086
rect 804 -346 1404 1850
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2936 -1522 -2754 -1286
rect -2518 -1522 -2336 -1286
rect -2936 -1606 -2336 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 -2336 -1606
rect -2936 -1864 -2336 -1842
rect 804 -1864 1404 -902
rect 4404 690054 5004 706162
rect 8004 698000 8604 708042
rect 11604 698000 12204 709922
rect 29604 711418 30204 711440
rect 29604 711182 29786 711418
rect 30022 711182 30204 711418
rect 29604 711098 30204 711182
rect 29604 710862 29786 711098
rect 30022 710862 30204 711098
rect 26004 709538 26604 709560
rect 26004 709302 26186 709538
rect 26422 709302 26604 709538
rect 26004 709218 26604 709302
rect 26004 708982 26186 709218
rect 26422 708982 26604 709218
rect 22404 707658 23004 707680
rect 22404 707422 22586 707658
rect 22822 707422 23004 707658
rect 22404 707338 23004 707422
rect 22404 707102 22586 707338
rect 22822 707102 23004 707338
rect 18804 705778 19404 705800
rect 18804 705542 18986 705778
rect 19222 705542 19404 705778
rect 18804 705458 19404 705542
rect 18804 705222 18986 705458
rect 19222 705222 19404 705458
rect 18804 701248 19404 705222
rect 18804 701184 18832 701248
rect 18896 701184 18912 701248
rect 18976 701184 18992 701248
rect 19056 701184 19072 701248
rect 19136 701184 19152 701248
rect 19216 701184 19232 701248
rect 19296 701184 19312 701248
rect 19376 701184 19404 701248
rect 18804 700160 19404 701184
rect 18804 700096 18832 700160
rect 18896 700096 18912 700160
rect 18976 700096 18992 700160
rect 19056 700096 19072 700160
rect 19136 700096 19152 700160
rect 19216 700096 19232 700160
rect 19296 700096 19312 700160
rect 19376 700096 19404 700160
rect 18804 699072 19404 700096
rect 18804 699008 18832 699072
rect 18896 699008 18912 699072
rect 18976 699008 18992 699072
rect 19056 699008 19072 699072
rect 19136 699008 19152 699072
rect 19216 699008 19232 699072
rect 19296 699008 19312 699072
rect 19376 699008 19404 699072
rect 18804 697952 19404 699008
rect 22404 698000 23004 707102
rect 26004 698000 26604 708982
rect 29604 698000 30204 710862
rect 47604 710478 48204 711440
rect 47604 710242 47786 710478
rect 48022 710242 48204 710478
rect 47604 710158 48204 710242
rect 47604 709922 47786 710158
rect 48022 709922 48204 710158
rect 44004 708598 44604 709560
rect 44004 708362 44186 708598
rect 44422 708362 44604 708598
rect 44004 708278 44604 708362
rect 44004 708042 44186 708278
rect 44422 708042 44604 708278
rect 40404 706718 41004 707680
rect 40404 706482 40586 706718
rect 40822 706482 41004 706718
rect 40404 706398 41004 706482
rect 40404 706162 40586 706398
rect 40822 706162 41004 706398
rect 36804 704838 37404 705800
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 701792 37404 704282
rect 36804 701728 36832 701792
rect 36896 701728 36912 701792
rect 36976 701728 36992 701792
rect 37056 701728 37072 701792
rect 37136 701728 37152 701792
rect 37216 701728 37232 701792
rect 37296 701728 37312 701792
rect 37376 701728 37404 701792
rect 36804 700704 37404 701728
rect 36804 700640 36832 700704
rect 36896 700640 36912 700704
rect 36976 700640 36992 700704
rect 37056 700640 37072 700704
rect 37136 700640 37152 700704
rect 37216 700640 37232 700704
rect 37296 700640 37312 700704
rect 37376 700640 37404 700704
rect 36804 699616 37404 700640
rect 36804 699552 36832 699616
rect 36896 699552 36912 699616
rect 36976 699552 36992 699616
rect 37056 699552 37072 699616
rect 37136 699552 37152 699616
rect 37216 699552 37232 699616
rect 37296 699552 37312 699616
rect 37376 699552 37404 699616
rect 36804 698528 37404 699552
rect 36804 698464 36832 698528
rect 36896 698464 36912 698528
rect 36976 698464 36992 698528
rect 37056 698464 37072 698528
rect 37136 698464 37152 698528
rect 37216 698464 37232 698528
rect 37296 698464 37312 698528
rect 37376 698464 37404 698528
rect 36804 697952 37404 698464
rect 40404 698000 41004 706162
rect 44004 698000 44604 708042
rect 47604 698000 48204 709922
rect 65604 711418 66204 711440
rect 65604 711182 65786 711418
rect 66022 711182 66204 711418
rect 65604 711098 66204 711182
rect 65604 710862 65786 711098
rect 66022 710862 66204 711098
rect 62004 709538 62604 709560
rect 62004 709302 62186 709538
rect 62422 709302 62604 709538
rect 62004 709218 62604 709302
rect 62004 708982 62186 709218
rect 62422 708982 62604 709218
rect 58404 707658 59004 707680
rect 58404 707422 58586 707658
rect 58822 707422 59004 707658
rect 58404 707338 59004 707422
rect 58404 707102 58586 707338
rect 58822 707102 59004 707338
rect 54804 705778 55404 705800
rect 54804 705542 54986 705778
rect 55222 705542 55404 705778
rect 54804 705458 55404 705542
rect 54804 705222 54986 705458
rect 55222 705222 55404 705458
rect 54804 701248 55404 705222
rect 54804 701184 54832 701248
rect 54896 701184 54912 701248
rect 54976 701184 54992 701248
rect 55056 701184 55072 701248
rect 55136 701184 55152 701248
rect 55216 701184 55232 701248
rect 55296 701184 55312 701248
rect 55376 701184 55404 701248
rect 54804 700160 55404 701184
rect 54804 700096 54832 700160
rect 54896 700096 54912 700160
rect 54976 700096 54992 700160
rect 55056 700096 55072 700160
rect 55136 700096 55152 700160
rect 55216 700096 55232 700160
rect 55296 700096 55312 700160
rect 55376 700096 55404 700160
rect 54804 699072 55404 700096
rect 54804 699008 54832 699072
rect 54896 699008 54912 699072
rect 54976 699008 54992 699072
rect 55056 699008 55072 699072
rect 55136 699008 55152 699072
rect 55216 699008 55232 699072
rect 55296 699008 55312 699072
rect 55376 699008 55404 699072
rect 54804 697952 55404 699008
rect 58404 698000 59004 707102
rect 62004 698000 62604 708982
rect 65604 698000 66204 710862
rect 83604 710478 84204 711440
rect 83604 710242 83786 710478
rect 84022 710242 84204 710478
rect 83604 710158 84204 710242
rect 83604 709922 83786 710158
rect 84022 709922 84204 710158
rect 80004 708598 80604 709560
rect 80004 708362 80186 708598
rect 80422 708362 80604 708598
rect 80004 708278 80604 708362
rect 80004 708042 80186 708278
rect 80422 708042 80604 708278
rect 76404 706718 77004 707680
rect 76404 706482 76586 706718
rect 76822 706482 77004 706718
rect 76404 706398 77004 706482
rect 76404 706162 76586 706398
rect 76822 706162 77004 706398
rect 72804 704838 73404 705800
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 701792 73404 704282
rect 72804 701728 72832 701792
rect 72896 701728 72912 701792
rect 72976 701728 72992 701792
rect 73056 701728 73072 701792
rect 73136 701728 73152 701792
rect 73216 701728 73232 701792
rect 73296 701728 73312 701792
rect 73376 701728 73404 701792
rect 72804 700704 73404 701728
rect 72804 700640 72832 700704
rect 72896 700640 72912 700704
rect 72976 700640 72992 700704
rect 73056 700640 73072 700704
rect 73136 700640 73152 700704
rect 73216 700640 73232 700704
rect 73296 700640 73312 700704
rect 73376 700640 73404 700704
rect 72804 699616 73404 700640
rect 72804 699552 72832 699616
rect 72896 699552 72912 699616
rect 72976 699552 72992 699616
rect 73056 699552 73072 699616
rect 73136 699552 73152 699616
rect 73216 699552 73232 699616
rect 73296 699552 73312 699616
rect 73376 699552 73404 699616
rect 72804 698528 73404 699552
rect 72804 698464 72832 698528
rect 72896 698464 72912 698528
rect 72976 698464 72992 698528
rect 73056 698464 73072 698528
rect 73136 698464 73152 698528
rect 73216 698464 73232 698528
rect 73296 698464 73312 698528
rect 73376 698464 73404 698528
rect 72804 697952 73404 698464
rect 76404 698000 77004 706162
rect 80004 698000 80604 708042
rect 83604 698000 84204 709922
rect 101604 711418 102204 711440
rect 101604 711182 101786 711418
rect 102022 711182 102204 711418
rect 101604 711098 102204 711182
rect 101604 710862 101786 711098
rect 102022 710862 102204 711098
rect 98004 709538 98604 709560
rect 98004 709302 98186 709538
rect 98422 709302 98604 709538
rect 98004 709218 98604 709302
rect 98004 708982 98186 709218
rect 98422 708982 98604 709218
rect 94404 707658 95004 707680
rect 94404 707422 94586 707658
rect 94822 707422 95004 707658
rect 94404 707338 95004 707422
rect 94404 707102 94586 707338
rect 94822 707102 95004 707338
rect 90804 705778 91404 705800
rect 90804 705542 90986 705778
rect 91222 705542 91404 705778
rect 90804 705458 91404 705542
rect 90804 705222 90986 705458
rect 91222 705222 91404 705458
rect 90804 701248 91404 705222
rect 90804 701184 90832 701248
rect 90896 701184 90912 701248
rect 90976 701184 90992 701248
rect 91056 701184 91072 701248
rect 91136 701184 91152 701248
rect 91216 701184 91232 701248
rect 91296 701184 91312 701248
rect 91376 701184 91404 701248
rect 90804 700160 91404 701184
rect 90804 700096 90832 700160
rect 90896 700096 90912 700160
rect 90976 700096 90992 700160
rect 91056 700096 91072 700160
rect 91136 700096 91152 700160
rect 91216 700096 91232 700160
rect 91296 700096 91312 700160
rect 91376 700096 91404 700160
rect 90804 699072 91404 700096
rect 90804 699008 90832 699072
rect 90896 699008 90912 699072
rect 90976 699008 90992 699072
rect 91056 699008 91072 699072
rect 91136 699008 91152 699072
rect 91216 699008 91232 699072
rect 91296 699008 91312 699072
rect 91376 699008 91404 699072
rect 90804 697952 91404 699008
rect 94404 698000 95004 707102
rect 98004 698000 98604 708982
rect 101604 698000 102204 710862
rect 119604 710478 120204 711440
rect 119604 710242 119786 710478
rect 120022 710242 120204 710478
rect 119604 710158 120204 710242
rect 119604 709922 119786 710158
rect 120022 709922 120204 710158
rect 116004 708598 116604 709560
rect 116004 708362 116186 708598
rect 116422 708362 116604 708598
rect 116004 708278 116604 708362
rect 116004 708042 116186 708278
rect 116422 708042 116604 708278
rect 112404 706718 113004 707680
rect 112404 706482 112586 706718
rect 112822 706482 113004 706718
rect 112404 706398 113004 706482
rect 112404 706162 112586 706398
rect 112822 706162 113004 706398
rect 108804 704838 109404 705800
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 701792 109404 704282
rect 108804 701728 108832 701792
rect 108896 701728 108912 701792
rect 108976 701728 108992 701792
rect 109056 701728 109072 701792
rect 109136 701728 109152 701792
rect 109216 701728 109232 701792
rect 109296 701728 109312 701792
rect 109376 701728 109404 701792
rect 108804 700704 109404 701728
rect 108804 700640 108832 700704
rect 108896 700640 108912 700704
rect 108976 700640 108992 700704
rect 109056 700640 109072 700704
rect 109136 700640 109152 700704
rect 109216 700640 109232 700704
rect 109296 700640 109312 700704
rect 109376 700640 109404 700704
rect 108804 699616 109404 700640
rect 108804 699552 108832 699616
rect 108896 699552 108912 699616
rect 108976 699552 108992 699616
rect 109056 699552 109072 699616
rect 109136 699552 109152 699616
rect 109216 699552 109232 699616
rect 109296 699552 109312 699616
rect 109376 699552 109404 699616
rect 108804 698528 109404 699552
rect 108804 698464 108832 698528
rect 108896 698464 108912 698528
rect 108976 698464 108992 698528
rect 109056 698464 109072 698528
rect 109136 698464 109152 698528
rect 109216 698464 109232 698528
rect 109296 698464 109312 698528
rect 109376 698464 109404 698528
rect 108804 697952 109404 698464
rect 112404 698000 113004 706162
rect 116004 698000 116604 708042
rect 119604 698000 120204 709922
rect 137604 711418 138204 711440
rect 137604 711182 137786 711418
rect 138022 711182 138204 711418
rect 137604 711098 138204 711182
rect 137604 710862 137786 711098
rect 138022 710862 138204 711098
rect 134004 709538 134604 709560
rect 134004 709302 134186 709538
rect 134422 709302 134604 709538
rect 134004 709218 134604 709302
rect 134004 708982 134186 709218
rect 134422 708982 134604 709218
rect 130404 707658 131004 707680
rect 130404 707422 130586 707658
rect 130822 707422 131004 707658
rect 130404 707338 131004 707422
rect 130404 707102 130586 707338
rect 130822 707102 131004 707338
rect 126804 705778 127404 705800
rect 126804 705542 126986 705778
rect 127222 705542 127404 705778
rect 126804 705458 127404 705542
rect 126804 705222 126986 705458
rect 127222 705222 127404 705458
rect 126804 701248 127404 705222
rect 126804 701184 126832 701248
rect 126896 701184 126912 701248
rect 126976 701184 126992 701248
rect 127056 701184 127072 701248
rect 127136 701184 127152 701248
rect 127216 701184 127232 701248
rect 127296 701184 127312 701248
rect 127376 701184 127404 701248
rect 126804 700160 127404 701184
rect 126804 700096 126832 700160
rect 126896 700096 126912 700160
rect 126976 700096 126992 700160
rect 127056 700096 127072 700160
rect 127136 700096 127152 700160
rect 127216 700096 127232 700160
rect 127296 700096 127312 700160
rect 127376 700096 127404 700160
rect 126804 699072 127404 700096
rect 126804 699008 126832 699072
rect 126896 699008 126912 699072
rect 126976 699008 126992 699072
rect 127056 699008 127072 699072
rect 127136 699008 127152 699072
rect 127216 699008 127232 699072
rect 127296 699008 127312 699072
rect 127376 699008 127404 699072
rect 126804 697952 127404 699008
rect 130404 698000 131004 707102
rect 134004 698000 134604 708982
rect 137604 698000 138204 710862
rect 155604 710478 156204 711440
rect 155604 710242 155786 710478
rect 156022 710242 156204 710478
rect 155604 710158 156204 710242
rect 155604 709922 155786 710158
rect 156022 709922 156204 710158
rect 152004 708598 152604 709560
rect 152004 708362 152186 708598
rect 152422 708362 152604 708598
rect 152004 708278 152604 708362
rect 152004 708042 152186 708278
rect 152422 708042 152604 708278
rect 148404 706718 149004 707680
rect 148404 706482 148586 706718
rect 148822 706482 149004 706718
rect 148404 706398 149004 706482
rect 148404 706162 148586 706398
rect 148822 706162 149004 706398
rect 144804 704838 145404 705800
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 701792 145404 704282
rect 144804 701728 144832 701792
rect 144896 701728 144912 701792
rect 144976 701728 144992 701792
rect 145056 701728 145072 701792
rect 145136 701728 145152 701792
rect 145216 701728 145232 701792
rect 145296 701728 145312 701792
rect 145376 701728 145404 701792
rect 144804 700704 145404 701728
rect 144804 700640 144832 700704
rect 144896 700640 144912 700704
rect 144976 700640 144992 700704
rect 145056 700640 145072 700704
rect 145136 700640 145152 700704
rect 145216 700640 145232 700704
rect 145296 700640 145312 700704
rect 145376 700640 145404 700704
rect 144804 699616 145404 700640
rect 144804 699552 144832 699616
rect 144896 699552 144912 699616
rect 144976 699552 144992 699616
rect 145056 699552 145072 699616
rect 145136 699552 145152 699616
rect 145216 699552 145232 699616
rect 145296 699552 145312 699616
rect 145376 699552 145404 699616
rect 144804 698528 145404 699552
rect 144804 698464 144832 698528
rect 144896 698464 144912 698528
rect 144976 698464 144992 698528
rect 145056 698464 145072 698528
rect 145136 698464 145152 698528
rect 145216 698464 145232 698528
rect 145296 698464 145312 698528
rect 145376 698464 145404 698528
rect 144804 697952 145404 698464
rect 148404 698000 149004 706162
rect 152004 698000 152604 708042
rect 155604 698000 156204 709922
rect 173604 711418 174204 711440
rect 173604 711182 173786 711418
rect 174022 711182 174204 711418
rect 173604 711098 174204 711182
rect 173604 710862 173786 711098
rect 174022 710862 174204 711098
rect 170004 709538 170604 709560
rect 170004 709302 170186 709538
rect 170422 709302 170604 709538
rect 170004 709218 170604 709302
rect 170004 708982 170186 709218
rect 170422 708982 170604 709218
rect 166404 707658 167004 707680
rect 166404 707422 166586 707658
rect 166822 707422 167004 707658
rect 166404 707338 167004 707422
rect 166404 707102 166586 707338
rect 166822 707102 167004 707338
rect 162804 705778 163404 705800
rect 162804 705542 162986 705778
rect 163222 705542 163404 705778
rect 162804 705458 163404 705542
rect 162804 705222 162986 705458
rect 163222 705222 163404 705458
rect 162804 701248 163404 705222
rect 162804 701184 162832 701248
rect 162896 701184 162912 701248
rect 162976 701184 162992 701248
rect 163056 701184 163072 701248
rect 163136 701184 163152 701248
rect 163216 701184 163232 701248
rect 163296 701184 163312 701248
rect 163376 701184 163404 701248
rect 162804 700160 163404 701184
rect 162804 700096 162832 700160
rect 162896 700096 162912 700160
rect 162976 700096 162992 700160
rect 163056 700096 163072 700160
rect 163136 700096 163152 700160
rect 163216 700096 163232 700160
rect 163296 700096 163312 700160
rect 163376 700096 163404 700160
rect 162804 699072 163404 700096
rect 162804 699008 162832 699072
rect 162896 699008 162912 699072
rect 162976 699008 162992 699072
rect 163056 699008 163072 699072
rect 163136 699008 163152 699072
rect 163216 699008 163232 699072
rect 163296 699008 163312 699072
rect 163376 699008 163404 699072
rect 162804 697952 163404 699008
rect 166404 698000 167004 707102
rect 170004 698000 170604 708982
rect 173604 698000 174204 710862
rect 191604 710478 192204 711440
rect 191604 710242 191786 710478
rect 192022 710242 192204 710478
rect 191604 710158 192204 710242
rect 191604 709922 191786 710158
rect 192022 709922 192204 710158
rect 188004 708598 188604 709560
rect 188004 708362 188186 708598
rect 188422 708362 188604 708598
rect 188004 708278 188604 708362
rect 188004 708042 188186 708278
rect 188422 708042 188604 708278
rect 184404 706718 185004 707680
rect 184404 706482 184586 706718
rect 184822 706482 185004 706718
rect 184404 706398 185004 706482
rect 184404 706162 184586 706398
rect 184822 706162 185004 706398
rect 180804 704838 181404 705800
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 701792 181404 704282
rect 180804 701728 180832 701792
rect 180896 701728 180912 701792
rect 180976 701728 180992 701792
rect 181056 701728 181072 701792
rect 181136 701728 181152 701792
rect 181216 701728 181232 701792
rect 181296 701728 181312 701792
rect 181376 701728 181404 701792
rect 180804 700704 181404 701728
rect 180804 700640 180832 700704
rect 180896 700640 180912 700704
rect 180976 700640 180992 700704
rect 181056 700640 181072 700704
rect 181136 700640 181152 700704
rect 181216 700640 181232 700704
rect 181296 700640 181312 700704
rect 181376 700640 181404 700704
rect 180804 699616 181404 700640
rect 180804 699552 180832 699616
rect 180896 699552 180912 699616
rect 180976 699552 180992 699616
rect 181056 699552 181072 699616
rect 181136 699552 181152 699616
rect 181216 699552 181232 699616
rect 181296 699552 181312 699616
rect 181376 699552 181404 699616
rect 180804 698528 181404 699552
rect 180804 698464 180832 698528
rect 180896 698464 180912 698528
rect 180976 698464 180992 698528
rect 181056 698464 181072 698528
rect 181136 698464 181152 698528
rect 181216 698464 181232 698528
rect 181296 698464 181312 698528
rect 181376 698464 181404 698528
rect 180804 697952 181404 698464
rect 184404 698000 185004 706162
rect 188004 698000 188604 708042
rect 191604 698000 192204 709922
rect 209604 711418 210204 711440
rect 209604 711182 209786 711418
rect 210022 711182 210204 711418
rect 209604 711098 210204 711182
rect 209604 710862 209786 711098
rect 210022 710862 210204 711098
rect 206004 709538 206604 709560
rect 206004 709302 206186 709538
rect 206422 709302 206604 709538
rect 206004 709218 206604 709302
rect 206004 708982 206186 709218
rect 206422 708982 206604 709218
rect 202404 707658 203004 707680
rect 202404 707422 202586 707658
rect 202822 707422 203004 707658
rect 202404 707338 203004 707422
rect 202404 707102 202586 707338
rect 202822 707102 203004 707338
rect 198804 705778 199404 705800
rect 198804 705542 198986 705778
rect 199222 705542 199404 705778
rect 198804 705458 199404 705542
rect 198804 705222 198986 705458
rect 199222 705222 199404 705458
rect 198804 701248 199404 705222
rect 198804 701184 198832 701248
rect 198896 701184 198912 701248
rect 198976 701184 198992 701248
rect 199056 701184 199072 701248
rect 199136 701184 199152 701248
rect 199216 701184 199232 701248
rect 199296 701184 199312 701248
rect 199376 701184 199404 701248
rect 198804 700160 199404 701184
rect 198804 700096 198832 700160
rect 198896 700096 198912 700160
rect 198976 700096 198992 700160
rect 199056 700096 199072 700160
rect 199136 700096 199152 700160
rect 199216 700096 199232 700160
rect 199296 700096 199312 700160
rect 199376 700096 199404 700160
rect 198804 699072 199404 700096
rect 198804 699008 198832 699072
rect 198896 699008 198912 699072
rect 198976 699008 198992 699072
rect 199056 699008 199072 699072
rect 199136 699008 199152 699072
rect 199216 699008 199232 699072
rect 199296 699008 199312 699072
rect 199376 699008 199404 699072
rect 198804 697952 199404 699008
rect 202404 698000 203004 707102
rect 206004 698000 206604 708982
rect 209604 698000 210204 710862
rect 227604 710478 228204 711440
rect 227604 710242 227786 710478
rect 228022 710242 228204 710478
rect 227604 710158 228204 710242
rect 227604 709922 227786 710158
rect 228022 709922 228204 710158
rect 224004 708598 224604 709560
rect 224004 708362 224186 708598
rect 224422 708362 224604 708598
rect 224004 708278 224604 708362
rect 224004 708042 224186 708278
rect 224422 708042 224604 708278
rect 220404 706718 221004 707680
rect 220404 706482 220586 706718
rect 220822 706482 221004 706718
rect 220404 706398 221004 706482
rect 220404 706162 220586 706398
rect 220822 706162 221004 706398
rect 216804 704838 217404 705800
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 701792 217404 704282
rect 216804 701728 216832 701792
rect 216896 701728 216912 701792
rect 216976 701728 216992 701792
rect 217056 701728 217072 701792
rect 217136 701728 217152 701792
rect 217216 701728 217232 701792
rect 217296 701728 217312 701792
rect 217376 701728 217404 701792
rect 216804 700704 217404 701728
rect 216804 700640 216832 700704
rect 216896 700640 216912 700704
rect 216976 700640 216992 700704
rect 217056 700640 217072 700704
rect 217136 700640 217152 700704
rect 217216 700640 217232 700704
rect 217296 700640 217312 700704
rect 217376 700640 217404 700704
rect 216804 699616 217404 700640
rect 216804 699552 216832 699616
rect 216896 699552 216912 699616
rect 216976 699552 216992 699616
rect 217056 699552 217072 699616
rect 217136 699552 217152 699616
rect 217216 699552 217232 699616
rect 217296 699552 217312 699616
rect 217376 699552 217404 699616
rect 216804 698528 217404 699552
rect 216804 698464 216832 698528
rect 216896 698464 216912 698528
rect 216976 698464 216992 698528
rect 217056 698464 217072 698528
rect 217136 698464 217152 698528
rect 217216 698464 217232 698528
rect 217296 698464 217312 698528
rect 217376 698464 217404 698528
rect 216804 697952 217404 698464
rect 220404 698000 221004 706162
rect 224004 698000 224604 708042
rect 227604 698000 228204 709922
rect 245604 711418 246204 711440
rect 245604 711182 245786 711418
rect 246022 711182 246204 711418
rect 245604 711098 246204 711182
rect 245604 710862 245786 711098
rect 246022 710862 246204 711098
rect 242004 709538 242604 709560
rect 242004 709302 242186 709538
rect 242422 709302 242604 709538
rect 242004 709218 242604 709302
rect 242004 708982 242186 709218
rect 242422 708982 242604 709218
rect 238404 707658 239004 707680
rect 238404 707422 238586 707658
rect 238822 707422 239004 707658
rect 238404 707338 239004 707422
rect 238404 707102 238586 707338
rect 238822 707102 239004 707338
rect 234804 705778 235404 705800
rect 234804 705542 234986 705778
rect 235222 705542 235404 705778
rect 234804 705458 235404 705542
rect 234804 705222 234986 705458
rect 235222 705222 235404 705458
rect 234804 701248 235404 705222
rect 234804 701184 234832 701248
rect 234896 701184 234912 701248
rect 234976 701184 234992 701248
rect 235056 701184 235072 701248
rect 235136 701184 235152 701248
rect 235216 701184 235232 701248
rect 235296 701184 235312 701248
rect 235376 701184 235404 701248
rect 234804 700160 235404 701184
rect 234804 700096 234832 700160
rect 234896 700096 234912 700160
rect 234976 700096 234992 700160
rect 235056 700096 235072 700160
rect 235136 700096 235152 700160
rect 235216 700096 235232 700160
rect 235296 700096 235312 700160
rect 235376 700096 235404 700160
rect 234804 699072 235404 700096
rect 234804 699008 234832 699072
rect 234896 699008 234912 699072
rect 234976 699008 234992 699072
rect 235056 699008 235072 699072
rect 235136 699008 235152 699072
rect 235216 699008 235232 699072
rect 235296 699008 235312 699072
rect 235376 699008 235404 699072
rect 234804 697952 235404 699008
rect 238404 698000 239004 707102
rect 242004 698000 242604 708982
rect 245604 698000 246204 710862
rect 263604 710478 264204 711440
rect 263604 710242 263786 710478
rect 264022 710242 264204 710478
rect 263604 710158 264204 710242
rect 263604 709922 263786 710158
rect 264022 709922 264204 710158
rect 260004 708598 260604 709560
rect 260004 708362 260186 708598
rect 260422 708362 260604 708598
rect 260004 708278 260604 708362
rect 260004 708042 260186 708278
rect 260422 708042 260604 708278
rect 256404 706718 257004 707680
rect 256404 706482 256586 706718
rect 256822 706482 257004 706718
rect 256404 706398 257004 706482
rect 256404 706162 256586 706398
rect 256822 706162 257004 706398
rect 252804 704838 253404 705800
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 701792 253404 704282
rect 252804 701728 252832 701792
rect 252896 701728 252912 701792
rect 252976 701728 252992 701792
rect 253056 701728 253072 701792
rect 253136 701728 253152 701792
rect 253216 701728 253232 701792
rect 253296 701728 253312 701792
rect 253376 701728 253404 701792
rect 252804 700704 253404 701728
rect 252804 700640 252832 700704
rect 252896 700640 252912 700704
rect 252976 700640 252992 700704
rect 253056 700640 253072 700704
rect 253136 700640 253152 700704
rect 253216 700640 253232 700704
rect 253296 700640 253312 700704
rect 253376 700640 253404 700704
rect 252804 699616 253404 700640
rect 252804 699552 252832 699616
rect 252896 699552 252912 699616
rect 252976 699552 252992 699616
rect 253056 699552 253072 699616
rect 253136 699552 253152 699616
rect 253216 699552 253232 699616
rect 253296 699552 253312 699616
rect 253376 699552 253404 699616
rect 252804 698528 253404 699552
rect 252804 698464 252832 698528
rect 252896 698464 252912 698528
rect 252976 698464 252992 698528
rect 253056 698464 253072 698528
rect 253136 698464 253152 698528
rect 253216 698464 253232 698528
rect 253296 698464 253312 698528
rect 253376 698464 253404 698528
rect 252804 697952 253404 698464
rect 256404 698000 257004 706162
rect 260004 698000 260604 708042
rect 263604 698000 264204 709922
rect 281604 711418 282204 711440
rect 281604 711182 281786 711418
rect 282022 711182 282204 711418
rect 281604 711098 282204 711182
rect 281604 710862 281786 711098
rect 282022 710862 282204 711098
rect 278004 709538 278604 709560
rect 278004 709302 278186 709538
rect 278422 709302 278604 709538
rect 278004 709218 278604 709302
rect 278004 708982 278186 709218
rect 278422 708982 278604 709218
rect 274404 707658 275004 707680
rect 274404 707422 274586 707658
rect 274822 707422 275004 707658
rect 274404 707338 275004 707422
rect 274404 707102 274586 707338
rect 274822 707102 275004 707338
rect 270804 705778 271404 705800
rect 270804 705542 270986 705778
rect 271222 705542 271404 705778
rect 270804 705458 271404 705542
rect 270804 705222 270986 705458
rect 271222 705222 271404 705458
rect 270804 701248 271404 705222
rect 270804 701184 270832 701248
rect 270896 701184 270912 701248
rect 270976 701184 270992 701248
rect 271056 701184 271072 701248
rect 271136 701184 271152 701248
rect 271216 701184 271232 701248
rect 271296 701184 271312 701248
rect 271376 701184 271404 701248
rect 270804 700160 271404 701184
rect 270804 700096 270832 700160
rect 270896 700096 270912 700160
rect 270976 700096 270992 700160
rect 271056 700096 271072 700160
rect 271136 700096 271152 700160
rect 271216 700096 271232 700160
rect 271296 700096 271312 700160
rect 271376 700096 271404 700160
rect 269067 699820 269133 699821
rect 269067 699756 269068 699820
rect 269132 699756 269133 699820
rect 269067 699755 269133 699756
rect 269070 699549 269130 699755
rect 269067 699548 269133 699549
rect 269067 699484 269068 699548
rect 269132 699484 269133 699548
rect 269067 699483 269133 699484
rect 270804 699072 271404 700096
rect 270804 699008 270832 699072
rect 270896 699008 270912 699072
rect 270976 699008 270992 699072
rect 271056 699008 271072 699072
rect 271136 699008 271152 699072
rect 271216 699008 271232 699072
rect 271296 699008 271312 699072
rect 271376 699008 271404 699072
rect 270804 697952 271404 699008
rect 274404 698000 275004 707102
rect 278004 698000 278604 708982
rect 281604 698000 282204 710862
rect 299604 710478 300204 711440
rect 299604 710242 299786 710478
rect 300022 710242 300204 710478
rect 299604 710158 300204 710242
rect 299604 709922 299786 710158
rect 300022 709922 300204 710158
rect 296004 708598 296604 709560
rect 296004 708362 296186 708598
rect 296422 708362 296604 708598
rect 296004 708278 296604 708362
rect 296004 708042 296186 708278
rect 296422 708042 296604 708278
rect 292404 706718 293004 707680
rect 292404 706482 292586 706718
rect 292822 706482 293004 706718
rect 292404 706398 293004 706482
rect 292404 706162 292586 706398
rect 292822 706162 293004 706398
rect 288804 704838 289404 705800
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 701792 289404 704282
rect 288804 701728 288832 701792
rect 288896 701728 288912 701792
rect 288976 701728 288992 701792
rect 289056 701728 289072 701792
rect 289136 701728 289152 701792
rect 289216 701728 289232 701792
rect 289296 701728 289312 701792
rect 289376 701728 289404 701792
rect 288804 700704 289404 701728
rect 288804 700640 288832 700704
rect 288896 700640 288912 700704
rect 288976 700640 288992 700704
rect 289056 700640 289072 700704
rect 289136 700640 289152 700704
rect 289216 700640 289232 700704
rect 289296 700640 289312 700704
rect 289376 700640 289404 700704
rect 288804 699616 289404 700640
rect 288804 699552 288832 699616
rect 288896 699552 288912 699616
rect 288976 699552 288992 699616
rect 289056 699552 289072 699616
rect 289136 699552 289152 699616
rect 289216 699552 289232 699616
rect 289296 699552 289312 699616
rect 289376 699552 289404 699616
rect 288804 698528 289404 699552
rect 288804 698464 288832 698528
rect 288896 698464 288912 698528
rect 288976 698464 288992 698528
rect 289056 698464 289072 698528
rect 289136 698464 289152 698528
rect 289216 698464 289232 698528
rect 289296 698464 289312 698528
rect 289376 698464 289404 698528
rect 288804 697952 289404 698464
rect 292404 698000 293004 706162
rect 296004 698000 296604 708042
rect 299604 698000 300204 709922
rect 317604 711418 318204 711440
rect 317604 711182 317786 711418
rect 318022 711182 318204 711418
rect 317604 711098 318204 711182
rect 317604 710862 317786 711098
rect 318022 710862 318204 711098
rect 314004 709538 314604 709560
rect 314004 709302 314186 709538
rect 314422 709302 314604 709538
rect 314004 709218 314604 709302
rect 314004 708982 314186 709218
rect 314422 708982 314604 709218
rect 310404 707658 311004 707680
rect 310404 707422 310586 707658
rect 310822 707422 311004 707658
rect 310404 707338 311004 707422
rect 310404 707102 310586 707338
rect 310822 707102 311004 707338
rect 306804 705778 307404 705800
rect 306804 705542 306986 705778
rect 307222 705542 307404 705778
rect 306804 705458 307404 705542
rect 306804 705222 306986 705458
rect 307222 705222 307404 705458
rect 306804 701248 307404 705222
rect 306804 701184 306832 701248
rect 306896 701184 306912 701248
rect 306976 701184 306992 701248
rect 307056 701184 307072 701248
rect 307136 701184 307152 701248
rect 307216 701184 307232 701248
rect 307296 701184 307312 701248
rect 307376 701184 307404 701248
rect 306804 700160 307404 701184
rect 306804 700096 306832 700160
rect 306896 700096 306912 700160
rect 306976 700096 306992 700160
rect 307056 700096 307072 700160
rect 307136 700096 307152 700160
rect 307216 700096 307232 700160
rect 307296 700096 307312 700160
rect 307376 700096 307404 700160
rect 306804 699072 307404 700096
rect 306804 699008 306832 699072
rect 306896 699008 306912 699072
rect 306976 699008 306992 699072
rect 307056 699008 307072 699072
rect 307136 699008 307152 699072
rect 307216 699008 307232 699072
rect 307296 699008 307312 699072
rect 307376 699008 307404 699072
rect 306804 697952 307404 699008
rect 310404 698000 311004 707102
rect 314004 698000 314604 708982
rect 317604 698000 318204 710862
rect 335604 710478 336204 711440
rect 335604 710242 335786 710478
rect 336022 710242 336204 710478
rect 335604 710158 336204 710242
rect 335604 709922 335786 710158
rect 336022 709922 336204 710158
rect 332004 708598 332604 709560
rect 332004 708362 332186 708598
rect 332422 708362 332604 708598
rect 332004 708278 332604 708362
rect 332004 708042 332186 708278
rect 332422 708042 332604 708278
rect 328404 706718 329004 707680
rect 328404 706482 328586 706718
rect 328822 706482 329004 706718
rect 328404 706398 329004 706482
rect 328404 706162 328586 706398
rect 328822 706162 329004 706398
rect 324804 704838 325404 705800
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 701792 325404 704282
rect 324804 701728 324832 701792
rect 324896 701728 324912 701792
rect 324976 701728 324992 701792
rect 325056 701728 325072 701792
rect 325136 701728 325152 701792
rect 325216 701728 325232 701792
rect 325296 701728 325312 701792
rect 325376 701728 325404 701792
rect 324804 700704 325404 701728
rect 324804 700640 324832 700704
rect 324896 700640 324912 700704
rect 324976 700640 324992 700704
rect 325056 700640 325072 700704
rect 325136 700640 325152 700704
rect 325216 700640 325232 700704
rect 325296 700640 325312 700704
rect 325376 700640 325404 700704
rect 324804 699616 325404 700640
rect 324804 699552 324832 699616
rect 324896 699552 324912 699616
rect 324976 699552 324992 699616
rect 325056 699552 325072 699616
rect 325136 699552 325152 699616
rect 325216 699552 325232 699616
rect 325296 699552 325312 699616
rect 325376 699552 325404 699616
rect 324804 698528 325404 699552
rect 324804 698464 324832 698528
rect 324896 698464 324912 698528
rect 324976 698464 324992 698528
rect 325056 698464 325072 698528
rect 325136 698464 325152 698528
rect 325216 698464 325232 698528
rect 325296 698464 325312 698528
rect 325376 698464 325404 698528
rect 324804 697952 325404 698464
rect 328404 698000 329004 706162
rect 332004 698000 332604 708042
rect 335604 698000 336204 709922
rect 353604 711418 354204 711440
rect 353604 711182 353786 711418
rect 354022 711182 354204 711418
rect 353604 711098 354204 711182
rect 353604 710862 353786 711098
rect 354022 710862 354204 711098
rect 350004 709538 350604 709560
rect 350004 709302 350186 709538
rect 350422 709302 350604 709538
rect 350004 709218 350604 709302
rect 350004 708982 350186 709218
rect 350422 708982 350604 709218
rect 346404 707658 347004 707680
rect 346404 707422 346586 707658
rect 346822 707422 347004 707658
rect 346404 707338 347004 707422
rect 346404 707102 346586 707338
rect 346822 707102 347004 707338
rect 342804 705778 343404 705800
rect 342804 705542 342986 705778
rect 343222 705542 343404 705778
rect 342804 705458 343404 705542
rect 342804 705222 342986 705458
rect 343222 705222 343404 705458
rect 342804 701248 343404 705222
rect 342804 701184 342832 701248
rect 342896 701184 342912 701248
rect 342976 701184 342992 701248
rect 343056 701184 343072 701248
rect 343136 701184 343152 701248
rect 343216 701184 343232 701248
rect 343296 701184 343312 701248
rect 343376 701184 343404 701248
rect 342804 700160 343404 701184
rect 342804 700096 342832 700160
rect 342896 700096 342912 700160
rect 342976 700096 342992 700160
rect 343056 700096 343072 700160
rect 343136 700096 343152 700160
rect 343216 700096 343232 700160
rect 343296 700096 343312 700160
rect 343376 700096 343404 700160
rect 342804 699072 343404 700096
rect 342804 699008 342832 699072
rect 342896 699008 342912 699072
rect 342976 699008 342992 699072
rect 343056 699008 343072 699072
rect 343136 699008 343152 699072
rect 343216 699008 343232 699072
rect 343296 699008 343312 699072
rect 343376 699008 343404 699072
rect 342804 697952 343404 699008
rect 346404 698000 347004 707102
rect 350004 698000 350604 708982
rect 353604 698000 354204 710862
rect 371604 710478 372204 711440
rect 371604 710242 371786 710478
rect 372022 710242 372204 710478
rect 371604 710158 372204 710242
rect 371604 709922 371786 710158
rect 372022 709922 372204 710158
rect 368004 708598 368604 709560
rect 368004 708362 368186 708598
rect 368422 708362 368604 708598
rect 368004 708278 368604 708362
rect 368004 708042 368186 708278
rect 368422 708042 368604 708278
rect 364404 706718 365004 707680
rect 364404 706482 364586 706718
rect 364822 706482 365004 706718
rect 364404 706398 365004 706482
rect 364404 706162 364586 706398
rect 364822 706162 365004 706398
rect 360804 704838 361404 705800
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 701792 361404 704282
rect 360804 701728 360832 701792
rect 360896 701728 360912 701792
rect 360976 701728 360992 701792
rect 361056 701728 361072 701792
rect 361136 701728 361152 701792
rect 361216 701728 361232 701792
rect 361296 701728 361312 701792
rect 361376 701728 361404 701792
rect 360804 700704 361404 701728
rect 360804 700640 360832 700704
rect 360896 700640 360912 700704
rect 360976 700640 360992 700704
rect 361056 700640 361072 700704
rect 361136 700640 361152 700704
rect 361216 700640 361232 700704
rect 361296 700640 361312 700704
rect 361376 700640 361404 700704
rect 360804 699616 361404 700640
rect 360804 699552 360832 699616
rect 360896 699552 360912 699616
rect 360976 699552 360992 699616
rect 361056 699552 361072 699616
rect 361136 699552 361152 699616
rect 361216 699552 361232 699616
rect 361296 699552 361312 699616
rect 361376 699552 361404 699616
rect 360804 698528 361404 699552
rect 360804 698464 360832 698528
rect 360896 698464 360912 698528
rect 360976 698464 360992 698528
rect 361056 698464 361072 698528
rect 361136 698464 361152 698528
rect 361216 698464 361232 698528
rect 361296 698464 361312 698528
rect 361376 698464 361404 698528
rect 360804 697952 361404 698464
rect 364404 698000 365004 706162
rect 368004 698000 368604 708042
rect 371604 698000 372204 709922
rect 389604 711418 390204 711440
rect 389604 711182 389786 711418
rect 390022 711182 390204 711418
rect 389604 711098 390204 711182
rect 389604 710862 389786 711098
rect 390022 710862 390204 711098
rect 386004 709538 386604 709560
rect 386004 709302 386186 709538
rect 386422 709302 386604 709538
rect 386004 709218 386604 709302
rect 386004 708982 386186 709218
rect 386422 708982 386604 709218
rect 382404 707658 383004 707680
rect 382404 707422 382586 707658
rect 382822 707422 383004 707658
rect 382404 707338 383004 707422
rect 382404 707102 382586 707338
rect 382822 707102 383004 707338
rect 378804 705778 379404 705800
rect 378804 705542 378986 705778
rect 379222 705542 379404 705778
rect 378804 705458 379404 705542
rect 378804 705222 378986 705458
rect 379222 705222 379404 705458
rect 378804 701248 379404 705222
rect 378804 701184 378832 701248
rect 378896 701184 378912 701248
rect 378976 701184 378992 701248
rect 379056 701184 379072 701248
rect 379136 701184 379152 701248
rect 379216 701184 379232 701248
rect 379296 701184 379312 701248
rect 379376 701184 379404 701248
rect 378804 700160 379404 701184
rect 378804 700096 378832 700160
rect 378896 700096 378912 700160
rect 378976 700096 378992 700160
rect 379056 700096 379072 700160
rect 379136 700096 379152 700160
rect 379216 700096 379232 700160
rect 379296 700096 379312 700160
rect 379376 700096 379404 700160
rect 378804 699072 379404 700096
rect 378804 699008 378832 699072
rect 378896 699008 378912 699072
rect 378976 699008 378992 699072
rect 379056 699008 379072 699072
rect 379136 699008 379152 699072
rect 379216 699008 379232 699072
rect 379296 699008 379312 699072
rect 379376 699008 379404 699072
rect 378804 697952 379404 699008
rect 382404 698000 383004 707102
rect 386004 698000 386604 708982
rect 389604 698000 390204 710862
rect 407604 710478 408204 711440
rect 407604 710242 407786 710478
rect 408022 710242 408204 710478
rect 407604 710158 408204 710242
rect 407604 709922 407786 710158
rect 408022 709922 408204 710158
rect 404004 708598 404604 709560
rect 404004 708362 404186 708598
rect 404422 708362 404604 708598
rect 404004 708278 404604 708362
rect 404004 708042 404186 708278
rect 404422 708042 404604 708278
rect 400404 706718 401004 707680
rect 400404 706482 400586 706718
rect 400822 706482 401004 706718
rect 400404 706398 401004 706482
rect 400404 706162 400586 706398
rect 400822 706162 401004 706398
rect 396804 704838 397404 705800
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 701792 397404 704282
rect 396804 701728 396832 701792
rect 396896 701728 396912 701792
rect 396976 701728 396992 701792
rect 397056 701728 397072 701792
rect 397136 701728 397152 701792
rect 397216 701728 397232 701792
rect 397296 701728 397312 701792
rect 397376 701728 397404 701792
rect 396804 700704 397404 701728
rect 396804 700640 396832 700704
rect 396896 700640 396912 700704
rect 396976 700640 396992 700704
rect 397056 700640 397072 700704
rect 397136 700640 397152 700704
rect 397216 700640 397232 700704
rect 397296 700640 397312 700704
rect 397376 700640 397404 700704
rect 396804 699616 397404 700640
rect 396804 699552 396832 699616
rect 396896 699552 396912 699616
rect 396976 699552 396992 699616
rect 397056 699552 397072 699616
rect 397136 699552 397152 699616
rect 397216 699552 397232 699616
rect 397296 699552 397312 699616
rect 397376 699552 397404 699616
rect 396804 698528 397404 699552
rect 396804 698464 396832 698528
rect 396896 698464 396912 698528
rect 396976 698464 396992 698528
rect 397056 698464 397072 698528
rect 397136 698464 397152 698528
rect 397216 698464 397232 698528
rect 397296 698464 397312 698528
rect 397376 698464 397404 698528
rect 396804 697952 397404 698464
rect 400404 698000 401004 706162
rect 404004 698000 404604 708042
rect 407604 698000 408204 709922
rect 425604 711418 426204 711440
rect 425604 711182 425786 711418
rect 426022 711182 426204 711418
rect 425604 711098 426204 711182
rect 425604 710862 425786 711098
rect 426022 710862 426204 711098
rect 422004 709538 422604 709560
rect 422004 709302 422186 709538
rect 422422 709302 422604 709538
rect 422004 709218 422604 709302
rect 422004 708982 422186 709218
rect 422422 708982 422604 709218
rect 418404 707658 419004 707680
rect 418404 707422 418586 707658
rect 418822 707422 419004 707658
rect 418404 707338 419004 707422
rect 418404 707102 418586 707338
rect 418822 707102 419004 707338
rect 414804 705778 415404 705800
rect 414804 705542 414986 705778
rect 415222 705542 415404 705778
rect 414804 705458 415404 705542
rect 414804 705222 414986 705458
rect 415222 705222 415404 705458
rect 414804 701248 415404 705222
rect 414804 701184 414832 701248
rect 414896 701184 414912 701248
rect 414976 701184 414992 701248
rect 415056 701184 415072 701248
rect 415136 701184 415152 701248
rect 415216 701184 415232 701248
rect 415296 701184 415312 701248
rect 415376 701184 415404 701248
rect 414804 700160 415404 701184
rect 414804 700096 414832 700160
rect 414896 700096 414912 700160
rect 414976 700096 414992 700160
rect 415056 700096 415072 700160
rect 415136 700096 415152 700160
rect 415216 700096 415232 700160
rect 415296 700096 415312 700160
rect 415376 700096 415404 700160
rect 414804 699072 415404 700096
rect 414804 699008 414832 699072
rect 414896 699008 414912 699072
rect 414976 699008 414992 699072
rect 415056 699008 415072 699072
rect 415136 699008 415152 699072
rect 415216 699008 415232 699072
rect 415296 699008 415312 699072
rect 415376 699008 415404 699072
rect 414804 697952 415404 699008
rect 418404 698000 419004 707102
rect 422004 698000 422604 708982
rect 425604 698000 426204 710862
rect 443604 710478 444204 711440
rect 443604 710242 443786 710478
rect 444022 710242 444204 710478
rect 443604 710158 444204 710242
rect 443604 709922 443786 710158
rect 444022 709922 444204 710158
rect 440004 708598 440604 709560
rect 440004 708362 440186 708598
rect 440422 708362 440604 708598
rect 440004 708278 440604 708362
rect 440004 708042 440186 708278
rect 440422 708042 440604 708278
rect 436404 706718 437004 707680
rect 436404 706482 436586 706718
rect 436822 706482 437004 706718
rect 436404 706398 437004 706482
rect 436404 706162 436586 706398
rect 436822 706162 437004 706398
rect 432804 704838 433404 705800
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 701792 433404 704282
rect 432804 701728 432832 701792
rect 432896 701728 432912 701792
rect 432976 701728 432992 701792
rect 433056 701728 433072 701792
rect 433136 701728 433152 701792
rect 433216 701728 433232 701792
rect 433296 701728 433312 701792
rect 433376 701728 433404 701792
rect 432804 700704 433404 701728
rect 432804 700640 432832 700704
rect 432896 700640 432912 700704
rect 432976 700640 432992 700704
rect 433056 700640 433072 700704
rect 433136 700640 433152 700704
rect 433216 700640 433232 700704
rect 433296 700640 433312 700704
rect 433376 700640 433404 700704
rect 432804 699616 433404 700640
rect 432804 699552 432832 699616
rect 432896 699552 432912 699616
rect 432976 699552 432992 699616
rect 433056 699552 433072 699616
rect 433136 699552 433152 699616
rect 433216 699552 433232 699616
rect 433296 699552 433312 699616
rect 433376 699552 433404 699616
rect 432804 698528 433404 699552
rect 432804 698464 432832 698528
rect 432896 698464 432912 698528
rect 432976 698464 432992 698528
rect 433056 698464 433072 698528
rect 433136 698464 433152 698528
rect 433216 698464 433232 698528
rect 433296 698464 433312 698528
rect 433376 698464 433404 698528
rect 432804 697952 433404 698464
rect 436404 698000 437004 706162
rect 440004 698000 440604 708042
rect 443604 698000 444204 709922
rect 461604 711418 462204 711440
rect 461604 711182 461786 711418
rect 462022 711182 462204 711418
rect 461604 711098 462204 711182
rect 461604 710862 461786 711098
rect 462022 710862 462204 711098
rect 458004 709538 458604 709560
rect 458004 709302 458186 709538
rect 458422 709302 458604 709538
rect 458004 709218 458604 709302
rect 458004 708982 458186 709218
rect 458422 708982 458604 709218
rect 454404 707658 455004 707680
rect 454404 707422 454586 707658
rect 454822 707422 455004 707658
rect 454404 707338 455004 707422
rect 454404 707102 454586 707338
rect 454822 707102 455004 707338
rect 450804 705778 451404 705800
rect 450804 705542 450986 705778
rect 451222 705542 451404 705778
rect 450804 705458 451404 705542
rect 450804 705222 450986 705458
rect 451222 705222 451404 705458
rect 450804 701248 451404 705222
rect 450804 701184 450832 701248
rect 450896 701184 450912 701248
rect 450976 701184 450992 701248
rect 451056 701184 451072 701248
rect 451136 701184 451152 701248
rect 451216 701184 451232 701248
rect 451296 701184 451312 701248
rect 451376 701184 451404 701248
rect 450804 700160 451404 701184
rect 450804 700096 450832 700160
rect 450896 700096 450912 700160
rect 450976 700096 450992 700160
rect 451056 700096 451072 700160
rect 451136 700096 451152 700160
rect 451216 700096 451232 700160
rect 451296 700096 451312 700160
rect 451376 700096 451404 700160
rect 450804 699072 451404 700096
rect 450804 699008 450832 699072
rect 450896 699008 450912 699072
rect 450976 699008 450992 699072
rect 451056 699008 451072 699072
rect 451136 699008 451152 699072
rect 451216 699008 451232 699072
rect 451296 699008 451312 699072
rect 451376 699008 451404 699072
rect 450804 697952 451404 699008
rect 454404 698000 455004 707102
rect 458004 698000 458604 708982
rect 461604 698000 462204 710862
rect 479604 710478 480204 711440
rect 479604 710242 479786 710478
rect 480022 710242 480204 710478
rect 479604 710158 480204 710242
rect 479604 709922 479786 710158
rect 480022 709922 480204 710158
rect 476004 708598 476604 709560
rect 476004 708362 476186 708598
rect 476422 708362 476604 708598
rect 476004 708278 476604 708362
rect 476004 708042 476186 708278
rect 476422 708042 476604 708278
rect 472404 706718 473004 707680
rect 472404 706482 472586 706718
rect 472822 706482 473004 706718
rect 472404 706398 473004 706482
rect 472404 706162 472586 706398
rect 472822 706162 473004 706398
rect 468804 704838 469404 705800
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 701792 469404 704282
rect 468804 701728 468832 701792
rect 468896 701728 468912 701792
rect 468976 701728 468992 701792
rect 469056 701728 469072 701792
rect 469136 701728 469152 701792
rect 469216 701728 469232 701792
rect 469296 701728 469312 701792
rect 469376 701728 469404 701792
rect 468804 700704 469404 701728
rect 468804 700640 468832 700704
rect 468896 700640 468912 700704
rect 468976 700640 468992 700704
rect 469056 700640 469072 700704
rect 469136 700640 469152 700704
rect 469216 700640 469232 700704
rect 469296 700640 469312 700704
rect 469376 700640 469404 700704
rect 468804 699616 469404 700640
rect 468804 699552 468832 699616
rect 468896 699552 468912 699616
rect 468976 699552 468992 699616
rect 469056 699552 469072 699616
rect 469136 699552 469152 699616
rect 469216 699552 469232 699616
rect 469296 699552 469312 699616
rect 469376 699552 469404 699616
rect 468804 698528 469404 699552
rect 468804 698464 468832 698528
rect 468896 698464 468912 698528
rect 468976 698464 468992 698528
rect 469056 698464 469072 698528
rect 469136 698464 469152 698528
rect 469216 698464 469232 698528
rect 469296 698464 469312 698528
rect 469376 698464 469404 698528
rect 468804 697952 469404 698464
rect 472404 698000 473004 706162
rect 476004 698000 476604 708042
rect 479604 698000 480204 709922
rect 497604 711418 498204 711440
rect 497604 711182 497786 711418
rect 498022 711182 498204 711418
rect 497604 711098 498204 711182
rect 497604 710862 497786 711098
rect 498022 710862 498204 711098
rect 494004 709538 494604 709560
rect 494004 709302 494186 709538
rect 494422 709302 494604 709538
rect 494004 709218 494604 709302
rect 494004 708982 494186 709218
rect 494422 708982 494604 709218
rect 490404 707658 491004 707680
rect 490404 707422 490586 707658
rect 490822 707422 491004 707658
rect 490404 707338 491004 707422
rect 490404 707102 490586 707338
rect 490822 707102 491004 707338
rect 486804 705778 487404 705800
rect 486804 705542 486986 705778
rect 487222 705542 487404 705778
rect 486804 705458 487404 705542
rect 486804 705222 486986 705458
rect 487222 705222 487404 705458
rect 486804 701248 487404 705222
rect 486804 701184 486832 701248
rect 486896 701184 486912 701248
rect 486976 701184 486992 701248
rect 487056 701184 487072 701248
rect 487136 701184 487152 701248
rect 487216 701184 487232 701248
rect 487296 701184 487312 701248
rect 487376 701184 487404 701248
rect 486804 700160 487404 701184
rect 486804 700096 486832 700160
rect 486896 700096 486912 700160
rect 486976 700096 486992 700160
rect 487056 700096 487072 700160
rect 487136 700096 487152 700160
rect 487216 700096 487232 700160
rect 487296 700096 487312 700160
rect 487376 700096 487404 700160
rect 486804 699072 487404 700096
rect 486804 699008 486832 699072
rect 486896 699008 486912 699072
rect 486976 699008 486992 699072
rect 487056 699008 487072 699072
rect 487136 699008 487152 699072
rect 487216 699008 487232 699072
rect 487296 699008 487312 699072
rect 487376 699008 487404 699072
rect 486804 697952 487404 699008
rect 490404 698000 491004 707102
rect 494004 698000 494604 708982
rect 497604 698000 498204 710862
rect 515604 710478 516204 711440
rect 515604 710242 515786 710478
rect 516022 710242 516204 710478
rect 515604 710158 516204 710242
rect 515604 709922 515786 710158
rect 516022 709922 516204 710158
rect 512004 708598 512604 709560
rect 512004 708362 512186 708598
rect 512422 708362 512604 708598
rect 512004 708278 512604 708362
rect 512004 708042 512186 708278
rect 512422 708042 512604 708278
rect 508404 706718 509004 707680
rect 508404 706482 508586 706718
rect 508822 706482 509004 706718
rect 508404 706398 509004 706482
rect 508404 706162 508586 706398
rect 508822 706162 509004 706398
rect 504804 704838 505404 705800
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 701792 505404 704282
rect 504804 701728 504832 701792
rect 504896 701728 504912 701792
rect 504976 701728 504992 701792
rect 505056 701728 505072 701792
rect 505136 701728 505152 701792
rect 505216 701728 505232 701792
rect 505296 701728 505312 701792
rect 505376 701728 505404 701792
rect 504804 700704 505404 701728
rect 504804 700640 504832 700704
rect 504896 700640 504912 700704
rect 504976 700640 504992 700704
rect 505056 700640 505072 700704
rect 505136 700640 505152 700704
rect 505216 700640 505232 700704
rect 505296 700640 505312 700704
rect 505376 700640 505404 700704
rect 504804 699616 505404 700640
rect 504804 699552 504832 699616
rect 504896 699552 504912 699616
rect 504976 699552 504992 699616
rect 505056 699552 505072 699616
rect 505136 699552 505152 699616
rect 505216 699552 505232 699616
rect 505296 699552 505312 699616
rect 505376 699552 505404 699616
rect 503483 699276 503549 699277
rect 503483 699212 503484 699276
rect 503548 699212 503549 699276
rect 503483 699211 503549 699212
rect 241467 696012 241533 696013
rect 241467 695948 241468 696012
rect 241532 695948 241533 696012
rect 241467 695947 241533 695948
rect 260787 696012 260853 696013
rect 260787 695948 260788 696012
rect 260852 695948 260853 696012
rect 260787 695947 260853 695948
rect 318747 696012 318813 696013
rect 318747 695948 318748 696012
rect 318812 695948 318813 696012
rect 318747 695947 318813 695948
rect 473307 696012 473373 696013
rect 473307 695948 473308 696012
rect 473372 695948 473373 696012
rect 473307 695947 473373 695948
rect 144867 695876 144933 695877
rect 144867 695812 144868 695876
rect 144932 695812 144933 695876
rect 144867 695811 144933 695812
rect 144870 695605 144930 695811
rect 241470 695741 241530 695947
rect 260790 695741 260850 695947
rect 318750 695741 318810 695947
rect 347635 695876 347701 695877
rect 347635 695812 347636 695876
rect 347700 695812 347701 695876
rect 347635 695811 347701 695812
rect 367139 695876 367205 695877
rect 367139 695812 367140 695876
rect 367204 695812 367205 695876
rect 367139 695811 367205 695812
rect 434667 695876 434733 695877
rect 434667 695812 434668 695876
rect 434732 695812 434733 695876
rect 434667 695811 434733 695812
rect 442947 695876 443013 695877
rect 442947 695812 442948 695876
rect 443012 695812 443013 695876
rect 442947 695811 443013 695812
rect 463739 695876 463805 695877
rect 463739 695812 463740 695876
rect 463804 695812 463805 695876
rect 463739 695811 463805 695812
rect 241467 695740 241533 695741
rect 241467 695676 241468 695740
rect 241532 695676 241533 695740
rect 241467 695675 241533 695676
rect 260787 695740 260853 695741
rect 260787 695676 260788 695740
rect 260852 695676 260853 695740
rect 260787 695675 260853 695676
rect 318747 695740 318813 695741
rect 318747 695676 318748 695740
rect 318812 695676 318813 695740
rect 318747 695675 318813 695676
rect 347638 695605 347698 695811
rect 367142 695741 367202 695811
rect 367139 695740 367205 695741
rect 367139 695676 367140 695740
rect 367204 695676 367205 695740
rect 367139 695675 367205 695676
rect 412587 695740 412653 695741
rect 412587 695676 412588 695740
rect 412652 695676 412653 695740
rect 412587 695675 412653 695676
rect 144867 695604 144933 695605
rect 144867 695540 144868 695604
rect 144932 695540 144933 695604
rect 144867 695539 144933 695540
rect 176515 695604 176581 695605
rect 176515 695540 176516 695604
rect 176580 695540 176581 695604
rect 176515 695539 176581 695540
rect 347635 695604 347701 695605
rect 347635 695540 347636 695604
rect 347700 695540 347701 695604
rect 347635 695539 347701 695540
rect 17171 695332 17237 695333
rect 17171 695268 17172 695332
rect 17236 695268 17237 695332
rect 17171 695267 17237 695268
rect 157011 695332 157077 695333
rect 157011 695268 157012 695332
rect 157076 695268 157077 695332
rect 157011 695267 157077 695268
rect 17174 694245 17234 695267
rect 124259 694788 124325 694789
rect 124259 694724 124260 694788
rect 124324 694724 124325 694788
rect 124259 694723 124325 694724
rect 133643 694788 133709 694789
rect 133643 694724 133644 694788
rect 133708 694724 133709 694788
rect 133643 694723 133709 694724
rect 153331 694788 153397 694789
rect 153331 694724 153332 694788
rect 153396 694724 153397 694788
rect 153331 694723 153397 694724
rect 111011 694516 111077 694517
rect 111011 694452 111012 694516
rect 111076 694452 111077 694516
rect 111011 694451 111077 694452
rect 115611 694516 115677 694517
rect 115611 694452 115612 694516
rect 115676 694452 115677 694516
rect 115611 694451 115677 694452
rect 17171 694244 17237 694245
rect 17171 694180 17172 694244
rect 17236 694180 17237 694244
rect 17171 694179 17237 694180
rect 9627 694108 9693 694109
rect 9627 694044 9628 694108
rect 9692 694044 9693 694108
rect 9627 694043 9693 694044
rect 31523 694108 31589 694109
rect 31523 694044 31524 694108
rect 31588 694044 31589 694108
rect 31523 694043 31589 694044
rect 89851 694108 89917 694109
rect 89851 694044 89852 694108
rect 89916 694044 89917 694108
rect 89851 694043 89917 694044
rect 96659 694108 96725 694109
rect 96659 694044 96660 694108
rect 96724 694044 96725 694108
rect 96659 694043 96725 694044
rect 9630 693970 9690 694043
rect 9811 693972 9877 693973
rect 9811 693970 9812 693972
rect 9630 693910 9812 693970
rect 9811 693908 9812 693910
rect 9876 693908 9877 693972
rect 31526 693970 31586 694043
rect 31891 693972 31957 693973
rect 31891 693970 31892 693972
rect 31526 693910 31892 693970
rect 9811 693907 9877 693908
rect 31891 693908 31892 693910
rect 31956 693908 31957 693972
rect 31891 693907 31957 693908
rect 37227 693972 37293 693973
rect 37227 693908 37228 693972
rect 37292 693908 37293 693972
rect 37227 693907 37293 693908
rect 46795 693972 46861 693973
rect 46795 693908 46796 693972
rect 46860 693908 46861 693972
rect 56547 693972 56613 693973
rect 46795 693907 46861 693908
rect 55630 693910 56426 693970
rect 37230 692698 37290 693907
rect 46798 692698 46858 693907
rect 55630 693837 55690 693910
rect 56366 693837 56426 693910
rect 56547 693908 56548 693972
rect 56612 693908 56613 693972
rect 56547 693907 56613 693908
rect 66115 693972 66181 693973
rect 66115 693908 66116 693972
rect 66180 693908 66181 693972
rect 75867 693972 75933 693973
rect 66115 693907 66181 693908
rect 74950 693910 75746 693970
rect 55627 693836 55693 693837
rect 55627 693772 55628 693836
rect 55692 693772 55693 693836
rect 55627 693771 55693 693772
rect 56363 693836 56429 693837
rect 56363 693772 56364 693836
rect 56428 693772 56429 693836
rect 56363 693771 56429 693772
rect 56550 692698 56610 693907
rect 66118 692698 66178 693907
rect 74950 693837 75010 693910
rect 75686 693837 75746 693910
rect 75867 693908 75868 693972
rect 75932 693908 75933 693972
rect 75867 693907 75933 693908
rect 85435 693972 85501 693973
rect 85435 693908 85436 693972
rect 85500 693908 85501 693972
rect 85435 693907 85501 693908
rect 89483 693972 89549 693973
rect 89483 693908 89484 693972
rect 89548 693970 89549 693972
rect 89854 693970 89914 694043
rect 89548 693910 89914 693970
rect 96662 693970 96722 694043
rect 111014 693973 111074 694451
rect 115614 693973 115674 694451
rect 124262 694245 124322 694723
rect 133646 694381 133706 694723
rect 133643 694380 133709 694381
rect 133643 694316 133644 694380
rect 133708 694316 133709 694380
rect 133643 694315 133709 694316
rect 153147 694380 153213 694381
rect 153147 694316 153148 694380
rect 153212 694378 153213 694380
rect 153334 694378 153394 694723
rect 153212 694318 153394 694378
rect 153212 694316 153213 694318
rect 153147 694315 153213 694316
rect 124259 694244 124325 694245
rect 124259 694180 124260 694244
rect 124324 694180 124325 694244
rect 124259 694179 124325 694180
rect 140819 694108 140885 694109
rect 140819 694044 140820 694108
rect 140884 694044 140885 694108
rect 140819 694043 140885 694044
rect 143579 694108 143645 694109
rect 143579 694044 143580 694108
rect 143644 694044 143645 694108
rect 143579 694043 143645 694044
rect 152963 694108 153029 694109
rect 152963 694044 152964 694108
rect 153028 694044 153029 694108
rect 152963 694043 153029 694044
rect 96843 693972 96909 693973
rect 96843 693970 96844 693972
rect 96662 693910 96844 693970
rect 89548 693908 89549 693910
rect 89483 693907 89549 693908
rect 96843 693908 96844 693910
rect 96908 693908 96909 693972
rect 96843 693907 96909 693908
rect 111011 693972 111077 693973
rect 111011 693908 111012 693972
rect 111076 693908 111077 693972
rect 111011 693907 111077 693908
rect 115611 693972 115677 693973
rect 115611 693908 115612 693972
rect 115676 693908 115677 693972
rect 124259 693972 124325 693973
rect 115611 693907 115677 693908
rect 123710 693910 124138 693970
rect 74947 693836 75013 693837
rect 74947 693772 74948 693836
rect 75012 693772 75013 693836
rect 74947 693771 75013 693772
rect 75683 693836 75749 693837
rect 75683 693772 75684 693836
rect 75748 693772 75749 693836
rect 75683 693771 75749 693772
rect 75870 692698 75930 693907
rect 85438 693834 85498 693907
rect 84334 693774 85498 693834
rect 108803 693836 108869 693837
rect 84334 692698 84394 693774
rect 108803 693772 108804 693836
rect 108868 693772 108869 693836
rect 108803 693771 108869 693772
rect 114139 693836 114205 693837
rect 114139 693772 114140 693836
rect 114204 693772 114205 693836
rect 114139 693771 114205 693772
rect 108806 692698 108866 693771
rect 114142 692698 114202 693771
rect 123710 693701 123770 693910
rect 124078 693701 124138 693910
rect 124259 693908 124260 693972
rect 124324 693908 124325 693972
rect 133643 693972 133709 693973
rect 133643 693970 133644 693972
rect 124259 693907 124325 693908
rect 133462 693910 133644 693970
rect 123707 693700 123773 693701
rect 123707 693636 123708 693700
rect 123772 693636 123773 693700
rect 123707 693635 123773 693636
rect 124075 693700 124141 693701
rect 124075 693636 124076 693700
rect 124140 693636 124141 693700
rect 124075 693635 124141 693636
rect 124262 692698 124322 693907
rect 133462 692698 133522 693910
rect 133643 693908 133644 693910
rect 133708 693908 133709 693972
rect 133643 693907 133709 693908
rect 140635 693972 140701 693973
rect 140635 693908 140636 693972
rect 140700 693970 140701 693972
rect 140822 693970 140882 694043
rect 140700 693910 140882 693970
rect 143582 693970 143642 694043
rect 152966 693970 153026 694043
rect 157014 693973 157074 695267
rect 176518 694925 176578 695539
rect 412590 695333 412650 695675
rect 434670 695605 434730 695811
rect 426387 695604 426453 695605
rect 426387 695540 426388 695604
rect 426452 695540 426453 695604
rect 426387 695539 426453 695540
rect 434667 695604 434733 695605
rect 434667 695540 434668 695604
rect 434732 695540 434733 695604
rect 434667 695539 434733 695540
rect 412587 695332 412653 695333
rect 412587 695268 412588 695332
rect 412652 695268 412653 695332
rect 412587 695267 412653 695268
rect 176515 694924 176581 694925
rect 176515 694860 176516 694924
rect 176580 694860 176581 694924
rect 176515 694859 176581 694860
rect 178907 694924 178973 694925
rect 178907 694860 178908 694924
rect 178972 694860 178973 694924
rect 178907 694859 178973 694860
rect 311571 694924 311637 694925
rect 311571 694860 311572 694924
rect 311636 694860 311637 694924
rect 311571 694859 311637 694860
rect 321507 694924 321573 694925
rect 321507 694860 321508 694924
rect 321572 694860 321573 694924
rect 321507 694859 321573 694860
rect 323715 694924 323781 694925
rect 323715 694860 323716 694924
rect 323780 694860 323781 694924
rect 323715 694859 323781 694860
rect 160875 694380 160941 694381
rect 160875 694316 160876 694380
rect 160940 694316 160941 694380
rect 160875 694315 160941 694316
rect 164187 694380 164253 694381
rect 164187 694316 164188 694380
rect 164252 694316 164253 694380
rect 164187 694315 164253 694316
rect 160878 694109 160938 694315
rect 164190 694109 164250 694315
rect 178910 694245 178970 694859
rect 273299 694788 273365 694789
rect 273299 694724 273300 694788
rect 273364 694724 273365 694788
rect 273299 694723 273365 694724
rect 279923 694788 279989 694789
rect 279923 694724 279924 694788
rect 279988 694724 279989 694788
rect 279923 694723 279989 694724
rect 299795 694788 299861 694789
rect 299795 694724 299796 694788
rect 299860 694724 299861 694788
rect 299795 694723 299861 694724
rect 311203 694788 311269 694789
rect 311203 694724 311204 694788
rect 311268 694724 311269 694788
rect 311203 694723 311269 694724
rect 186267 694652 186333 694653
rect 186267 694588 186268 694652
rect 186332 694588 186333 694652
rect 186267 694587 186333 694588
rect 256003 694652 256069 694653
rect 256003 694588 256004 694652
rect 256068 694588 256069 694652
rect 256003 694587 256069 694588
rect 185899 694380 185965 694381
rect 185899 694316 185900 694380
rect 185964 694316 185965 694380
rect 185899 694315 185965 694316
rect 178907 694244 178973 694245
rect 178907 694180 178908 694244
rect 178972 694180 178973 694244
rect 178907 694179 178973 694180
rect 185902 694109 185962 694315
rect 186270 694109 186330 694587
rect 196019 694516 196085 694517
rect 196019 694514 196020 694516
rect 195838 694454 196020 694514
rect 195838 694381 195898 694454
rect 196019 694452 196020 694454
rect 196084 694452 196085 694516
rect 215339 694516 215405 694517
rect 215339 694514 215340 694516
rect 196019 694451 196085 694452
rect 215158 694454 215340 694514
rect 215158 694381 215218 694454
rect 215339 694452 215340 694454
rect 215404 694452 215405 694516
rect 215339 694451 215405 694452
rect 195835 694380 195901 694381
rect 195835 694316 195836 694380
rect 195900 694316 195901 694380
rect 195835 694315 195901 694316
rect 215155 694380 215221 694381
rect 215155 694316 215156 694380
rect 215220 694316 215221 694380
rect 215155 694315 215221 694316
rect 253795 694380 253861 694381
rect 253795 694316 253796 694380
rect 253860 694316 253861 694380
rect 253795 694315 253861 694316
rect 254347 694380 254413 694381
rect 254347 694316 254348 694380
rect 254412 694316 254413 694380
rect 254347 694315 254413 694316
rect 160875 694108 160941 694109
rect 160875 694044 160876 694108
rect 160940 694044 160941 694108
rect 160875 694043 160941 694044
rect 164187 694108 164253 694109
rect 164187 694044 164188 694108
rect 164252 694044 164253 694108
rect 164187 694043 164253 694044
rect 185899 694108 185965 694109
rect 185899 694044 185900 694108
rect 185964 694044 185965 694108
rect 185899 694043 185965 694044
rect 186267 694108 186333 694109
rect 186267 694044 186268 694108
rect 186332 694044 186333 694108
rect 186267 694043 186333 694044
rect 195835 694108 195901 694109
rect 195835 694044 195836 694108
rect 195900 694106 195901 694108
rect 196019 694108 196085 694109
rect 196019 694106 196020 694108
rect 195900 694046 196020 694106
rect 195900 694044 195901 694046
rect 195835 694043 195901 694044
rect 196019 694044 196020 694046
rect 196084 694044 196085 694108
rect 196019 694043 196085 694044
rect 205403 694108 205469 694109
rect 205403 694044 205404 694108
rect 205468 694106 205469 694108
rect 205955 694108 206021 694109
rect 205955 694106 205956 694108
rect 205468 694046 205956 694106
rect 205468 694044 205469 694046
rect 205403 694043 205469 694044
rect 205955 694044 205956 694046
rect 206020 694044 206021 694108
rect 205955 694043 206021 694044
rect 215155 694108 215221 694109
rect 215155 694044 215156 694108
rect 215220 694106 215221 694108
rect 215339 694108 215405 694109
rect 215339 694106 215340 694108
rect 215220 694046 215340 694106
rect 215220 694044 215221 694046
rect 215155 694043 215221 694044
rect 215339 694044 215340 694046
rect 215404 694044 215405 694108
rect 215339 694043 215405 694044
rect 224723 694108 224789 694109
rect 224723 694044 224724 694108
rect 224788 694106 224789 694108
rect 225275 694108 225341 694109
rect 225275 694106 225276 694108
rect 224788 694046 225276 694106
rect 224788 694044 224789 694046
rect 224723 694043 224789 694044
rect 225275 694044 225276 694046
rect 225340 694044 225341 694108
rect 225275 694043 225341 694044
rect 244043 694108 244109 694109
rect 244043 694044 244044 694108
rect 244108 694106 244109 694108
rect 244595 694108 244661 694109
rect 244595 694106 244596 694108
rect 244108 694046 244596 694106
rect 244108 694044 244109 694046
rect 244043 694043 244109 694044
rect 244595 694044 244596 694046
rect 244660 694044 244661 694108
rect 253798 694106 253858 694315
rect 254350 694106 254410 694315
rect 256006 694245 256066 694587
rect 263547 694516 263613 694517
rect 263547 694452 263548 694516
rect 263612 694452 263613 694516
rect 263547 694451 263613 694452
rect 256003 694244 256069 694245
rect 256003 694180 256004 694244
rect 256068 694180 256069 694244
rect 256003 694179 256069 694180
rect 263550 694109 263610 694451
rect 273302 694245 273362 694723
rect 275323 694652 275389 694653
rect 275323 694588 275324 694652
rect 275388 694588 275389 694652
rect 275323 694587 275389 694588
rect 273667 694516 273733 694517
rect 273667 694452 273668 694516
rect 273732 694452 273733 694516
rect 273667 694451 273733 694452
rect 273299 694244 273365 694245
rect 273299 694180 273300 694244
rect 273364 694180 273365 694244
rect 273299 694179 273365 694180
rect 273670 694109 273730 694451
rect 275326 694245 275386 694587
rect 279926 694514 279986 694723
rect 284891 694652 284957 694653
rect 282686 694590 283298 694650
rect 279926 694454 280124 694514
rect 280064 694381 280124 694454
rect 282686 694381 282746 694590
rect 283051 694516 283117 694517
rect 283051 694452 283052 694516
rect 283116 694452 283117 694516
rect 283051 694451 283117 694452
rect 280061 694380 280127 694381
rect 280061 694316 280062 694380
rect 280126 694316 280127 694380
rect 280061 694315 280127 694316
rect 282683 694380 282749 694381
rect 282683 694316 282684 694380
rect 282748 694316 282749 694380
rect 282683 694315 282749 694316
rect 275323 694244 275389 694245
rect 275323 694180 275324 694244
rect 275388 694180 275389 694244
rect 275323 694179 275389 694180
rect 253798 694046 254410 694106
rect 263547 694108 263613 694109
rect 244595 694043 244661 694044
rect 263547 694044 263548 694108
rect 263612 694044 263613 694108
rect 263547 694043 263613 694044
rect 273667 694108 273733 694109
rect 273667 694044 273668 694108
rect 273732 694044 273733 694108
rect 273667 694043 273733 694044
rect 282867 694108 282933 694109
rect 282867 694044 282868 694108
rect 282932 694106 282933 694108
rect 283054 694106 283114 694451
rect 283238 694381 283298 694590
rect 284891 694588 284892 694652
rect 284956 694588 284957 694652
rect 284891 694587 284957 694588
rect 283235 694380 283301 694381
rect 283235 694316 283236 694380
rect 283300 694316 283301 694380
rect 283235 694315 283301 694316
rect 284894 694109 284954 694587
rect 282932 694046 283114 694106
rect 284891 694108 284957 694109
rect 282932 694044 282933 694046
rect 282867 694043 282933 694044
rect 284891 694044 284892 694108
rect 284956 694044 284957 694108
rect 284891 694043 284957 694044
rect 299243 694108 299309 694109
rect 299243 694044 299244 694108
rect 299308 694044 299309 694108
rect 299243 694043 299309 694044
rect 143582 693910 143826 693970
rect 140700 693908 140701 693910
rect 140635 693907 140701 693908
rect 143766 692698 143826 693910
rect 152782 693910 153026 693970
rect 157011 693972 157077 693973
rect 152782 692698 152842 693910
rect 157011 693908 157012 693972
rect 157076 693908 157077 693972
rect 157011 693907 157077 693908
rect 173939 693972 174005 693973
rect 173939 693908 173940 693972
rect 174004 693970 174005 693972
rect 174123 693972 174189 693973
rect 174123 693970 174124 693972
rect 174004 693910 174124 693970
rect 174004 693908 174005 693910
rect 173939 693907 174005 693908
rect 174123 693908 174124 693910
rect 174188 693908 174189 693972
rect 299246 693970 299306 694043
rect 299798 693970 299858 694723
rect 311206 694109 311266 694723
rect 311574 694381 311634 694859
rect 318747 694788 318813 694789
rect 318747 694724 318748 694788
rect 318812 694724 318813 694788
rect 318747 694723 318813 694724
rect 311755 694652 311821 694653
rect 311755 694588 311756 694652
rect 311820 694588 311821 694652
rect 318750 694650 318810 694723
rect 318931 694652 318997 694653
rect 318931 694650 318932 694652
rect 318750 694590 318932 694650
rect 311755 694587 311821 694588
rect 318931 694588 318932 694590
rect 318996 694588 318997 694652
rect 318931 694587 318997 694588
rect 311758 694381 311818 694587
rect 311571 694380 311637 694381
rect 311571 694316 311572 694380
rect 311636 694316 311637 694380
rect 311571 694315 311637 694316
rect 311755 694380 311821 694381
rect 311755 694316 311756 694380
rect 311820 694316 311821 694380
rect 311755 694315 311821 694316
rect 321510 694109 321570 694859
rect 323718 694517 323778 694859
rect 331075 694788 331141 694789
rect 331075 694724 331076 694788
rect 331140 694724 331141 694788
rect 331075 694723 331141 694724
rect 424915 694788 424981 694789
rect 424915 694724 424916 694788
rect 424980 694724 424981 694788
rect 424915 694723 424981 694724
rect 425099 694788 425165 694789
rect 425099 694724 425100 694788
rect 425164 694724 425165 694788
rect 425099 694723 425165 694724
rect 331078 694650 331138 694723
rect 331259 694652 331325 694653
rect 331259 694650 331260 694652
rect 331078 694590 331260 694650
rect 331259 694588 331260 694590
rect 331324 694588 331325 694652
rect 331259 694587 331325 694588
rect 340827 694652 340893 694653
rect 340827 694588 340828 694652
rect 340892 694588 340893 694652
rect 340827 694587 340893 694588
rect 371923 694652 371989 694653
rect 371923 694588 371924 694652
rect 371988 694588 371989 694652
rect 371923 694587 371989 694588
rect 379099 694652 379165 694653
rect 379099 694588 379100 694652
rect 379164 694588 379165 694652
rect 379099 694587 379165 694588
rect 391243 694652 391309 694653
rect 391243 694588 391244 694652
rect 391308 694588 391309 694652
rect 391243 694587 391309 694588
rect 398419 694652 398485 694653
rect 398419 694588 398420 694652
rect 398484 694588 398485 694652
rect 398419 694587 398485 694588
rect 323531 694516 323597 694517
rect 323531 694452 323532 694516
rect 323596 694452 323597 694516
rect 323531 694451 323597 694452
rect 323715 694516 323781 694517
rect 323715 694452 323716 694516
rect 323780 694452 323781 694516
rect 323715 694451 323781 694452
rect 330707 694516 330773 694517
rect 330707 694452 330708 694516
rect 330772 694452 330773 694516
rect 330707 694451 330773 694452
rect 323534 694109 323594 694451
rect 330710 694109 330770 694451
rect 340830 694109 340890 694587
rect 359963 694516 360029 694517
rect 359963 694452 359964 694516
rect 360028 694452 360029 694516
rect 369899 694516 369965 694517
rect 369899 694514 369900 694516
rect 359963 694451 360029 694452
rect 369718 694454 369900 694514
rect 359966 694378 360026 694451
rect 369718 694381 369778 694454
rect 369899 694452 369900 694454
rect 369964 694452 369965 694516
rect 369899 694451 369965 694452
rect 360331 694380 360397 694381
rect 360331 694378 360332 694380
rect 359966 694318 360332 694378
rect 360331 694316 360332 694318
rect 360396 694316 360397 694380
rect 360331 694315 360397 694316
rect 369715 694380 369781 694381
rect 369715 694316 369716 694380
rect 369780 694316 369781 694380
rect 369715 694315 369781 694316
rect 371926 694245 371986 694587
rect 379102 694245 379162 694587
rect 390139 694516 390205 694517
rect 390139 694514 390140 694516
rect 389222 694454 390140 694514
rect 389222 694381 389282 694454
rect 390139 694452 390140 694454
rect 390204 694452 390205 694516
rect 390139 694451 390205 694452
rect 389219 694380 389285 694381
rect 389219 694316 389220 694380
rect 389284 694316 389285 694380
rect 389219 694315 389285 694316
rect 391246 694245 391306 694587
rect 398422 694245 398482 694587
rect 420131 694516 420197 694517
rect 420131 694452 420132 694516
rect 420196 694452 420197 694516
rect 420131 694451 420197 694452
rect 371923 694244 371989 694245
rect 371923 694180 371924 694244
rect 371988 694180 371989 694244
rect 371923 694179 371989 694180
rect 379099 694244 379165 694245
rect 379099 694180 379100 694244
rect 379164 694180 379165 694244
rect 379099 694179 379165 694180
rect 391243 694244 391309 694245
rect 391243 694180 391244 694244
rect 391308 694180 391309 694244
rect 391243 694179 391309 694180
rect 398419 694244 398485 694245
rect 398419 694180 398420 694244
rect 398484 694180 398485 694244
rect 398419 694179 398485 694180
rect 420134 694109 420194 694451
rect 424918 694245 424978 694723
rect 420315 694244 420381 694245
rect 420315 694180 420316 694244
rect 420380 694180 420381 694244
rect 420315 694179 420381 694180
rect 424731 694244 424797 694245
rect 424731 694180 424732 694244
rect 424796 694180 424797 694244
rect 424731 694179 424797 694180
rect 424915 694244 424981 694245
rect 424915 694180 424916 694244
rect 424980 694180 424981 694244
rect 424915 694179 424981 694180
rect 311203 694108 311269 694109
rect 311203 694044 311204 694108
rect 311268 694044 311269 694108
rect 311203 694043 311269 694044
rect 321507 694108 321573 694109
rect 321507 694044 321508 694108
rect 321572 694044 321573 694108
rect 321507 694043 321573 694044
rect 323531 694108 323597 694109
rect 323531 694044 323532 694108
rect 323596 694044 323597 694108
rect 323531 694043 323597 694044
rect 330707 694108 330773 694109
rect 330707 694044 330708 694108
rect 330772 694044 330773 694108
rect 330707 694043 330773 694044
rect 340827 694108 340893 694109
rect 340827 694044 340828 694108
rect 340892 694044 340893 694108
rect 340827 694043 340893 694044
rect 359963 694108 360029 694109
rect 359963 694044 359964 694108
rect 360028 694106 360029 694108
rect 360331 694108 360397 694109
rect 360331 694106 360332 694108
rect 360028 694046 360332 694106
rect 360028 694044 360029 694046
rect 359963 694043 360029 694044
rect 360331 694044 360332 694046
rect 360396 694044 360397 694108
rect 360331 694043 360397 694044
rect 369715 694108 369781 694109
rect 369715 694044 369716 694108
rect 369780 694106 369781 694108
rect 369899 694108 369965 694109
rect 369899 694106 369900 694108
rect 369780 694046 369900 694106
rect 369780 694044 369781 694046
rect 369715 694043 369781 694044
rect 369899 694044 369900 694046
rect 369964 694044 369965 694108
rect 369899 694043 369965 694044
rect 420131 694108 420197 694109
rect 420131 694044 420132 694108
rect 420196 694044 420197 694108
rect 420131 694043 420197 694044
rect 420318 693973 420378 694179
rect 424734 694106 424794 694179
rect 425102 694109 425162 694723
rect 426390 694517 426450 695539
rect 442950 695469 443010 695811
rect 463742 695741 463802 695811
rect 463739 695740 463805 695741
rect 463739 695676 463740 695740
rect 463804 695676 463805 695740
rect 463739 695675 463805 695676
rect 473310 695605 473370 695947
rect 473307 695604 473373 695605
rect 473307 695540 473308 695604
rect 473372 695540 473373 695604
rect 473307 695539 473373 695540
rect 442947 695468 443013 695469
rect 442947 695404 442948 695468
rect 443012 695404 443013 695468
rect 442947 695403 443013 695404
rect 489683 694924 489749 694925
rect 489683 694922 489684 694924
rect 489502 694862 489684 694922
rect 434299 694788 434365 694789
rect 434299 694724 434300 694788
rect 434364 694724 434365 694788
rect 434299 694723 434365 694724
rect 461163 694788 461229 694789
rect 461163 694724 461164 694788
rect 461228 694724 461229 694788
rect 461163 694723 461229 694724
rect 470363 694788 470429 694789
rect 470363 694724 470364 694788
rect 470428 694724 470429 694788
rect 470363 694723 470429 694724
rect 426387 694516 426453 694517
rect 426387 694452 426388 694516
rect 426452 694452 426453 694516
rect 434302 694514 434362 694723
rect 434302 694454 434546 694514
rect 426387 694451 426453 694452
rect 434486 694109 434546 694454
rect 460979 694244 461045 694245
rect 460979 694180 460980 694244
rect 461044 694180 461045 694244
rect 460979 694179 461045 694180
rect 425099 694108 425165 694109
rect 424734 694046 424978 694106
rect 424918 693973 424978 694046
rect 425099 694044 425100 694108
rect 425164 694044 425165 694108
rect 425099 694043 425165 694044
rect 434483 694108 434549 694109
rect 434483 694044 434484 694108
rect 434548 694044 434549 694108
rect 434483 694043 434549 694044
rect 434667 694108 434733 694109
rect 434667 694044 434668 694108
rect 434732 694106 434733 694108
rect 435035 694108 435101 694109
rect 435035 694106 435036 694108
rect 434732 694046 435036 694106
rect 434732 694044 434733 694046
rect 434667 694043 434733 694044
rect 435035 694044 435036 694046
rect 435100 694044 435101 694108
rect 435035 694043 435101 694044
rect 299246 693910 299858 693970
rect 420315 693972 420381 693973
rect 174123 693907 174189 693908
rect 420315 693908 420316 693972
rect 420380 693908 420381 693972
rect 424915 693972 424981 693973
rect 420315 693907 420381 693908
rect 423998 693910 424794 693970
rect 162899 693836 162965 693837
rect 162899 693772 162900 693836
rect 162964 693772 162965 693836
rect 162899 693771 162965 693772
rect 163819 693836 163885 693837
rect 163819 693772 163820 693836
rect 163884 693772 163885 693836
rect 163819 693771 163885 693772
rect 162902 691930 162962 693771
rect 163083 693700 163149 693701
rect 163083 693636 163084 693700
rect 163148 693636 163149 693700
rect 163083 693635 163149 693636
rect 163635 693700 163701 693701
rect 163635 693636 163636 693700
rect 163700 693636 163701 693700
rect 163635 693635 163701 693636
rect 163086 692610 163146 693635
rect 163638 692610 163698 693635
rect 163086 692550 163698 692610
rect 163822 691930 163882 693771
rect 423998 693701 424058 693910
rect 424179 693836 424245 693837
rect 424179 693772 424180 693836
rect 424244 693772 424245 693836
rect 424179 693771 424245 693772
rect 423995 693700 424061 693701
rect 423995 693636 423996 693700
rect 424060 693636 424061 693700
rect 423995 693635 424061 693636
rect 424182 693290 424242 693771
rect 424734 693701 424794 693910
rect 424915 693908 424916 693972
rect 424980 693908 424981 693972
rect 434667 693972 434733 693973
rect 424915 693907 424981 693908
rect 434118 693910 434546 693970
rect 434118 693837 434178 693910
rect 434486 693837 434546 693910
rect 434667 693908 434668 693972
rect 434732 693970 434733 693972
rect 435035 693972 435101 693973
rect 435035 693970 435036 693972
rect 434732 693910 435036 693970
rect 434732 693908 434733 693910
rect 434667 693907 434733 693908
rect 435035 693908 435036 693910
rect 435100 693908 435101 693972
rect 460982 693970 461042 694179
rect 461166 693970 461226 694723
rect 470366 694381 470426 694723
rect 470547 694652 470613 694653
rect 470547 694588 470548 694652
rect 470612 694588 470613 694652
rect 470547 694587 470613 694588
rect 470550 694381 470610 694587
rect 489502 694381 489562 694862
rect 489683 694860 489684 694862
rect 489748 694860 489749 694924
rect 489683 694859 489749 694860
rect 500907 694516 500973 694517
rect 500907 694452 500908 694516
rect 500972 694452 500973 694516
rect 500907 694451 500973 694452
rect 470363 694380 470429 694381
rect 470363 694316 470364 694380
rect 470428 694316 470429 694380
rect 470363 694315 470429 694316
rect 470547 694380 470613 694381
rect 470547 694316 470548 694380
rect 470612 694316 470613 694380
rect 470547 694315 470613 694316
rect 489499 694380 489565 694381
rect 489499 694316 489500 694380
rect 489564 694316 489565 694380
rect 489499 694315 489565 694316
rect 500910 694245 500970 694451
rect 500907 694244 500973 694245
rect 500907 694180 500908 694244
rect 500972 694180 500973 694244
rect 500907 694179 500973 694180
rect 460982 693910 461226 693970
rect 435035 693907 435101 693908
rect 503486 693837 503546 699211
rect 504804 698528 505404 699552
rect 504804 698464 504832 698528
rect 504896 698464 504912 698528
rect 504976 698464 504992 698528
rect 505056 698464 505072 698528
rect 505136 698464 505152 698528
rect 505216 698464 505232 698528
rect 505296 698464 505312 698528
rect 505376 698464 505404 698528
rect 504804 697952 505404 698464
rect 508404 698000 509004 706162
rect 512004 698000 512604 708042
rect 515604 698000 516204 709922
rect 533604 711418 534204 711440
rect 533604 711182 533786 711418
rect 534022 711182 534204 711418
rect 533604 711098 534204 711182
rect 533604 710862 533786 711098
rect 534022 710862 534204 711098
rect 530004 709538 530604 709560
rect 530004 709302 530186 709538
rect 530422 709302 530604 709538
rect 530004 709218 530604 709302
rect 530004 708982 530186 709218
rect 530422 708982 530604 709218
rect 526404 707658 527004 707680
rect 526404 707422 526586 707658
rect 526822 707422 527004 707658
rect 526404 707338 527004 707422
rect 526404 707102 526586 707338
rect 526822 707102 527004 707338
rect 522804 705778 523404 705800
rect 522804 705542 522986 705778
rect 523222 705542 523404 705778
rect 522804 705458 523404 705542
rect 522804 705222 522986 705458
rect 523222 705222 523404 705458
rect 522804 701248 523404 705222
rect 522804 701184 522832 701248
rect 522896 701184 522912 701248
rect 522976 701184 522992 701248
rect 523056 701184 523072 701248
rect 523136 701184 523152 701248
rect 523216 701184 523232 701248
rect 523296 701184 523312 701248
rect 523376 701184 523404 701248
rect 522804 700160 523404 701184
rect 522804 700096 522832 700160
rect 522896 700096 522912 700160
rect 522976 700096 522992 700160
rect 523056 700096 523072 700160
rect 523136 700096 523152 700160
rect 523216 700096 523232 700160
rect 523296 700096 523312 700160
rect 523376 700096 523404 700160
rect 522804 699072 523404 700096
rect 522804 699008 522832 699072
rect 522896 699008 522912 699072
rect 522976 699008 522992 699072
rect 523056 699008 523072 699072
rect 523136 699008 523152 699072
rect 523216 699008 523232 699072
rect 523296 699008 523312 699072
rect 523376 699008 523404 699072
rect 522804 697952 523404 699008
rect 526404 698000 527004 707102
rect 530004 698000 530604 708982
rect 533604 698000 534204 710862
rect 551604 710478 552204 711440
rect 551604 710242 551786 710478
rect 552022 710242 552204 710478
rect 551604 710158 552204 710242
rect 551604 709922 551786 710158
rect 552022 709922 552204 710158
rect 548004 708598 548604 709560
rect 548004 708362 548186 708598
rect 548422 708362 548604 708598
rect 548004 708278 548604 708362
rect 548004 708042 548186 708278
rect 548422 708042 548604 708278
rect 544404 706718 545004 707680
rect 544404 706482 544586 706718
rect 544822 706482 545004 706718
rect 544404 706398 545004 706482
rect 544404 706162 544586 706398
rect 544822 706162 545004 706398
rect 540804 704838 541404 705800
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 701792 541404 704282
rect 540804 701728 540832 701792
rect 540896 701728 540912 701792
rect 540976 701728 540992 701792
rect 541056 701728 541072 701792
rect 541136 701728 541152 701792
rect 541216 701728 541232 701792
rect 541296 701728 541312 701792
rect 541376 701728 541404 701792
rect 540804 700704 541404 701728
rect 540804 700640 540832 700704
rect 540896 700640 540912 700704
rect 540976 700640 540992 700704
rect 541056 700640 541072 700704
rect 541136 700640 541152 700704
rect 541216 700640 541232 700704
rect 541296 700640 541312 700704
rect 541376 700640 541404 700704
rect 540804 699616 541404 700640
rect 540804 699552 540832 699616
rect 540896 699552 540912 699616
rect 540976 699552 540992 699616
rect 541056 699552 541072 699616
rect 541136 699552 541152 699616
rect 541216 699552 541232 699616
rect 541296 699552 541312 699616
rect 541376 699552 541404 699616
rect 540804 698528 541404 699552
rect 540804 698464 540832 698528
rect 540896 698464 540912 698528
rect 540976 698464 540992 698528
rect 541056 698464 541072 698528
rect 541136 698464 541152 698528
rect 541216 698464 541232 698528
rect 541296 698464 541312 698528
rect 541376 698464 541404 698528
rect 540804 697952 541404 698464
rect 544404 698000 545004 706162
rect 548004 698000 548604 708042
rect 551604 698000 552204 709922
rect 569604 711418 570204 711440
rect 569604 711182 569786 711418
rect 570022 711182 570204 711418
rect 569604 711098 570204 711182
rect 569604 710862 569786 711098
rect 570022 710862 570204 711098
rect 566004 709538 566604 709560
rect 566004 709302 566186 709538
rect 566422 709302 566604 709538
rect 566004 709218 566604 709302
rect 566004 708982 566186 709218
rect 566422 708982 566604 709218
rect 562404 707658 563004 707680
rect 562404 707422 562586 707658
rect 562822 707422 563004 707658
rect 562404 707338 563004 707422
rect 562404 707102 562586 707338
rect 562822 707102 563004 707338
rect 558804 705778 559404 705800
rect 558804 705542 558986 705778
rect 559222 705542 559404 705778
rect 558804 705458 559404 705542
rect 558804 705222 558986 705458
rect 559222 705222 559404 705458
rect 558804 701248 559404 705222
rect 558804 701184 558832 701248
rect 558896 701184 558912 701248
rect 558976 701184 558992 701248
rect 559056 701184 559072 701248
rect 559136 701184 559152 701248
rect 559216 701184 559232 701248
rect 559296 701184 559312 701248
rect 559376 701184 559404 701248
rect 558804 700160 559404 701184
rect 558804 700096 558832 700160
rect 558896 700096 558912 700160
rect 558976 700096 558992 700160
rect 559056 700096 559072 700160
rect 559136 700096 559152 700160
rect 559216 700096 559232 700160
rect 559296 700096 559312 700160
rect 559376 700096 559404 700160
rect 558804 699072 559404 700096
rect 558804 699008 558832 699072
rect 558896 699008 558912 699072
rect 558976 699008 558992 699072
rect 559056 699008 559072 699072
rect 559136 699008 559152 699072
rect 559216 699008 559232 699072
rect 559296 699008 559312 699072
rect 559376 699008 559404 699072
rect 558804 697952 559404 699008
rect 562404 698000 563004 707102
rect 566004 698000 566604 708982
rect 569604 698000 570204 710862
rect 591900 711418 592500 711440
rect 591900 711182 592082 711418
rect 592318 711182 592500 711418
rect 591900 711098 592500 711182
rect 591900 710862 592082 711098
rect 592318 710862 592500 711098
rect 590960 710478 591560 710500
rect 590960 710242 591142 710478
rect 591378 710242 591560 710478
rect 590960 710158 591560 710242
rect 590960 709922 591142 710158
rect 591378 709922 591560 710158
rect 590020 709538 590620 709560
rect 590020 709302 590202 709538
rect 590438 709302 590620 709538
rect 590020 709218 590620 709302
rect 590020 708982 590202 709218
rect 590438 708982 590620 709218
rect 589080 708598 589680 708620
rect 589080 708362 589262 708598
rect 589498 708362 589680 708598
rect 589080 708278 589680 708362
rect 589080 708042 589262 708278
rect 589498 708042 589680 708278
rect 580404 706718 581004 707680
rect 588140 707658 588740 707680
rect 588140 707422 588322 707658
rect 588558 707422 588740 707658
rect 588140 707338 588740 707422
rect 588140 707102 588322 707338
rect 588558 707102 588740 707338
rect 580404 706482 580586 706718
rect 580822 706482 581004 706718
rect 580404 706398 581004 706482
rect 580404 706162 580586 706398
rect 580822 706162 581004 706398
rect 576804 704838 577404 705800
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 701792 577404 704282
rect 576804 701728 576832 701792
rect 576896 701728 576912 701792
rect 576976 701728 576992 701792
rect 577056 701728 577072 701792
rect 577136 701728 577152 701792
rect 577216 701728 577232 701792
rect 577296 701728 577312 701792
rect 577376 701728 577404 701792
rect 576804 700704 577404 701728
rect 576804 700640 576832 700704
rect 576896 700640 576912 700704
rect 576976 700640 576992 700704
rect 577056 700640 577072 700704
rect 577136 700640 577152 700704
rect 577216 700640 577232 700704
rect 577296 700640 577312 700704
rect 577376 700640 577404 700704
rect 576804 699616 577404 700640
rect 576804 699552 576832 699616
rect 576896 699552 576912 699616
rect 576976 699552 576992 699616
rect 577056 699552 577072 699616
rect 577136 699552 577152 699616
rect 577216 699552 577232 699616
rect 577296 699552 577312 699616
rect 577376 699552 577404 699616
rect 576804 698528 577404 699552
rect 576804 698464 576832 698528
rect 576896 698464 576912 698528
rect 576976 698464 576992 698528
rect 577056 698464 577072 698528
rect 577136 698464 577152 698528
rect 577216 698464 577232 698528
rect 577296 698464 577312 698528
rect 577376 698464 577404 698528
rect 576804 697952 577404 698464
rect 521331 695332 521397 695333
rect 521331 695268 521332 695332
rect 521396 695268 521397 695332
rect 521331 695267 521397 695268
rect 511947 694652 512013 694653
rect 511947 694588 511948 694652
rect 512012 694588 512013 694652
rect 511947 694587 512013 694588
rect 511950 694109 512010 694587
rect 511947 694108 512013 694109
rect 511947 694044 511948 694108
rect 512012 694044 512013 694108
rect 511947 694043 512013 694044
rect 424915 693836 424981 693837
rect 424915 693772 424916 693836
rect 424980 693772 424981 693836
rect 424915 693771 424981 693772
rect 434115 693836 434181 693837
rect 434115 693772 434116 693836
rect 434180 693772 434181 693836
rect 434115 693771 434181 693772
rect 434483 693836 434549 693837
rect 434483 693772 434484 693836
rect 434548 693772 434549 693836
rect 434483 693771 434549 693772
rect 434667 693836 434733 693837
rect 434667 693772 434668 693836
rect 434732 693834 434733 693836
rect 435219 693836 435285 693837
rect 435219 693834 435220 693836
rect 434732 693774 435220 693834
rect 434732 693772 434733 693774
rect 434667 693771 434733 693772
rect 435219 693772 435220 693774
rect 435284 693772 435285 693836
rect 435219 693771 435285 693772
rect 503483 693836 503549 693837
rect 503483 693772 503484 693836
rect 503548 693772 503549 693836
rect 503483 693771 503549 693772
rect 424731 693700 424797 693701
rect 424731 693636 424732 693700
rect 424796 693636 424797 693700
rect 424731 693635 424797 693636
rect 424918 693290 424978 693771
rect 521334 693701 521394 695267
rect 531267 694788 531333 694789
rect 531267 694724 531268 694788
rect 531332 694724 531333 694788
rect 531267 694723 531333 694724
rect 521515 694652 521581 694653
rect 521515 694588 521516 694652
rect 521580 694588 521581 694652
rect 521515 694587 521581 694588
rect 521518 694109 521578 694587
rect 531270 694517 531330 694723
rect 521699 694516 521765 694517
rect 521699 694452 521700 694516
rect 521764 694452 521765 694516
rect 521699 694451 521765 694452
rect 531267 694516 531333 694517
rect 531267 694452 531268 694516
rect 531332 694452 531333 694516
rect 531267 694451 531333 694452
rect 550587 694516 550653 694517
rect 550587 694452 550588 694516
rect 550652 694452 550653 694516
rect 550587 694451 550653 694452
rect 521702 694245 521762 694451
rect 550590 694245 550650 694451
rect 521699 694244 521765 694245
rect 521699 694180 521700 694244
rect 521764 694180 521765 694244
rect 521699 694179 521765 694180
rect 550587 694244 550653 694245
rect 550587 694180 550588 694244
rect 550652 694180 550653 694244
rect 550587 694179 550653 694180
rect 521515 694108 521581 694109
rect 521515 694044 521516 694108
rect 521580 694044 521581 694108
rect 521515 694043 521581 694044
rect 521699 694108 521765 694109
rect 521699 694044 521700 694108
rect 521764 694044 521765 694108
rect 521699 694043 521765 694044
rect 524459 694108 524525 694109
rect 524459 694044 524460 694108
rect 524524 694044 524525 694108
rect 524459 694043 524525 694044
rect 539547 694108 539613 694109
rect 539547 694044 539548 694108
rect 539612 694044 539613 694108
rect 539547 694043 539613 694044
rect 521702 693837 521762 694043
rect 524462 693837 524522 694043
rect 521699 693836 521765 693837
rect 521699 693772 521700 693836
rect 521764 693772 521765 693836
rect 521699 693771 521765 693772
rect 524459 693836 524525 693837
rect 524459 693772 524460 693836
rect 524524 693772 524525 693836
rect 524459 693771 524525 693772
rect 433931 693700 433997 693701
rect 433931 693636 433932 693700
rect 433996 693636 433997 693700
rect 433931 693635 433997 693636
rect 434483 693700 434549 693701
rect 434483 693636 434484 693700
rect 434548 693636 434549 693700
rect 434483 693635 434549 693636
rect 473491 693700 473557 693701
rect 473491 693636 473492 693700
rect 473556 693636 473557 693700
rect 473491 693635 473557 693636
rect 474043 693700 474109 693701
rect 474043 693636 474044 693700
rect 474108 693636 474109 693700
rect 474043 693635 474109 693636
rect 521331 693700 521397 693701
rect 521331 693636 521332 693700
rect 521396 693636 521397 693700
rect 521331 693635 521397 693636
rect 424182 693230 424978 693290
rect 433934 692610 433994 693635
rect 434486 692610 434546 693635
rect 473494 693290 473554 693635
rect 474046 693290 474106 693635
rect 473494 693230 474106 693290
rect 539550 692698 539610 694043
rect 543595 693972 543661 693973
rect 543595 693908 543596 693972
rect 543660 693970 543661 693972
rect 543779 693972 543845 693973
rect 543779 693970 543780 693972
rect 543660 693910 543780 693970
rect 543660 693908 543661 693910
rect 543595 693907 543661 693908
rect 543779 693908 543780 693910
rect 543844 693908 543845 693972
rect 562915 693972 562981 693973
rect 543779 693907 543845 693908
rect 550590 693910 550834 693970
rect 549115 693836 549181 693837
rect 549115 693772 549116 693836
rect 549180 693772 549181 693836
rect 549115 693771 549181 693772
rect 549118 692698 549178 693771
rect 550590 693701 550650 693910
rect 550774 693701 550834 693910
rect 562915 693908 562916 693972
rect 562980 693970 562981 693972
rect 563099 693972 563165 693973
rect 563099 693970 563100 693972
rect 562980 693910 563100 693970
rect 562980 693908 562981 693910
rect 562915 693907 562981 693908
rect 563099 693908 563100 693910
rect 563164 693908 563165 693972
rect 563099 693907 563165 693908
rect 550587 693700 550653 693701
rect 550587 693636 550588 693700
rect 550652 693636 550653 693700
rect 550587 693635 550653 693636
rect 550771 693700 550837 693701
rect 550771 693636 550772 693700
rect 550836 693636 550837 693700
rect 550771 693635 550837 693636
rect 558867 693700 558933 693701
rect 558867 693636 558868 693700
rect 558932 693636 558933 693700
rect 558867 693635 558933 693636
rect 558870 692698 558930 693635
rect 565675 693428 565741 693429
rect 565675 693364 565676 693428
rect 565740 693364 565741 693428
rect 565675 693363 565741 693364
rect 565678 692698 565738 693363
rect 433934 692550 434546 692610
rect 162902 691870 163882 691930
rect 4404 689818 4586 690054
rect 4822 689818 5004 690054
rect 4404 689734 5004 689818
rect 4404 689498 4586 689734
rect 4822 689498 5004 689734
rect 4404 654054 5004 689498
rect 4404 653818 4586 654054
rect 4822 653818 5004 654054
rect 4404 653734 5004 653818
rect 4404 653498 4586 653734
rect 4822 653498 5004 653734
rect 4404 618054 5004 653498
rect 4404 617818 4586 618054
rect 4822 617818 5004 618054
rect 4404 617734 5004 617818
rect 4404 617498 4586 617734
rect 4822 617498 5004 617734
rect 4404 582054 5004 617498
rect 4404 581818 4586 582054
rect 4822 581818 5004 582054
rect 4404 581734 5004 581818
rect 4404 581498 4586 581734
rect 4822 581498 5004 581734
rect 4404 546054 5004 581498
rect 4404 545818 4586 546054
rect 4822 545818 5004 546054
rect 4404 545734 5004 545818
rect 4404 545498 4586 545734
rect 4822 545498 5004 545734
rect 4404 510054 5004 545498
rect 4404 509818 4586 510054
rect 4822 509818 5004 510054
rect 4404 509734 5004 509818
rect 4404 509498 4586 509734
rect 4822 509498 5004 509734
rect 4404 474054 5004 509498
rect 4404 473818 4586 474054
rect 4822 473818 5004 474054
rect 4404 473734 5004 473818
rect 4404 473498 4586 473734
rect 4822 473498 5004 473734
rect 4404 438054 5004 473498
rect 4404 437818 4586 438054
rect 4822 437818 5004 438054
rect 4404 437734 5004 437818
rect 4404 437498 4586 437734
rect 4822 437498 5004 437734
rect 4404 402054 5004 437498
rect 4404 401818 4586 402054
rect 4822 401818 5004 402054
rect 4404 401734 5004 401818
rect 4404 401498 4586 401734
rect 4822 401498 5004 401734
rect 4404 366054 5004 401498
rect 4404 365818 4586 366054
rect 4822 365818 5004 366054
rect 4404 365734 5004 365818
rect 4404 365498 4586 365734
rect 4822 365498 5004 365734
rect 4404 330054 5004 365498
rect 4404 329818 4586 330054
rect 4822 329818 5004 330054
rect 4404 329734 5004 329818
rect 4404 329498 4586 329734
rect 4822 329498 5004 329734
rect 4404 294054 5004 329498
rect 4404 293818 4586 294054
rect 4822 293818 5004 294054
rect 4404 293734 5004 293818
rect 4404 293498 4586 293734
rect 4822 293498 5004 293734
rect 4404 258054 5004 293498
rect 4404 257818 4586 258054
rect 4822 257818 5004 258054
rect 4404 257734 5004 257818
rect 4404 257498 4586 257734
rect 4822 257498 5004 257734
rect 4404 222054 5004 257498
rect 4404 221818 4586 222054
rect 4822 221818 5004 222054
rect 4404 221734 5004 221818
rect 4404 221498 4586 221734
rect 4822 221498 5004 221734
rect 4404 186054 5004 221498
rect 4404 185818 4586 186054
rect 4822 185818 5004 186054
rect 4404 185734 5004 185818
rect 4404 185498 4586 185734
rect 4822 185498 5004 185734
rect 4404 150054 5004 185498
rect 4404 149818 4586 150054
rect 4822 149818 5004 150054
rect 4404 149734 5004 149818
rect 4404 149498 4586 149734
rect 4822 149498 5004 149734
rect 4404 114054 5004 149498
rect 4404 113818 4586 114054
rect 4822 113818 5004 114054
rect 4404 113734 5004 113818
rect 4404 113498 4586 113734
rect 4822 113498 5004 113734
rect 4404 78054 5004 113498
rect 4404 77818 4586 78054
rect 4822 77818 5004 78054
rect 4404 77734 5004 77818
rect 4404 77498 4586 77734
rect 4822 77498 5004 77734
rect 4404 42054 5004 77498
rect 4404 41818 4586 42054
rect 4822 41818 5004 42054
rect 4404 41734 5004 41818
rect 4404 41498 4586 41734
rect 4822 41498 5004 41734
rect 4404 6054 5004 41498
rect 4404 5818 4586 6054
rect 4822 5818 5004 6054
rect 580404 690054 581004 706162
rect 587200 706718 587800 706740
rect 587200 706482 587382 706718
rect 587618 706482 587800 706718
rect 587200 706398 587800 706482
rect 587200 706162 587382 706398
rect 587618 706162 587800 706398
rect 586260 705778 586860 705800
rect 586260 705542 586442 705778
rect 586678 705542 586860 705778
rect 586260 705458 586860 705542
rect 586260 705222 586442 705458
rect 586678 705222 586860 705458
rect 580404 689818 580586 690054
rect 580822 689818 581004 690054
rect 580404 689734 581004 689818
rect 580404 689498 580586 689734
rect 580822 689498 581004 689734
rect 580404 654054 581004 689498
rect 580404 653818 580586 654054
rect 580822 653818 581004 654054
rect 580404 653734 581004 653818
rect 580404 653498 580586 653734
rect 580822 653498 581004 653734
rect 580404 618054 581004 653498
rect 580404 617818 580586 618054
rect 580822 617818 581004 618054
rect 580404 617734 581004 617818
rect 580404 617498 580586 617734
rect 580822 617498 581004 617734
rect 580404 582054 581004 617498
rect 580404 581818 580586 582054
rect 580822 581818 581004 582054
rect 580404 581734 581004 581818
rect 580404 581498 580586 581734
rect 580822 581498 581004 581734
rect 580404 546054 581004 581498
rect 580404 545818 580586 546054
rect 580822 545818 581004 546054
rect 580404 545734 581004 545818
rect 580404 545498 580586 545734
rect 580822 545498 581004 545734
rect 580404 510054 581004 545498
rect 580404 509818 580586 510054
rect 580822 509818 581004 510054
rect 580404 509734 581004 509818
rect 580404 509498 580586 509734
rect 580822 509498 581004 509734
rect 580404 474054 581004 509498
rect 580404 473818 580586 474054
rect 580822 473818 581004 474054
rect 580404 473734 581004 473818
rect 580404 473498 580586 473734
rect 580822 473498 581004 473734
rect 580404 438054 581004 473498
rect 580404 437818 580586 438054
rect 580822 437818 581004 438054
rect 580404 437734 581004 437818
rect 580404 437498 580586 437734
rect 580822 437498 581004 437734
rect 580404 402054 581004 437498
rect 580404 401818 580586 402054
rect 580822 401818 581004 402054
rect 580404 401734 581004 401818
rect 580404 401498 580586 401734
rect 580822 401498 581004 401734
rect 580404 366054 581004 401498
rect 580404 365818 580586 366054
rect 580822 365818 581004 366054
rect 580404 365734 581004 365818
rect 580404 365498 580586 365734
rect 580822 365498 581004 365734
rect 580404 330054 581004 365498
rect 580404 329818 580586 330054
rect 580822 329818 581004 330054
rect 580404 329734 581004 329818
rect 580404 329498 580586 329734
rect 580822 329498 581004 329734
rect 580404 294054 581004 329498
rect 580404 293818 580586 294054
rect 580822 293818 581004 294054
rect 580404 293734 581004 293818
rect 580404 293498 580586 293734
rect 580822 293498 581004 293734
rect 580404 258054 581004 293498
rect 580404 257818 580586 258054
rect 580822 257818 581004 258054
rect 580404 257734 581004 257818
rect 580404 257498 580586 257734
rect 580822 257498 581004 257734
rect 580404 222054 581004 257498
rect 580404 221818 580586 222054
rect 580822 221818 581004 222054
rect 580404 221734 581004 221818
rect 580404 221498 580586 221734
rect 580822 221498 581004 221734
rect 580404 186054 581004 221498
rect 580404 185818 580586 186054
rect 580822 185818 581004 186054
rect 580404 185734 581004 185818
rect 580404 185498 580586 185734
rect 580822 185498 581004 185734
rect 580404 150054 581004 185498
rect 580404 149818 580586 150054
rect 580822 149818 581004 150054
rect 580404 149734 581004 149818
rect 580404 149498 580586 149734
rect 580822 149498 581004 149734
rect 580404 114054 581004 149498
rect 580404 113818 580586 114054
rect 580822 113818 581004 114054
rect 580404 113734 581004 113818
rect 580404 113498 580586 113734
rect 580822 113498 581004 113734
rect 580404 78054 581004 113498
rect 580404 77818 580586 78054
rect 580822 77818 581004 78054
rect 580404 77734 581004 77818
rect 580404 77498 580586 77734
rect 580822 77498 581004 77734
rect 580404 42054 581004 77498
rect 580404 41818 580586 42054
rect 580822 41818 581004 42054
rect 580404 41734 581004 41818
rect 580404 41498 580586 41734
rect 580822 41498 581004 41734
rect 580404 6054 581004 41498
rect 18804 6016 19404 6048
rect 4404 5734 5004 5818
rect 4404 5498 4586 5734
rect 4822 5498 5004 5734
rect -3876 -2462 -3694 -2226
rect -3458 -2462 -3276 -2226
rect -3876 -2546 -3276 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 -3276 -2546
rect -3876 -2804 -3276 -2782
rect 4404 -2226 5004 5498
rect 4404 -2462 4586 -2226
rect 4822 -2462 5004 -2226
rect 4404 -2546 5004 -2462
rect 4404 -2782 4586 -2546
rect 4822 -2782 5004 -2546
rect -4816 -3402 -4634 -3166
rect -4398 -3402 -4216 -3166
rect -4816 -3486 -4216 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 -4216 -3486
rect -4816 -3744 -4216 -3722
rect 4404 -3744 5004 -2782
rect -5756 -4342 -5574 -4106
rect -5338 -4342 -5156 -4106
rect -5756 -4426 -5156 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 -5156 -4426
rect -5756 -4684 -5156 -4662
rect 8004 -4106 8604 6000
rect 8004 -4342 8186 -4106
rect 8422 -4342 8604 -4106
rect 8004 -4426 8604 -4342
rect 8004 -4662 8186 -4426
rect 8422 -4662 8604 -4426
rect -6696 -5282 -6514 -5046
rect -6278 -5282 -6096 -5046
rect -6696 -5366 -6096 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 -6096 -5366
rect -6696 -5624 -6096 -5602
rect 8004 -5624 8604 -4662
rect -7636 -6222 -7454 -5986
rect -7218 -6222 -7036 -5986
rect -7636 -6306 -7036 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 -7036 -6306
rect -7636 -6564 -7036 -6542
rect 11604 -5986 12204 6000
rect 18804 5952 18832 6016
rect 18896 5952 18912 6016
rect 18976 5952 18992 6016
rect 19056 5952 19072 6016
rect 19136 5952 19152 6016
rect 19216 5952 19232 6016
rect 19296 5952 19312 6016
rect 19376 5952 19404 6016
rect 18804 4928 19404 5952
rect 18804 4864 18832 4928
rect 18896 4864 18912 4928
rect 18976 4864 18992 4928
rect 19056 4864 19072 4928
rect 19136 4864 19152 4928
rect 19216 4864 19232 4928
rect 19296 4864 19312 4928
rect 19376 4864 19404 4928
rect 18804 3840 19404 4864
rect 18804 3776 18832 3840
rect 18896 3776 18912 3840
rect 18976 3776 18992 3840
rect 19056 3776 19072 3840
rect 19136 3776 19152 3840
rect 19216 3776 19232 3840
rect 19296 3776 19312 3840
rect 19376 3776 19404 3840
rect 18804 2752 19404 3776
rect 18804 2688 18832 2752
rect 18896 2688 18912 2752
rect 18976 2688 18992 2752
rect 19056 2688 19072 2752
rect 19136 2688 19152 2752
rect 19216 2688 19232 2752
rect 19296 2688 19312 2752
rect 19376 2688 19404 2752
rect 18804 -1286 19404 2688
rect 18804 -1522 18986 -1286
rect 19222 -1522 19404 -1286
rect 18804 -1606 19404 -1522
rect 18804 -1842 18986 -1606
rect 19222 -1842 19404 -1606
rect 18804 -1864 19404 -1842
rect 22404 -3166 23004 6000
rect 22404 -3402 22586 -3166
rect 22822 -3402 23004 -3166
rect 22404 -3486 23004 -3402
rect 22404 -3722 22586 -3486
rect 22822 -3722 23004 -3486
rect 22404 -3744 23004 -3722
rect 26004 -5046 26604 6000
rect 26004 -5282 26186 -5046
rect 26422 -5282 26604 -5046
rect 26004 -5366 26604 -5282
rect 26004 -5602 26186 -5366
rect 26422 -5602 26604 -5366
rect 26004 -5624 26604 -5602
rect 11604 -6222 11786 -5986
rect 12022 -6222 12204 -5986
rect 11604 -6306 12204 -6222
rect 11604 -6542 11786 -6306
rect 12022 -6542 12204 -6306
rect -8576 -7162 -8394 -6926
rect -8158 -7162 -7976 -6926
rect -8576 -7246 -7976 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 -7976 -7246
rect -8576 -7504 -7976 -7482
rect 11604 -7504 12204 -6542
rect 29604 -6926 30204 6000
rect 36804 5472 37404 6048
rect 54804 6016 55404 6048
rect 36804 5408 36832 5472
rect 36896 5408 36912 5472
rect 36976 5408 36992 5472
rect 37056 5408 37072 5472
rect 37136 5408 37152 5472
rect 37216 5408 37232 5472
rect 37296 5408 37312 5472
rect 37376 5408 37404 5472
rect 36804 4384 37404 5408
rect 36804 4320 36832 4384
rect 36896 4320 36912 4384
rect 36976 4320 36992 4384
rect 37056 4320 37072 4384
rect 37136 4320 37152 4384
rect 37216 4320 37232 4384
rect 37296 4320 37312 4384
rect 37376 4320 37404 4384
rect 36804 3296 37404 4320
rect 36804 3232 36832 3296
rect 36896 3232 36912 3296
rect 36976 3232 36992 3296
rect 37056 3232 37072 3296
rect 37136 3232 37152 3296
rect 37216 3232 37232 3296
rect 37296 3232 37312 3296
rect 37376 3232 37404 3296
rect 36804 2406 37404 3232
rect 36804 2208 36986 2406
rect 37222 2208 37404 2406
rect 36804 2144 36832 2208
rect 36896 2144 36912 2208
rect 36976 2170 36986 2208
rect 37222 2170 37232 2208
rect 36976 2144 36992 2170
rect 37056 2144 37072 2170
rect 37136 2144 37152 2170
rect 37216 2144 37232 2170
rect 37296 2144 37312 2208
rect 37376 2144 37404 2208
rect 36804 2086 37404 2144
rect 36804 1850 36986 2086
rect 37222 1850 37404 2086
rect 36804 -346 37404 1850
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1864 37404 -902
rect 40404 -2226 41004 6000
rect 40404 -2462 40586 -2226
rect 40822 -2462 41004 -2226
rect 40404 -2546 41004 -2462
rect 40404 -2782 40586 -2546
rect 40822 -2782 41004 -2546
rect 40404 -3744 41004 -2782
rect 44004 -4106 44604 6000
rect 44004 -4342 44186 -4106
rect 44422 -4342 44604 -4106
rect 44004 -4426 44604 -4342
rect 44004 -4662 44186 -4426
rect 44422 -4662 44604 -4426
rect 44004 -5624 44604 -4662
rect 29604 -7162 29786 -6926
rect 30022 -7162 30204 -6926
rect 29604 -7246 30204 -7162
rect 29604 -7482 29786 -7246
rect 30022 -7482 30204 -7246
rect 29604 -7504 30204 -7482
rect 47604 -5986 48204 6000
rect 54804 5952 54832 6016
rect 54896 5952 54912 6016
rect 54976 5952 54992 6016
rect 55056 5952 55072 6016
rect 55136 5952 55152 6016
rect 55216 5952 55232 6016
rect 55296 5952 55312 6016
rect 55376 5952 55404 6016
rect 54804 4928 55404 5952
rect 54804 4864 54832 4928
rect 54896 4864 54912 4928
rect 54976 4864 54992 4928
rect 55056 4864 55072 4928
rect 55136 4864 55152 4928
rect 55216 4864 55232 4928
rect 55296 4864 55312 4928
rect 55376 4864 55404 4928
rect 54804 3840 55404 4864
rect 54804 3776 54832 3840
rect 54896 3776 54912 3840
rect 54976 3776 54992 3840
rect 55056 3776 55072 3840
rect 55136 3776 55152 3840
rect 55216 3776 55232 3840
rect 55296 3776 55312 3840
rect 55376 3776 55404 3840
rect 54804 2752 55404 3776
rect 54804 2688 54832 2752
rect 54896 2688 54912 2752
rect 54976 2688 54992 2752
rect 55056 2688 55072 2752
rect 55136 2688 55152 2752
rect 55216 2688 55232 2752
rect 55296 2688 55312 2752
rect 55376 2688 55404 2752
rect 54804 -1286 55404 2688
rect 54804 -1522 54986 -1286
rect 55222 -1522 55404 -1286
rect 54804 -1606 55404 -1522
rect 54804 -1842 54986 -1606
rect 55222 -1842 55404 -1606
rect 54804 -1864 55404 -1842
rect 58404 -3166 59004 6000
rect 58404 -3402 58586 -3166
rect 58822 -3402 59004 -3166
rect 58404 -3486 59004 -3402
rect 58404 -3722 58586 -3486
rect 58822 -3722 59004 -3486
rect 58404 -3744 59004 -3722
rect 62004 -5046 62604 6000
rect 62004 -5282 62186 -5046
rect 62422 -5282 62604 -5046
rect 62004 -5366 62604 -5282
rect 62004 -5602 62186 -5366
rect 62422 -5602 62604 -5366
rect 62004 -5624 62604 -5602
rect 47604 -6222 47786 -5986
rect 48022 -6222 48204 -5986
rect 47604 -6306 48204 -6222
rect 47604 -6542 47786 -6306
rect 48022 -6542 48204 -6306
rect 47604 -7504 48204 -6542
rect 65604 -6926 66204 6000
rect 72804 5472 73404 6048
rect 90804 6016 91404 6048
rect 72804 5408 72832 5472
rect 72896 5408 72912 5472
rect 72976 5408 72992 5472
rect 73056 5408 73072 5472
rect 73136 5408 73152 5472
rect 73216 5408 73232 5472
rect 73296 5408 73312 5472
rect 73376 5408 73404 5472
rect 72804 4384 73404 5408
rect 72804 4320 72832 4384
rect 72896 4320 72912 4384
rect 72976 4320 72992 4384
rect 73056 4320 73072 4384
rect 73136 4320 73152 4384
rect 73216 4320 73232 4384
rect 73296 4320 73312 4384
rect 73376 4320 73404 4384
rect 72804 3296 73404 4320
rect 72804 3232 72832 3296
rect 72896 3232 72912 3296
rect 72976 3232 72992 3296
rect 73056 3232 73072 3296
rect 73136 3232 73152 3296
rect 73216 3232 73232 3296
rect 73296 3232 73312 3296
rect 73376 3232 73404 3296
rect 72804 2406 73404 3232
rect 72804 2208 72986 2406
rect 73222 2208 73404 2406
rect 72804 2144 72832 2208
rect 72896 2144 72912 2208
rect 72976 2170 72986 2208
rect 73222 2170 73232 2208
rect 72976 2144 72992 2170
rect 73056 2144 73072 2170
rect 73136 2144 73152 2170
rect 73216 2144 73232 2170
rect 73296 2144 73312 2208
rect 73376 2144 73404 2208
rect 72804 2086 73404 2144
rect 72804 1850 72986 2086
rect 73222 1850 73404 2086
rect 72804 -346 73404 1850
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1864 73404 -902
rect 76404 -2226 77004 6000
rect 76404 -2462 76586 -2226
rect 76822 -2462 77004 -2226
rect 76404 -2546 77004 -2462
rect 76404 -2782 76586 -2546
rect 76822 -2782 77004 -2546
rect 76404 -3744 77004 -2782
rect 80004 -4106 80604 6000
rect 80004 -4342 80186 -4106
rect 80422 -4342 80604 -4106
rect 80004 -4426 80604 -4342
rect 80004 -4662 80186 -4426
rect 80422 -4662 80604 -4426
rect 80004 -5624 80604 -4662
rect 65604 -7162 65786 -6926
rect 66022 -7162 66204 -6926
rect 65604 -7246 66204 -7162
rect 65604 -7482 65786 -7246
rect 66022 -7482 66204 -7246
rect 65604 -7504 66204 -7482
rect 83604 -5986 84204 6000
rect 90804 5952 90832 6016
rect 90896 5952 90912 6016
rect 90976 5952 90992 6016
rect 91056 5952 91072 6016
rect 91136 5952 91152 6016
rect 91216 5952 91232 6016
rect 91296 5952 91312 6016
rect 91376 5952 91404 6016
rect 90804 4928 91404 5952
rect 90804 4864 90832 4928
rect 90896 4864 90912 4928
rect 90976 4864 90992 4928
rect 91056 4864 91072 4928
rect 91136 4864 91152 4928
rect 91216 4864 91232 4928
rect 91296 4864 91312 4928
rect 91376 4864 91404 4928
rect 90804 3840 91404 4864
rect 90804 3776 90832 3840
rect 90896 3776 90912 3840
rect 90976 3776 90992 3840
rect 91056 3776 91072 3840
rect 91136 3776 91152 3840
rect 91216 3776 91232 3840
rect 91296 3776 91312 3840
rect 91376 3776 91404 3840
rect 90804 2752 91404 3776
rect 90804 2688 90832 2752
rect 90896 2688 90912 2752
rect 90976 2688 90992 2752
rect 91056 2688 91072 2752
rect 91136 2688 91152 2752
rect 91216 2688 91232 2752
rect 91296 2688 91312 2752
rect 91376 2688 91404 2752
rect 90804 -1286 91404 2688
rect 90804 -1522 90986 -1286
rect 91222 -1522 91404 -1286
rect 90804 -1606 91404 -1522
rect 90804 -1842 90986 -1606
rect 91222 -1842 91404 -1606
rect 90804 -1864 91404 -1842
rect 94404 -3166 95004 6000
rect 94404 -3402 94586 -3166
rect 94822 -3402 95004 -3166
rect 94404 -3486 95004 -3402
rect 94404 -3722 94586 -3486
rect 94822 -3722 95004 -3486
rect 94404 -3744 95004 -3722
rect 98004 -5046 98604 6000
rect 98004 -5282 98186 -5046
rect 98422 -5282 98604 -5046
rect 98004 -5366 98604 -5282
rect 98004 -5602 98186 -5366
rect 98422 -5602 98604 -5366
rect 98004 -5624 98604 -5602
rect 83604 -6222 83786 -5986
rect 84022 -6222 84204 -5986
rect 83604 -6306 84204 -6222
rect 83604 -6542 83786 -6306
rect 84022 -6542 84204 -6306
rect 83604 -7504 84204 -6542
rect 101604 -6926 102204 6000
rect 108804 5472 109404 6048
rect 126804 6016 127404 6048
rect 108804 5408 108832 5472
rect 108896 5408 108912 5472
rect 108976 5408 108992 5472
rect 109056 5408 109072 5472
rect 109136 5408 109152 5472
rect 109216 5408 109232 5472
rect 109296 5408 109312 5472
rect 109376 5408 109404 5472
rect 108804 4384 109404 5408
rect 108804 4320 108832 4384
rect 108896 4320 108912 4384
rect 108976 4320 108992 4384
rect 109056 4320 109072 4384
rect 109136 4320 109152 4384
rect 109216 4320 109232 4384
rect 109296 4320 109312 4384
rect 109376 4320 109404 4384
rect 108804 3296 109404 4320
rect 108804 3232 108832 3296
rect 108896 3232 108912 3296
rect 108976 3232 108992 3296
rect 109056 3232 109072 3296
rect 109136 3232 109152 3296
rect 109216 3232 109232 3296
rect 109296 3232 109312 3296
rect 109376 3232 109404 3296
rect 108804 2406 109404 3232
rect 108804 2208 108986 2406
rect 109222 2208 109404 2406
rect 108804 2144 108832 2208
rect 108896 2144 108912 2208
rect 108976 2170 108986 2208
rect 109222 2170 109232 2208
rect 108976 2144 108992 2170
rect 109056 2144 109072 2170
rect 109136 2144 109152 2170
rect 109216 2144 109232 2170
rect 109296 2144 109312 2208
rect 109376 2144 109404 2208
rect 108804 2086 109404 2144
rect 108804 1850 108986 2086
rect 109222 1850 109404 2086
rect 108804 -346 109404 1850
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1864 109404 -902
rect 112404 -2226 113004 6000
rect 112404 -2462 112586 -2226
rect 112822 -2462 113004 -2226
rect 112404 -2546 113004 -2462
rect 112404 -2782 112586 -2546
rect 112822 -2782 113004 -2546
rect 112404 -3744 113004 -2782
rect 116004 -4106 116604 6000
rect 116004 -4342 116186 -4106
rect 116422 -4342 116604 -4106
rect 116004 -4426 116604 -4342
rect 116004 -4662 116186 -4426
rect 116422 -4662 116604 -4426
rect 116004 -5624 116604 -4662
rect 101604 -7162 101786 -6926
rect 102022 -7162 102204 -6926
rect 101604 -7246 102204 -7162
rect 101604 -7482 101786 -7246
rect 102022 -7482 102204 -7246
rect 101604 -7504 102204 -7482
rect 119604 -5986 120204 6000
rect 126804 5952 126832 6016
rect 126896 5952 126912 6016
rect 126976 5952 126992 6016
rect 127056 5952 127072 6016
rect 127136 5952 127152 6016
rect 127216 5952 127232 6016
rect 127296 5952 127312 6016
rect 127376 5952 127404 6016
rect 126804 4928 127404 5952
rect 126804 4864 126832 4928
rect 126896 4864 126912 4928
rect 126976 4864 126992 4928
rect 127056 4864 127072 4928
rect 127136 4864 127152 4928
rect 127216 4864 127232 4928
rect 127296 4864 127312 4928
rect 127376 4864 127404 4928
rect 126804 3840 127404 4864
rect 126804 3776 126832 3840
rect 126896 3776 126912 3840
rect 126976 3776 126992 3840
rect 127056 3776 127072 3840
rect 127136 3776 127152 3840
rect 127216 3776 127232 3840
rect 127296 3776 127312 3840
rect 127376 3776 127404 3840
rect 126804 2752 127404 3776
rect 126804 2688 126832 2752
rect 126896 2688 126912 2752
rect 126976 2688 126992 2752
rect 127056 2688 127072 2752
rect 127136 2688 127152 2752
rect 127216 2688 127232 2752
rect 127296 2688 127312 2752
rect 127376 2688 127404 2752
rect 126804 -1286 127404 2688
rect 126804 -1522 126986 -1286
rect 127222 -1522 127404 -1286
rect 126804 -1606 127404 -1522
rect 126804 -1842 126986 -1606
rect 127222 -1842 127404 -1606
rect 126804 -1864 127404 -1842
rect 130404 -3166 131004 6000
rect 130404 -3402 130586 -3166
rect 130822 -3402 131004 -3166
rect 130404 -3486 131004 -3402
rect 130404 -3722 130586 -3486
rect 130822 -3722 131004 -3486
rect 130404 -3744 131004 -3722
rect 134004 -5046 134604 6000
rect 134004 -5282 134186 -5046
rect 134422 -5282 134604 -5046
rect 134004 -5366 134604 -5282
rect 134004 -5602 134186 -5366
rect 134422 -5602 134604 -5366
rect 134004 -5624 134604 -5602
rect 119604 -6222 119786 -5986
rect 120022 -6222 120204 -5986
rect 119604 -6306 120204 -6222
rect 119604 -6542 119786 -6306
rect 120022 -6542 120204 -6306
rect 119604 -7504 120204 -6542
rect 137604 -6926 138204 6000
rect 144804 5472 145404 6048
rect 162804 6016 163404 6048
rect 144804 5408 144832 5472
rect 144896 5408 144912 5472
rect 144976 5408 144992 5472
rect 145056 5408 145072 5472
rect 145136 5408 145152 5472
rect 145216 5408 145232 5472
rect 145296 5408 145312 5472
rect 145376 5408 145404 5472
rect 144804 4384 145404 5408
rect 144804 4320 144832 4384
rect 144896 4320 144912 4384
rect 144976 4320 144992 4384
rect 145056 4320 145072 4384
rect 145136 4320 145152 4384
rect 145216 4320 145232 4384
rect 145296 4320 145312 4384
rect 145376 4320 145404 4384
rect 144804 3296 145404 4320
rect 144804 3232 144832 3296
rect 144896 3232 144912 3296
rect 144976 3232 144992 3296
rect 145056 3232 145072 3296
rect 145136 3232 145152 3296
rect 145216 3232 145232 3296
rect 145296 3232 145312 3296
rect 145376 3232 145404 3296
rect 144804 2406 145404 3232
rect 144804 2208 144986 2406
rect 145222 2208 145404 2406
rect 144804 2144 144832 2208
rect 144896 2144 144912 2208
rect 144976 2170 144986 2208
rect 145222 2170 145232 2208
rect 144976 2144 144992 2170
rect 145056 2144 145072 2170
rect 145136 2144 145152 2170
rect 145216 2144 145232 2170
rect 145296 2144 145312 2208
rect 145376 2144 145404 2208
rect 144804 2086 145404 2144
rect 144804 1850 144986 2086
rect 145222 1850 145404 2086
rect 144804 -346 145404 1850
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1864 145404 -902
rect 148404 -2226 149004 6000
rect 148404 -2462 148586 -2226
rect 148822 -2462 149004 -2226
rect 148404 -2546 149004 -2462
rect 148404 -2782 148586 -2546
rect 148822 -2782 149004 -2546
rect 148404 -3744 149004 -2782
rect 152004 -4106 152604 6000
rect 152004 -4342 152186 -4106
rect 152422 -4342 152604 -4106
rect 152004 -4426 152604 -4342
rect 152004 -4662 152186 -4426
rect 152422 -4662 152604 -4426
rect 152004 -5624 152604 -4662
rect 137604 -7162 137786 -6926
rect 138022 -7162 138204 -6926
rect 137604 -7246 138204 -7162
rect 137604 -7482 137786 -7246
rect 138022 -7482 138204 -7246
rect 137604 -7504 138204 -7482
rect 155604 -5986 156204 6000
rect 162804 5952 162832 6016
rect 162896 5952 162912 6016
rect 162976 5952 162992 6016
rect 163056 5952 163072 6016
rect 163136 5952 163152 6016
rect 163216 5952 163232 6016
rect 163296 5952 163312 6016
rect 163376 5952 163404 6016
rect 162804 4928 163404 5952
rect 162804 4864 162832 4928
rect 162896 4864 162912 4928
rect 162976 4864 162992 4928
rect 163056 4864 163072 4928
rect 163136 4864 163152 4928
rect 163216 4864 163232 4928
rect 163296 4864 163312 4928
rect 163376 4864 163404 4928
rect 162804 3840 163404 4864
rect 162804 3776 162832 3840
rect 162896 3776 162912 3840
rect 162976 3776 162992 3840
rect 163056 3776 163072 3840
rect 163136 3776 163152 3840
rect 163216 3776 163232 3840
rect 163296 3776 163312 3840
rect 163376 3776 163404 3840
rect 162804 2752 163404 3776
rect 162804 2688 162832 2752
rect 162896 2688 162912 2752
rect 162976 2688 162992 2752
rect 163056 2688 163072 2752
rect 163136 2688 163152 2752
rect 163216 2688 163232 2752
rect 163296 2688 163312 2752
rect 163376 2688 163404 2752
rect 162804 -1286 163404 2688
rect 162804 -1522 162986 -1286
rect 163222 -1522 163404 -1286
rect 162804 -1606 163404 -1522
rect 162804 -1842 162986 -1606
rect 163222 -1842 163404 -1606
rect 162804 -1864 163404 -1842
rect 166404 -3166 167004 6000
rect 166404 -3402 166586 -3166
rect 166822 -3402 167004 -3166
rect 166404 -3486 167004 -3402
rect 166404 -3722 166586 -3486
rect 166822 -3722 167004 -3486
rect 166404 -3744 167004 -3722
rect 170004 -5046 170604 6000
rect 170004 -5282 170186 -5046
rect 170422 -5282 170604 -5046
rect 170004 -5366 170604 -5282
rect 170004 -5602 170186 -5366
rect 170422 -5602 170604 -5366
rect 170004 -5624 170604 -5602
rect 155604 -6222 155786 -5986
rect 156022 -6222 156204 -5986
rect 155604 -6306 156204 -6222
rect 155604 -6542 155786 -6306
rect 156022 -6542 156204 -6306
rect 155604 -7504 156204 -6542
rect 173604 -6926 174204 6000
rect 180804 5472 181404 6048
rect 198804 6016 199404 6048
rect 180804 5408 180832 5472
rect 180896 5408 180912 5472
rect 180976 5408 180992 5472
rect 181056 5408 181072 5472
rect 181136 5408 181152 5472
rect 181216 5408 181232 5472
rect 181296 5408 181312 5472
rect 181376 5408 181404 5472
rect 180804 4384 181404 5408
rect 180804 4320 180832 4384
rect 180896 4320 180912 4384
rect 180976 4320 180992 4384
rect 181056 4320 181072 4384
rect 181136 4320 181152 4384
rect 181216 4320 181232 4384
rect 181296 4320 181312 4384
rect 181376 4320 181404 4384
rect 180804 3296 181404 4320
rect 180804 3232 180832 3296
rect 180896 3232 180912 3296
rect 180976 3232 180992 3296
rect 181056 3232 181072 3296
rect 181136 3232 181152 3296
rect 181216 3232 181232 3296
rect 181296 3232 181312 3296
rect 181376 3232 181404 3296
rect 180804 2406 181404 3232
rect 180804 2208 180986 2406
rect 181222 2208 181404 2406
rect 180804 2144 180832 2208
rect 180896 2144 180912 2208
rect 180976 2170 180986 2208
rect 181222 2170 181232 2208
rect 180976 2144 180992 2170
rect 181056 2144 181072 2170
rect 181136 2144 181152 2170
rect 181216 2144 181232 2170
rect 181296 2144 181312 2208
rect 181376 2144 181404 2208
rect 180804 2086 181404 2144
rect 180804 1850 180986 2086
rect 181222 1850 181404 2086
rect 180804 -346 181404 1850
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1864 181404 -902
rect 184404 -2226 185004 6000
rect 184404 -2462 184586 -2226
rect 184822 -2462 185004 -2226
rect 184404 -2546 185004 -2462
rect 184404 -2782 184586 -2546
rect 184822 -2782 185004 -2546
rect 184404 -3744 185004 -2782
rect 188004 -4106 188604 6000
rect 188004 -4342 188186 -4106
rect 188422 -4342 188604 -4106
rect 188004 -4426 188604 -4342
rect 188004 -4662 188186 -4426
rect 188422 -4662 188604 -4426
rect 188004 -5624 188604 -4662
rect 173604 -7162 173786 -6926
rect 174022 -7162 174204 -6926
rect 173604 -7246 174204 -7162
rect 173604 -7482 173786 -7246
rect 174022 -7482 174204 -7246
rect 173604 -7504 174204 -7482
rect 191604 -5986 192204 6000
rect 198804 5952 198832 6016
rect 198896 5952 198912 6016
rect 198976 5952 198992 6016
rect 199056 5952 199072 6016
rect 199136 5952 199152 6016
rect 199216 5952 199232 6016
rect 199296 5952 199312 6016
rect 199376 5952 199404 6016
rect 198804 4928 199404 5952
rect 198804 4864 198832 4928
rect 198896 4864 198912 4928
rect 198976 4864 198992 4928
rect 199056 4864 199072 4928
rect 199136 4864 199152 4928
rect 199216 4864 199232 4928
rect 199296 4864 199312 4928
rect 199376 4864 199404 4928
rect 198804 3840 199404 4864
rect 198804 3776 198832 3840
rect 198896 3776 198912 3840
rect 198976 3776 198992 3840
rect 199056 3776 199072 3840
rect 199136 3776 199152 3840
rect 199216 3776 199232 3840
rect 199296 3776 199312 3840
rect 199376 3776 199404 3840
rect 198804 2752 199404 3776
rect 198804 2688 198832 2752
rect 198896 2688 198912 2752
rect 198976 2688 198992 2752
rect 199056 2688 199072 2752
rect 199136 2688 199152 2752
rect 199216 2688 199232 2752
rect 199296 2688 199312 2752
rect 199376 2688 199404 2752
rect 198804 -1286 199404 2688
rect 198804 -1522 198986 -1286
rect 199222 -1522 199404 -1286
rect 198804 -1606 199404 -1522
rect 198804 -1842 198986 -1606
rect 199222 -1842 199404 -1606
rect 198804 -1864 199404 -1842
rect 202404 -3166 203004 6000
rect 202404 -3402 202586 -3166
rect 202822 -3402 203004 -3166
rect 202404 -3486 203004 -3402
rect 202404 -3722 202586 -3486
rect 202822 -3722 203004 -3486
rect 202404 -3744 203004 -3722
rect 206004 -5046 206604 6000
rect 206004 -5282 206186 -5046
rect 206422 -5282 206604 -5046
rect 206004 -5366 206604 -5282
rect 206004 -5602 206186 -5366
rect 206422 -5602 206604 -5366
rect 206004 -5624 206604 -5602
rect 191604 -6222 191786 -5986
rect 192022 -6222 192204 -5986
rect 191604 -6306 192204 -6222
rect 191604 -6542 191786 -6306
rect 192022 -6542 192204 -6306
rect 191604 -7504 192204 -6542
rect 209604 -6926 210204 6000
rect 216804 5472 217404 6048
rect 234804 6016 235404 6048
rect 216804 5408 216832 5472
rect 216896 5408 216912 5472
rect 216976 5408 216992 5472
rect 217056 5408 217072 5472
rect 217136 5408 217152 5472
rect 217216 5408 217232 5472
rect 217296 5408 217312 5472
rect 217376 5408 217404 5472
rect 216804 4384 217404 5408
rect 216804 4320 216832 4384
rect 216896 4320 216912 4384
rect 216976 4320 216992 4384
rect 217056 4320 217072 4384
rect 217136 4320 217152 4384
rect 217216 4320 217232 4384
rect 217296 4320 217312 4384
rect 217376 4320 217404 4384
rect 216804 3296 217404 4320
rect 216804 3232 216832 3296
rect 216896 3232 216912 3296
rect 216976 3232 216992 3296
rect 217056 3232 217072 3296
rect 217136 3232 217152 3296
rect 217216 3232 217232 3296
rect 217296 3232 217312 3296
rect 217376 3232 217404 3296
rect 216804 2406 217404 3232
rect 216804 2208 216986 2406
rect 217222 2208 217404 2406
rect 216804 2144 216832 2208
rect 216896 2144 216912 2208
rect 216976 2170 216986 2208
rect 217222 2170 217232 2208
rect 216976 2144 216992 2170
rect 217056 2144 217072 2170
rect 217136 2144 217152 2170
rect 217216 2144 217232 2170
rect 217296 2144 217312 2208
rect 217376 2144 217404 2208
rect 216804 2086 217404 2144
rect 216804 1850 216986 2086
rect 217222 1850 217404 2086
rect 216804 -346 217404 1850
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1864 217404 -902
rect 220404 -2226 221004 6000
rect 220404 -2462 220586 -2226
rect 220822 -2462 221004 -2226
rect 220404 -2546 221004 -2462
rect 220404 -2782 220586 -2546
rect 220822 -2782 221004 -2546
rect 220404 -3744 221004 -2782
rect 224004 -4106 224604 6000
rect 224004 -4342 224186 -4106
rect 224422 -4342 224604 -4106
rect 224004 -4426 224604 -4342
rect 224004 -4662 224186 -4426
rect 224422 -4662 224604 -4426
rect 224004 -5624 224604 -4662
rect 209604 -7162 209786 -6926
rect 210022 -7162 210204 -6926
rect 209604 -7246 210204 -7162
rect 209604 -7482 209786 -7246
rect 210022 -7482 210204 -7246
rect 209604 -7504 210204 -7482
rect 227604 -5986 228204 6000
rect 234804 5952 234832 6016
rect 234896 5952 234912 6016
rect 234976 5952 234992 6016
rect 235056 5952 235072 6016
rect 235136 5952 235152 6016
rect 235216 5952 235232 6016
rect 235296 5952 235312 6016
rect 235376 5952 235404 6016
rect 234804 4928 235404 5952
rect 234804 4864 234832 4928
rect 234896 4864 234912 4928
rect 234976 4864 234992 4928
rect 235056 4864 235072 4928
rect 235136 4864 235152 4928
rect 235216 4864 235232 4928
rect 235296 4864 235312 4928
rect 235376 4864 235404 4928
rect 234804 3840 235404 4864
rect 234804 3776 234832 3840
rect 234896 3776 234912 3840
rect 234976 3776 234992 3840
rect 235056 3776 235072 3840
rect 235136 3776 235152 3840
rect 235216 3776 235232 3840
rect 235296 3776 235312 3840
rect 235376 3776 235404 3840
rect 234804 2752 235404 3776
rect 234804 2688 234832 2752
rect 234896 2688 234912 2752
rect 234976 2688 234992 2752
rect 235056 2688 235072 2752
rect 235136 2688 235152 2752
rect 235216 2688 235232 2752
rect 235296 2688 235312 2752
rect 235376 2688 235404 2752
rect 234804 -1286 235404 2688
rect 234804 -1522 234986 -1286
rect 235222 -1522 235404 -1286
rect 234804 -1606 235404 -1522
rect 234804 -1842 234986 -1606
rect 235222 -1842 235404 -1606
rect 234804 -1864 235404 -1842
rect 238404 -3166 239004 6000
rect 238404 -3402 238586 -3166
rect 238822 -3402 239004 -3166
rect 238404 -3486 239004 -3402
rect 238404 -3722 238586 -3486
rect 238822 -3722 239004 -3486
rect 238404 -3744 239004 -3722
rect 242004 -5046 242604 6000
rect 242004 -5282 242186 -5046
rect 242422 -5282 242604 -5046
rect 242004 -5366 242604 -5282
rect 242004 -5602 242186 -5366
rect 242422 -5602 242604 -5366
rect 242004 -5624 242604 -5602
rect 227604 -6222 227786 -5986
rect 228022 -6222 228204 -5986
rect 227604 -6306 228204 -6222
rect 227604 -6542 227786 -6306
rect 228022 -6542 228204 -6306
rect 227604 -7504 228204 -6542
rect 245604 -6926 246204 6000
rect 252804 5472 253404 6048
rect 270804 6016 271404 6048
rect 252804 5408 252832 5472
rect 252896 5408 252912 5472
rect 252976 5408 252992 5472
rect 253056 5408 253072 5472
rect 253136 5408 253152 5472
rect 253216 5408 253232 5472
rect 253296 5408 253312 5472
rect 253376 5408 253404 5472
rect 252804 4384 253404 5408
rect 252804 4320 252832 4384
rect 252896 4320 252912 4384
rect 252976 4320 252992 4384
rect 253056 4320 253072 4384
rect 253136 4320 253152 4384
rect 253216 4320 253232 4384
rect 253296 4320 253312 4384
rect 253376 4320 253404 4384
rect 252804 3296 253404 4320
rect 252804 3232 252832 3296
rect 252896 3232 252912 3296
rect 252976 3232 252992 3296
rect 253056 3232 253072 3296
rect 253136 3232 253152 3296
rect 253216 3232 253232 3296
rect 253296 3232 253312 3296
rect 253376 3232 253404 3296
rect 252804 2406 253404 3232
rect 252804 2208 252986 2406
rect 253222 2208 253404 2406
rect 252804 2144 252832 2208
rect 252896 2144 252912 2208
rect 252976 2170 252986 2208
rect 253222 2170 253232 2208
rect 252976 2144 252992 2170
rect 253056 2144 253072 2170
rect 253136 2144 253152 2170
rect 253216 2144 253232 2170
rect 253296 2144 253312 2208
rect 253376 2144 253404 2208
rect 252804 2086 253404 2144
rect 252804 1850 252986 2086
rect 253222 1850 253404 2086
rect 252804 -346 253404 1850
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1864 253404 -902
rect 256404 -2226 257004 6000
rect 256404 -2462 256586 -2226
rect 256822 -2462 257004 -2226
rect 256404 -2546 257004 -2462
rect 256404 -2782 256586 -2546
rect 256822 -2782 257004 -2546
rect 256404 -3744 257004 -2782
rect 260004 -4106 260604 6000
rect 260004 -4342 260186 -4106
rect 260422 -4342 260604 -4106
rect 260004 -4426 260604 -4342
rect 260004 -4662 260186 -4426
rect 260422 -4662 260604 -4426
rect 260004 -5624 260604 -4662
rect 245604 -7162 245786 -6926
rect 246022 -7162 246204 -6926
rect 245604 -7246 246204 -7162
rect 245604 -7482 245786 -7246
rect 246022 -7482 246204 -7246
rect 245604 -7504 246204 -7482
rect 263604 -5986 264204 6000
rect 270804 5952 270832 6016
rect 270896 5952 270912 6016
rect 270976 5952 270992 6016
rect 271056 5952 271072 6016
rect 271136 5952 271152 6016
rect 271216 5952 271232 6016
rect 271296 5952 271312 6016
rect 271376 5952 271404 6016
rect 270804 4928 271404 5952
rect 270804 4864 270832 4928
rect 270896 4864 270912 4928
rect 270976 4864 270992 4928
rect 271056 4864 271072 4928
rect 271136 4864 271152 4928
rect 271216 4864 271232 4928
rect 271296 4864 271312 4928
rect 271376 4864 271404 4928
rect 270804 3840 271404 4864
rect 270804 3776 270832 3840
rect 270896 3776 270912 3840
rect 270976 3776 270992 3840
rect 271056 3776 271072 3840
rect 271136 3776 271152 3840
rect 271216 3776 271232 3840
rect 271296 3776 271312 3840
rect 271376 3776 271404 3840
rect 270804 2752 271404 3776
rect 270804 2688 270832 2752
rect 270896 2688 270912 2752
rect 270976 2688 270992 2752
rect 271056 2688 271072 2752
rect 271136 2688 271152 2752
rect 271216 2688 271232 2752
rect 271296 2688 271312 2752
rect 271376 2688 271404 2752
rect 270804 -1286 271404 2688
rect 270804 -1522 270986 -1286
rect 271222 -1522 271404 -1286
rect 270804 -1606 271404 -1522
rect 270804 -1842 270986 -1606
rect 271222 -1842 271404 -1606
rect 270804 -1864 271404 -1842
rect 274404 -3166 275004 6000
rect 274404 -3402 274586 -3166
rect 274822 -3402 275004 -3166
rect 274404 -3486 275004 -3402
rect 274404 -3722 274586 -3486
rect 274822 -3722 275004 -3486
rect 274404 -3744 275004 -3722
rect 278004 -5046 278604 6000
rect 278004 -5282 278186 -5046
rect 278422 -5282 278604 -5046
rect 278004 -5366 278604 -5282
rect 278004 -5602 278186 -5366
rect 278422 -5602 278604 -5366
rect 278004 -5624 278604 -5602
rect 263604 -6222 263786 -5986
rect 264022 -6222 264204 -5986
rect 263604 -6306 264204 -6222
rect 263604 -6542 263786 -6306
rect 264022 -6542 264204 -6306
rect 263604 -7504 264204 -6542
rect 281604 -6926 282204 6000
rect 288804 5472 289404 6048
rect 306804 6016 307404 6048
rect 288804 5408 288832 5472
rect 288896 5408 288912 5472
rect 288976 5408 288992 5472
rect 289056 5408 289072 5472
rect 289136 5408 289152 5472
rect 289216 5408 289232 5472
rect 289296 5408 289312 5472
rect 289376 5408 289404 5472
rect 288804 4384 289404 5408
rect 288804 4320 288832 4384
rect 288896 4320 288912 4384
rect 288976 4320 288992 4384
rect 289056 4320 289072 4384
rect 289136 4320 289152 4384
rect 289216 4320 289232 4384
rect 289296 4320 289312 4384
rect 289376 4320 289404 4384
rect 288804 3296 289404 4320
rect 288804 3232 288832 3296
rect 288896 3232 288912 3296
rect 288976 3232 288992 3296
rect 289056 3232 289072 3296
rect 289136 3232 289152 3296
rect 289216 3232 289232 3296
rect 289296 3232 289312 3296
rect 289376 3232 289404 3296
rect 288804 2406 289404 3232
rect 288804 2208 288986 2406
rect 289222 2208 289404 2406
rect 288804 2144 288832 2208
rect 288896 2144 288912 2208
rect 288976 2170 288986 2208
rect 289222 2170 289232 2208
rect 288976 2144 288992 2170
rect 289056 2144 289072 2170
rect 289136 2144 289152 2170
rect 289216 2144 289232 2170
rect 289296 2144 289312 2208
rect 289376 2144 289404 2208
rect 288804 2086 289404 2144
rect 288804 1850 288986 2086
rect 289222 1850 289404 2086
rect 288804 -346 289404 1850
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1864 289404 -902
rect 292404 -2226 293004 6000
rect 292404 -2462 292586 -2226
rect 292822 -2462 293004 -2226
rect 292404 -2546 293004 -2462
rect 292404 -2782 292586 -2546
rect 292822 -2782 293004 -2546
rect 292404 -3744 293004 -2782
rect 296004 -4106 296604 6000
rect 296004 -4342 296186 -4106
rect 296422 -4342 296604 -4106
rect 296004 -4426 296604 -4342
rect 296004 -4662 296186 -4426
rect 296422 -4662 296604 -4426
rect 296004 -5624 296604 -4662
rect 281604 -7162 281786 -6926
rect 282022 -7162 282204 -6926
rect 281604 -7246 282204 -7162
rect 281604 -7482 281786 -7246
rect 282022 -7482 282204 -7246
rect 281604 -7504 282204 -7482
rect 299604 -5986 300204 6000
rect 306804 5952 306832 6016
rect 306896 5952 306912 6016
rect 306976 5952 306992 6016
rect 307056 5952 307072 6016
rect 307136 5952 307152 6016
rect 307216 5952 307232 6016
rect 307296 5952 307312 6016
rect 307376 5952 307404 6016
rect 306804 4928 307404 5952
rect 306804 4864 306832 4928
rect 306896 4864 306912 4928
rect 306976 4864 306992 4928
rect 307056 4864 307072 4928
rect 307136 4864 307152 4928
rect 307216 4864 307232 4928
rect 307296 4864 307312 4928
rect 307376 4864 307404 4928
rect 306804 3840 307404 4864
rect 306804 3776 306832 3840
rect 306896 3776 306912 3840
rect 306976 3776 306992 3840
rect 307056 3776 307072 3840
rect 307136 3776 307152 3840
rect 307216 3776 307232 3840
rect 307296 3776 307312 3840
rect 307376 3776 307404 3840
rect 306804 2752 307404 3776
rect 306804 2688 306832 2752
rect 306896 2688 306912 2752
rect 306976 2688 306992 2752
rect 307056 2688 307072 2752
rect 307136 2688 307152 2752
rect 307216 2688 307232 2752
rect 307296 2688 307312 2752
rect 307376 2688 307404 2752
rect 306804 -1286 307404 2688
rect 306804 -1522 306986 -1286
rect 307222 -1522 307404 -1286
rect 306804 -1606 307404 -1522
rect 306804 -1842 306986 -1606
rect 307222 -1842 307404 -1606
rect 306804 -1864 307404 -1842
rect 310404 -3166 311004 6000
rect 310404 -3402 310586 -3166
rect 310822 -3402 311004 -3166
rect 310404 -3486 311004 -3402
rect 310404 -3722 310586 -3486
rect 310822 -3722 311004 -3486
rect 310404 -3744 311004 -3722
rect 314004 -5046 314604 6000
rect 314004 -5282 314186 -5046
rect 314422 -5282 314604 -5046
rect 314004 -5366 314604 -5282
rect 314004 -5602 314186 -5366
rect 314422 -5602 314604 -5366
rect 314004 -5624 314604 -5602
rect 299604 -6222 299786 -5986
rect 300022 -6222 300204 -5986
rect 299604 -6306 300204 -6222
rect 299604 -6542 299786 -6306
rect 300022 -6542 300204 -6306
rect 299604 -7504 300204 -6542
rect 317604 -6926 318204 6000
rect 324804 5472 325404 6048
rect 342804 6016 343404 6048
rect 324804 5408 324832 5472
rect 324896 5408 324912 5472
rect 324976 5408 324992 5472
rect 325056 5408 325072 5472
rect 325136 5408 325152 5472
rect 325216 5408 325232 5472
rect 325296 5408 325312 5472
rect 325376 5408 325404 5472
rect 324804 4384 325404 5408
rect 324804 4320 324832 4384
rect 324896 4320 324912 4384
rect 324976 4320 324992 4384
rect 325056 4320 325072 4384
rect 325136 4320 325152 4384
rect 325216 4320 325232 4384
rect 325296 4320 325312 4384
rect 325376 4320 325404 4384
rect 324804 3296 325404 4320
rect 324804 3232 324832 3296
rect 324896 3232 324912 3296
rect 324976 3232 324992 3296
rect 325056 3232 325072 3296
rect 325136 3232 325152 3296
rect 325216 3232 325232 3296
rect 325296 3232 325312 3296
rect 325376 3232 325404 3296
rect 324804 2406 325404 3232
rect 324804 2208 324986 2406
rect 325222 2208 325404 2406
rect 324804 2144 324832 2208
rect 324896 2144 324912 2208
rect 324976 2170 324986 2208
rect 325222 2170 325232 2208
rect 324976 2144 324992 2170
rect 325056 2144 325072 2170
rect 325136 2144 325152 2170
rect 325216 2144 325232 2170
rect 325296 2144 325312 2208
rect 325376 2144 325404 2208
rect 324804 2086 325404 2144
rect 324804 1850 324986 2086
rect 325222 1850 325404 2086
rect 324804 -346 325404 1850
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1864 325404 -902
rect 328404 -2226 329004 6000
rect 328404 -2462 328586 -2226
rect 328822 -2462 329004 -2226
rect 328404 -2546 329004 -2462
rect 328404 -2782 328586 -2546
rect 328822 -2782 329004 -2546
rect 328404 -3744 329004 -2782
rect 332004 -4106 332604 6000
rect 332004 -4342 332186 -4106
rect 332422 -4342 332604 -4106
rect 332004 -4426 332604 -4342
rect 332004 -4662 332186 -4426
rect 332422 -4662 332604 -4426
rect 332004 -5624 332604 -4662
rect 317604 -7162 317786 -6926
rect 318022 -7162 318204 -6926
rect 317604 -7246 318204 -7162
rect 317604 -7482 317786 -7246
rect 318022 -7482 318204 -7246
rect 317604 -7504 318204 -7482
rect 335604 -5986 336204 6000
rect 342804 5952 342832 6016
rect 342896 5952 342912 6016
rect 342976 5952 342992 6016
rect 343056 5952 343072 6016
rect 343136 5952 343152 6016
rect 343216 5952 343232 6016
rect 343296 5952 343312 6016
rect 343376 5952 343404 6016
rect 342804 4928 343404 5952
rect 342804 4864 342832 4928
rect 342896 4864 342912 4928
rect 342976 4864 342992 4928
rect 343056 4864 343072 4928
rect 343136 4864 343152 4928
rect 343216 4864 343232 4928
rect 343296 4864 343312 4928
rect 343376 4864 343404 4928
rect 342804 3840 343404 4864
rect 342804 3776 342832 3840
rect 342896 3776 342912 3840
rect 342976 3776 342992 3840
rect 343056 3776 343072 3840
rect 343136 3776 343152 3840
rect 343216 3776 343232 3840
rect 343296 3776 343312 3840
rect 343376 3776 343404 3840
rect 342804 2752 343404 3776
rect 342804 2688 342832 2752
rect 342896 2688 342912 2752
rect 342976 2688 342992 2752
rect 343056 2688 343072 2752
rect 343136 2688 343152 2752
rect 343216 2688 343232 2752
rect 343296 2688 343312 2752
rect 343376 2688 343404 2752
rect 342804 -1286 343404 2688
rect 342804 -1522 342986 -1286
rect 343222 -1522 343404 -1286
rect 342804 -1606 343404 -1522
rect 342804 -1842 342986 -1606
rect 343222 -1842 343404 -1606
rect 342804 -1864 343404 -1842
rect 346404 -3166 347004 6000
rect 346404 -3402 346586 -3166
rect 346822 -3402 347004 -3166
rect 346404 -3486 347004 -3402
rect 346404 -3722 346586 -3486
rect 346822 -3722 347004 -3486
rect 346404 -3744 347004 -3722
rect 350004 -5046 350604 6000
rect 350004 -5282 350186 -5046
rect 350422 -5282 350604 -5046
rect 350004 -5366 350604 -5282
rect 350004 -5602 350186 -5366
rect 350422 -5602 350604 -5366
rect 350004 -5624 350604 -5602
rect 335604 -6222 335786 -5986
rect 336022 -6222 336204 -5986
rect 335604 -6306 336204 -6222
rect 335604 -6542 335786 -6306
rect 336022 -6542 336204 -6306
rect 335604 -7504 336204 -6542
rect 353604 -6926 354204 6000
rect 360804 5472 361404 6048
rect 378804 6016 379404 6048
rect 360804 5408 360832 5472
rect 360896 5408 360912 5472
rect 360976 5408 360992 5472
rect 361056 5408 361072 5472
rect 361136 5408 361152 5472
rect 361216 5408 361232 5472
rect 361296 5408 361312 5472
rect 361376 5408 361404 5472
rect 360804 4384 361404 5408
rect 360804 4320 360832 4384
rect 360896 4320 360912 4384
rect 360976 4320 360992 4384
rect 361056 4320 361072 4384
rect 361136 4320 361152 4384
rect 361216 4320 361232 4384
rect 361296 4320 361312 4384
rect 361376 4320 361404 4384
rect 360804 3296 361404 4320
rect 360804 3232 360832 3296
rect 360896 3232 360912 3296
rect 360976 3232 360992 3296
rect 361056 3232 361072 3296
rect 361136 3232 361152 3296
rect 361216 3232 361232 3296
rect 361296 3232 361312 3296
rect 361376 3232 361404 3296
rect 360804 2406 361404 3232
rect 360804 2208 360986 2406
rect 361222 2208 361404 2406
rect 360804 2144 360832 2208
rect 360896 2144 360912 2208
rect 360976 2170 360986 2208
rect 361222 2170 361232 2208
rect 360976 2144 360992 2170
rect 361056 2144 361072 2170
rect 361136 2144 361152 2170
rect 361216 2144 361232 2170
rect 361296 2144 361312 2208
rect 361376 2144 361404 2208
rect 360804 2086 361404 2144
rect 360804 1850 360986 2086
rect 361222 1850 361404 2086
rect 360804 -346 361404 1850
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1864 361404 -902
rect 364404 -2226 365004 6000
rect 364404 -2462 364586 -2226
rect 364822 -2462 365004 -2226
rect 364404 -2546 365004 -2462
rect 364404 -2782 364586 -2546
rect 364822 -2782 365004 -2546
rect 364404 -3744 365004 -2782
rect 368004 -4106 368604 6000
rect 368004 -4342 368186 -4106
rect 368422 -4342 368604 -4106
rect 368004 -4426 368604 -4342
rect 368004 -4662 368186 -4426
rect 368422 -4662 368604 -4426
rect 368004 -5624 368604 -4662
rect 353604 -7162 353786 -6926
rect 354022 -7162 354204 -6926
rect 353604 -7246 354204 -7162
rect 353604 -7482 353786 -7246
rect 354022 -7482 354204 -7246
rect 353604 -7504 354204 -7482
rect 371604 -5986 372204 6000
rect 378804 5952 378832 6016
rect 378896 5952 378912 6016
rect 378976 5952 378992 6016
rect 379056 5952 379072 6016
rect 379136 5952 379152 6016
rect 379216 5952 379232 6016
rect 379296 5952 379312 6016
rect 379376 5952 379404 6016
rect 378804 4928 379404 5952
rect 378804 4864 378832 4928
rect 378896 4864 378912 4928
rect 378976 4864 378992 4928
rect 379056 4864 379072 4928
rect 379136 4864 379152 4928
rect 379216 4864 379232 4928
rect 379296 4864 379312 4928
rect 379376 4864 379404 4928
rect 378804 3840 379404 4864
rect 378804 3776 378832 3840
rect 378896 3776 378912 3840
rect 378976 3776 378992 3840
rect 379056 3776 379072 3840
rect 379136 3776 379152 3840
rect 379216 3776 379232 3840
rect 379296 3776 379312 3840
rect 379376 3776 379404 3840
rect 378804 2752 379404 3776
rect 378804 2688 378832 2752
rect 378896 2688 378912 2752
rect 378976 2688 378992 2752
rect 379056 2688 379072 2752
rect 379136 2688 379152 2752
rect 379216 2688 379232 2752
rect 379296 2688 379312 2752
rect 379376 2688 379404 2752
rect 378804 -1286 379404 2688
rect 378804 -1522 378986 -1286
rect 379222 -1522 379404 -1286
rect 378804 -1606 379404 -1522
rect 378804 -1842 378986 -1606
rect 379222 -1842 379404 -1606
rect 378804 -1864 379404 -1842
rect 382404 -3166 383004 6000
rect 382404 -3402 382586 -3166
rect 382822 -3402 383004 -3166
rect 382404 -3486 383004 -3402
rect 382404 -3722 382586 -3486
rect 382822 -3722 383004 -3486
rect 382404 -3744 383004 -3722
rect 386004 -5046 386604 6000
rect 386004 -5282 386186 -5046
rect 386422 -5282 386604 -5046
rect 386004 -5366 386604 -5282
rect 386004 -5602 386186 -5366
rect 386422 -5602 386604 -5366
rect 386004 -5624 386604 -5602
rect 371604 -6222 371786 -5986
rect 372022 -6222 372204 -5986
rect 371604 -6306 372204 -6222
rect 371604 -6542 371786 -6306
rect 372022 -6542 372204 -6306
rect 371604 -7504 372204 -6542
rect 389604 -6926 390204 6000
rect 396804 5472 397404 6048
rect 414804 6016 415404 6048
rect 396804 5408 396832 5472
rect 396896 5408 396912 5472
rect 396976 5408 396992 5472
rect 397056 5408 397072 5472
rect 397136 5408 397152 5472
rect 397216 5408 397232 5472
rect 397296 5408 397312 5472
rect 397376 5408 397404 5472
rect 396804 4384 397404 5408
rect 396804 4320 396832 4384
rect 396896 4320 396912 4384
rect 396976 4320 396992 4384
rect 397056 4320 397072 4384
rect 397136 4320 397152 4384
rect 397216 4320 397232 4384
rect 397296 4320 397312 4384
rect 397376 4320 397404 4384
rect 396804 3296 397404 4320
rect 396804 3232 396832 3296
rect 396896 3232 396912 3296
rect 396976 3232 396992 3296
rect 397056 3232 397072 3296
rect 397136 3232 397152 3296
rect 397216 3232 397232 3296
rect 397296 3232 397312 3296
rect 397376 3232 397404 3296
rect 396804 2406 397404 3232
rect 396804 2208 396986 2406
rect 397222 2208 397404 2406
rect 396804 2144 396832 2208
rect 396896 2144 396912 2208
rect 396976 2170 396986 2208
rect 397222 2170 397232 2208
rect 396976 2144 396992 2170
rect 397056 2144 397072 2170
rect 397136 2144 397152 2170
rect 397216 2144 397232 2170
rect 397296 2144 397312 2208
rect 397376 2144 397404 2208
rect 396804 2086 397404 2144
rect 396804 1850 396986 2086
rect 397222 1850 397404 2086
rect 396804 -346 397404 1850
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1864 397404 -902
rect 400404 -2226 401004 6000
rect 400404 -2462 400586 -2226
rect 400822 -2462 401004 -2226
rect 400404 -2546 401004 -2462
rect 400404 -2782 400586 -2546
rect 400822 -2782 401004 -2546
rect 400404 -3744 401004 -2782
rect 404004 -4106 404604 6000
rect 404004 -4342 404186 -4106
rect 404422 -4342 404604 -4106
rect 404004 -4426 404604 -4342
rect 404004 -4662 404186 -4426
rect 404422 -4662 404604 -4426
rect 404004 -5624 404604 -4662
rect 389604 -7162 389786 -6926
rect 390022 -7162 390204 -6926
rect 389604 -7246 390204 -7162
rect 389604 -7482 389786 -7246
rect 390022 -7482 390204 -7246
rect 389604 -7504 390204 -7482
rect 407604 -5986 408204 6000
rect 414804 5952 414832 6016
rect 414896 5952 414912 6016
rect 414976 5952 414992 6016
rect 415056 5952 415072 6016
rect 415136 5952 415152 6016
rect 415216 5952 415232 6016
rect 415296 5952 415312 6016
rect 415376 5952 415404 6016
rect 414804 4928 415404 5952
rect 414804 4864 414832 4928
rect 414896 4864 414912 4928
rect 414976 4864 414992 4928
rect 415056 4864 415072 4928
rect 415136 4864 415152 4928
rect 415216 4864 415232 4928
rect 415296 4864 415312 4928
rect 415376 4864 415404 4928
rect 414804 3840 415404 4864
rect 414804 3776 414832 3840
rect 414896 3776 414912 3840
rect 414976 3776 414992 3840
rect 415056 3776 415072 3840
rect 415136 3776 415152 3840
rect 415216 3776 415232 3840
rect 415296 3776 415312 3840
rect 415376 3776 415404 3840
rect 414804 2752 415404 3776
rect 414804 2688 414832 2752
rect 414896 2688 414912 2752
rect 414976 2688 414992 2752
rect 415056 2688 415072 2752
rect 415136 2688 415152 2752
rect 415216 2688 415232 2752
rect 415296 2688 415312 2752
rect 415376 2688 415404 2752
rect 414804 -1286 415404 2688
rect 414804 -1522 414986 -1286
rect 415222 -1522 415404 -1286
rect 414804 -1606 415404 -1522
rect 414804 -1842 414986 -1606
rect 415222 -1842 415404 -1606
rect 414804 -1864 415404 -1842
rect 418404 -3166 419004 6000
rect 418404 -3402 418586 -3166
rect 418822 -3402 419004 -3166
rect 418404 -3486 419004 -3402
rect 418404 -3722 418586 -3486
rect 418822 -3722 419004 -3486
rect 418404 -3744 419004 -3722
rect 422004 -5046 422604 6000
rect 422004 -5282 422186 -5046
rect 422422 -5282 422604 -5046
rect 422004 -5366 422604 -5282
rect 422004 -5602 422186 -5366
rect 422422 -5602 422604 -5366
rect 422004 -5624 422604 -5602
rect 407604 -6222 407786 -5986
rect 408022 -6222 408204 -5986
rect 407604 -6306 408204 -6222
rect 407604 -6542 407786 -6306
rect 408022 -6542 408204 -6306
rect 407604 -7504 408204 -6542
rect 425604 -6926 426204 6000
rect 432804 5472 433404 6048
rect 450804 6016 451404 6048
rect 432804 5408 432832 5472
rect 432896 5408 432912 5472
rect 432976 5408 432992 5472
rect 433056 5408 433072 5472
rect 433136 5408 433152 5472
rect 433216 5408 433232 5472
rect 433296 5408 433312 5472
rect 433376 5408 433404 5472
rect 432804 4384 433404 5408
rect 432804 4320 432832 4384
rect 432896 4320 432912 4384
rect 432976 4320 432992 4384
rect 433056 4320 433072 4384
rect 433136 4320 433152 4384
rect 433216 4320 433232 4384
rect 433296 4320 433312 4384
rect 433376 4320 433404 4384
rect 432804 3296 433404 4320
rect 432804 3232 432832 3296
rect 432896 3232 432912 3296
rect 432976 3232 432992 3296
rect 433056 3232 433072 3296
rect 433136 3232 433152 3296
rect 433216 3232 433232 3296
rect 433296 3232 433312 3296
rect 433376 3232 433404 3296
rect 432804 2406 433404 3232
rect 432804 2208 432986 2406
rect 433222 2208 433404 2406
rect 432804 2144 432832 2208
rect 432896 2144 432912 2208
rect 432976 2170 432986 2208
rect 433222 2170 433232 2208
rect 432976 2144 432992 2170
rect 433056 2144 433072 2170
rect 433136 2144 433152 2170
rect 433216 2144 433232 2170
rect 433296 2144 433312 2208
rect 433376 2144 433404 2208
rect 432804 2086 433404 2144
rect 432804 1850 432986 2086
rect 433222 1850 433404 2086
rect 432804 -346 433404 1850
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1864 433404 -902
rect 436404 -2226 437004 6000
rect 436404 -2462 436586 -2226
rect 436822 -2462 437004 -2226
rect 436404 -2546 437004 -2462
rect 436404 -2782 436586 -2546
rect 436822 -2782 437004 -2546
rect 436404 -3744 437004 -2782
rect 440004 -4106 440604 6000
rect 440004 -4342 440186 -4106
rect 440422 -4342 440604 -4106
rect 440004 -4426 440604 -4342
rect 440004 -4662 440186 -4426
rect 440422 -4662 440604 -4426
rect 440004 -5624 440604 -4662
rect 425604 -7162 425786 -6926
rect 426022 -7162 426204 -6926
rect 425604 -7246 426204 -7162
rect 425604 -7482 425786 -7246
rect 426022 -7482 426204 -7246
rect 425604 -7504 426204 -7482
rect 443604 -5986 444204 6000
rect 450804 5952 450832 6016
rect 450896 5952 450912 6016
rect 450976 5952 450992 6016
rect 451056 5952 451072 6016
rect 451136 5952 451152 6016
rect 451216 5952 451232 6016
rect 451296 5952 451312 6016
rect 451376 5952 451404 6016
rect 450804 4928 451404 5952
rect 450804 4864 450832 4928
rect 450896 4864 450912 4928
rect 450976 4864 450992 4928
rect 451056 4864 451072 4928
rect 451136 4864 451152 4928
rect 451216 4864 451232 4928
rect 451296 4864 451312 4928
rect 451376 4864 451404 4928
rect 450804 3840 451404 4864
rect 450804 3776 450832 3840
rect 450896 3776 450912 3840
rect 450976 3776 450992 3840
rect 451056 3776 451072 3840
rect 451136 3776 451152 3840
rect 451216 3776 451232 3840
rect 451296 3776 451312 3840
rect 451376 3776 451404 3840
rect 450804 2752 451404 3776
rect 450804 2688 450832 2752
rect 450896 2688 450912 2752
rect 450976 2688 450992 2752
rect 451056 2688 451072 2752
rect 451136 2688 451152 2752
rect 451216 2688 451232 2752
rect 451296 2688 451312 2752
rect 451376 2688 451404 2752
rect 450804 -1286 451404 2688
rect 450804 -1522 450986 -1286
rect 451222 -1522 451404 -1286
rect 450804 -1606 451404 -1522
rect 450804 -1842 450986 -1606
rect 451222 -1842 451404 -1606
rect 450804 -1864 451404 -1842
rect 454404 -3166 455004 6000
rect 454404 -3402 454586 -3166
rect 454822 -3402 455004 -3166
rect 454404 -3486 455004 -3402
rect 454404 -3722 454586 -3486
rect 454822 -3722 455004 -3486
rect 454404 -3744 455004 -3722
rect 458004 -5046 458604 6000
rect 458004 -5282 458186 -5046
rect 458422 -5282 458604 -5046
rect 458004 -5366 458604 -5282
rect 458004 -5602 458186 -5366
rect 458422 -5602 458604 -5366
rect 458004 -5624 458604 -5602
rect 443604 -6222 443786 -5986
rect 444022 -6222 444204 -5986
rect 443604 -6306 444204 -6222
rect 443604 -6542 443786 -6306
rect 444022 -6542 444204 -6306
rect 443604 -7504 444204 -6542
rect 461604 -6926 462204 6000
rect 468804 5472 469404 6048
rect 486804 6016 487404 6048
rect 468804 5408 468832 5472
rect 468896 5408 468912 5472
rect 468976 5408 468992 5472
rect 469056 5408 469072 5472
rect 469136 5408 469152 5472
rect 469216 5408 469232 5472
rect 469296 5408 469312 5472
rect 469376 5408 469404 5472
rect 468804 4384 469404 5408
rect 468804 4320 468832 4384
rect 468896 4320 468912 4384
rect 468976 4320 468992 4384
rect 469056 4320 469072 4384
rect 469136 4320 469152 4384
rect 469216 4320 469232 4384
rect 469296 4320 469312 4384
rect 469376 4320 469404 4384
rect 468804 3296 469404 4320
rect 468804 3232 468832 3296
rect 468896 3232 468912 3296
rect 468976 3232 468992 3296
rect 469056 3232 469072 3296
rect 469136 3232 469152 3296
rect 469216 3232 469232 3296
rect 469296 3232 469312 3296
rect 469376 3232 469404 3296
rect 468804 2406 469404 3232
rect 468804 2208 468986 2406
rect 469222 2208 469404 2406
rect 468804 2144 468832 2208
rect 468896 2144 468912 2208
rect 468976 2170 468986 2208
rect 469222 2170 469232 2208
rect 468976 2144 468992 2170
rect 469056 2144 469072 2170
rect 469136 2144 469152 2170
rect 469216 2144 469232 2170
rect 469296 2144 469312 2208
rect 469376 2144 469404 2208
rect 468804 2086 469404 2144
rect 468804 1850 468986 2086
rect 469222 1850 469404 2086
rect 468804 -346 469404 1850
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1864 469404 -902
rect 472404 -2226 473004 6000
rect 472404 -2462 472586 -2226
rect 472822 -2462 473004 -2226
rect 472404 -2546 473004 -2462
rect 472404 -2782 472586 -2546
rect 472822 -2782 473004 -2546
rect 472404 -3744 473004 -2782
rect 476004 -4106 476604 6000
rect 476004 -4342 476186 -4106
rect 476422 -4342 476604 -4106
rect 476004 -4426 476604 -4342
rect 476004 -4662 476186 -4426
rect 476422 -4662 476604 -4426
rect 476004 -5624 476604 -4662
rect 461604 -7162 461786 -6926
rect 462022 -7162 462204 -6926
rect 461604 -7246 462204 -7162
rect 461604 -7482 461786 -7246
rect 462022 -7482 462204 -7246
rect 461604 -7504 462204 -7482
rect 479604 -5986 480204 6000
rect 486804 5952 486832 6016
rect 486896 5952 486912 6016
rect 486976 5952 486992 6016
rect 487056 5952 487072 6016
rect 487136 5952 487152 6016
rect 487216 5952 487232 6016
rect 487296 5952 487312 6016
rect 487376 5952 487404 6016
rect 486804 4928 487404 5952
rect 486804 4864 486832 4928
rect 486896 4864 486912 4928
rect 486976 4864 486992 4928
rect 487056 4864 487072 4928
rect 487136 4864 487152 4928
rect 487216 4864 487232 4928
rect 487296 4864 487312 4928
rect 487376 4864 487404 4928
rect 486804 3840 487404 4864
rect 486804 3776 486832 3840
rect 486896 3776 486912 3840
rect 486976 3776 486992 3840
rect 487056 3776 487072 3840
rect 487136 3776 487152 3840
rect 487216 3776 487232 3840
rect 487296 3776 487312 3840
rect 487376 3776 487404 3840
rect 486804 2752 487404 3776
rect 486804 2688 486832 2752
rect 486896 2688 486912 2752
rect 486976 2688 486992 2752
rect 487056 2688 487072 2752
rect 487136 2688 487152 2752
rect 487216 2688 487232 2752
rect 487296 2688 487312 2752
rect 487376 2688 487404 2752
rect 486804 -1286 487404 2688
rect 486804 -1522 486986 -1286
rect 487222 -1522 487404 -1286
rect 486804 -1606 487404 -1522
rect 486804 -1842 486986 -1606
rect 487222 -1842 487404 -1606
rect 486804 -1864 487404 -1842
rect 490404 -3166 491004 6000
rect 490404 -3402 490586 -3166
rect 490822 -3402 491004 -3166
rect 490404 -3486 491004 -3402
rect 490404 -3722 490586 -3486
rect 490822 -3722 491004 -3486
rect 490404 -3744 491004 -3722
rect 494004 -5046 494604 6000
rect 494004 -5282 494186 -5046
rect 494422 -5282 494604 -5046
rect 494004 -5366 494604 -5282
rect 494004 -5602 494186 -5366
rect 494422 -5602 494604 -5366
rect 494004 -5624 494604 -5602
rect 479604 -6222 479786 -5986
rect 480022 -6222 480204 -5986
rect 479604 -6306 480204 -6222
rect 479604 -6542 479786 -6306
rect 480022 -6542 480204 -6306
rect 479604 -7504 480204 -6542
rect 497604 -6926 498204 6000
rect 504804 5472 505404 6048
rect 522804 6016 523404 6048
rect 504804 5408 504832 5472
rect 504896 5408 504912 5472
rect 504976 5408 504992 5472
rect 505056 5408 505072 5472
rect 505136 5408 505152 5472
rect 505216 5408 505232 5472
rect 505296 5408 505312 5472
rect 505376 5408 505404 5472
rect 504804 4384 505404 5408
rect 504804 4320 504832 4384
rect 504896 4320 504912 4384
rect 504976 4320 504992 4384
rect 505056 4320 505072 4384
rect 505136 4320 505152 4384
rect 505216 4320 505232 4384
rect 505296 4320 505312 4384
rect 505376 4320 505404 4384
rect 504804 3296 505404 4320
rect 504804 3232 504832 3296
rect 504896 3232 504912 3296
rect 504976 3232 504992 3296
rect 505056 3232 505072 3296
rect 505136 3232 505152 3296
rect 505216 3232 505232 3296
rect 505296 3232 505312 3296
rect 505376 3232 505404 3296
rect 504804 2406 505404 3232
rect 504804 2208 504986 2406
rect 505222 2208 505404 2406
rect 504804 2144 504832 2208
rect 504896 2144 504912 2208
rect 504976 2170 504986 2208
rect 505222 2170 505232 2208
rect 504976 2144 504992 2170
rect 505056 2144 505072 2170
rect 505136 2144 505152 2170
rect 505216 2144 505232 2170
rect 505296 2144 505312 2208
rect 505376 2144 505404 2208
rect 504804 2086 505404 2144
rect 504804 1850 504986 2086
rect 505222 1850 505404 2086
rect 504804 -346 505404 1850
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1864 505404 -902
rect 508404 -2226 509004 6000
rect 508404 -2462 508586 -2226
rect 508822 -2462 509004 -2226
rect 508404 -2546 509004 -2462
rect 508404 -2782 508586 -2546
rect 508822 -2782 509004 -2546
rect 508404 -3744 509004 -2782
rect 512004 -4106 512604 6000
rect 512004 -4342 512186 -4106
rect 512422 -4342 512604 -4106
rect 512004 -4426 512604 -4342
rect 512004 -4662 512186 -4426
rect 512422 -4662 512604 -4426
rect 512004 -5624 512604 -4662
rect 497604 -7162 497786 -6926
rect 498022 -7162 498204 -6926
rect 497604 -7246 498204 -7162
rect 497604 -7482 497786 -7246
rect 498022 -7482 498204 -7246
rect 497604 -7504 498204 -7482
rect 515604 -5986 516204 6000
rect 522804 5952 522832 6016
rect 522896 5952 522912 6016
rect 522976 5952 522992 6016
rect 523056 5952 523072 6016
rect 523136 5952 523152 6016
rect 523216 5952 523232 6016
rect 523296 5952 523312 6016
rect 523376 5952 523404 6016
rect 522804 4928 523404 5952
rect 522804 4864 522832 4928
rect 522896 4864 522912 4928
rect 522976 4864 522992 4928
rect 523056 4864 523072 4928
rect 523136 4864 523152 4928
rect 523216 4864 523232 4928
rect 523296 4864 523312 4928
rect 523376 4864 523404 4928
rect 522804 3840 523404 4864
rect 522804 3776 522832 3840
rect 522896 3776 522912 3840
rect 522976 3776 522992 3840
rect 523056 3776 523072 3840
rect 523136 3776 523152 3840
rect 523216 3776 523232 3840
rect 523296 3776 523312 3840
rect 523376 3776 523404 3840
rect 522804 2752 523404 3776
rect 522804 2688 522832 2752
rect 522896 2688 522912 2752
rect 522976 2688 522992 2752
rect 523056 2688 523072 2752
rect 523136 2688 523152 2752
rect 523216 2688 523232 2752
rect 523296 2688 523312 2752
rect 523376 2688 523404 2752
rect 522804 -1286 523404 2688
rect 522804 -1522 522986 -1286
rect 523222 -1522 523404 -1286
rect 522804 -1606 523404 -1522
rect 522804 -1842 522986 -1606
rect 523222 -1842 523404 -1606
rect 522804 -1864 523404 -1842
rect 526404 -3166 527004 6000
rect 526404 -3402 526586 -3166
rect 526822 -3402 527004 -3166
rect 526404 -3486 527004 -3402
rect 526404 -3722 526586 -3486
rect 526822 -3722 527004 -3486
rect 526404 -3744 527004 -3722
rect 530004 -5046 530604 6000
rect 530004 -5282 530186 -5046
rect 530422 -5282 530604 -5046
rect 530004 -5366 530604 -5282
rect 530004 -5602 530186 -5366
rect 530422 -5602 530604 -5366
rect 530004 -5624 530604 -5602
rect 515604 -6222 515786 -5986
rect 516022 -6222 516204 -5986
rect 515604 -6306 516204 -6222
rect 515604 -6542 515786 -6306
rect 516022 -6542 516204 -6306
rect 515604 -7504 516204 -6542
rect 533604 -6926 534204 6000
rect 540804 5472 541404 6048
rect 558804 6016 559404 6048
rect 540804 5408 540832 5472
rect 540896 5408 540912 5472
rect 540976 5408 540992 5472
rect 541056 5408 541072 5472
rect 541136 5408 541152 5472
rect 541216 5408 541232 5472
rect 541296 5408 541312 5472
rect 541376 5408 541404 5472
rect 540804 4384 541404 5408
rect 540804 4320 540832 4384
rect 540896 4320 540912 4384
rect 540976 4320 540992 4384
rect 541056 4320 541072 4384
rect 541136 4320 541152 4384
rect 541216 4320 541232 4384
rect 541296 4320 541312 4384
rect 541376 4320 541404 4384
rect 540804 3296 541404 4320
rect 540804 3232 540832 3296
rect 540896 3232 540912 3296
rect 540976 3232 540992 3296
rect 541056 3232 541072 3296
rect 541136 3232 541152 3296
rect 541216 3232 541232 3296
rect 541296 3232 541312 3296
rect 541376 3232 541404 3296
rect 540804 2406 541404 3232
rect 540804 2208 540986 2406
rect 541222 2208 541404 2406
rect 540804 2144 540832 2208
rect 540896 2144 540912 2208
rect 540976 2170 540986 2208
rect 541222 2170 541232 2208
rect 540976 2144 540992 2170
rect 541056 2144 541072 2170
rect 541136 2144 541152 2170
rect 541216 2144 541232 2170
rect 541296 2144 541312 2208
rect 541376 2144 541404 2208
rect 540804 2086 541404 2144
rect 540804 1850 540986 2086
rect 541222 1850 541404 2086
rect 540804 -346 541404 1850
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1864 541404 -902
rect 544404 -2226 545004 6000
rect 544404 -2462 544586 -2226
rect 544822 -2462 545004 -2226
rect 544404 -2546 545004 -2462
rect 544404 -2782 544586 -2546
rect 544822 -2782 545004 -2546
rect 544404 -3744 545004 -2782
rect 548004 -4106 548604 6000
rect 548004 -4342 548186 -4106
rect 548422 -4342 548604 -4106
rect 548004 -4426 548604 -4342
rect 548004 -4662 548186 -4426
rect 548422 -4662 548604 -4426
rect 548004 -5624 548604 -4662
rect 533604 -7162 533786 -6926
rect 534022 -7162 534204 -6926
rect 533604 -7246 534204 -7162
rect 533604 -7482 533786 -7246
rect 534022 -7482 534204 -7246
rect 533604 -7504 534204 -7482
rect 551604 -5986 552204 6000
rect 558804 5952 558832 6016
rect 558896 5952 558912 6016
rect 558976 5952 558992 6016
rect 559056 5952 559072 6016
rect 559136 5952 559152 6016
rect 559216 5952 559232 6016
rect 559296 5952 559312 6016
rect 559376 5952 559404 6016
rect 558804 4928 559404 5952
rect 558804 4864 558832 4928
rect 558896 4864 558912 4928
rect 558976 4864 558992 4928
rect 559056 4864 559072 4928
rect 559136 4864 559152 4928
rect 559216 4864 559232 4928
rect 559296 4864 559312 4928
rect 559376 4864 559404 4928
rect 558804 3840 559404 4864
rect 558804 3776 558832 3840
rect 558896 3776 558912 3840
rect 558976 3776 558992 3840
rect 559056 3776 559072 3840
rect 559136 3776 559152 3840
rect 559216 3776 559232 3840
rect 559296 3776 559312 3840
rect 559376 3776 559404 3840
rect 558804 2752 559404 3776
rect 558804 2688 558832 2752
rect 558896 2688 558912 2752
rect 558976 2688 558992 2752
rect 559056 2688 559072 2752
rect 559136 2688 559152 2752
rect 559216 2688 559232 2752
rect 559296 2688 559312 2752
rect 559376 2688 559404 2752
rect 558804 -1286 559404 2688
rect 558804 -1522 558986 -1286
rect 559222 -1522 559404 -1286
rect 558804 -1606 559404 -1522
rect 558804 -1842 558986 -1606
rect 559222 -1842 559404 -1606
rect 558804 -1864 559404 -1842
rect 562404 -3166 563004 6000
rect 562404 -3402 562586 -3166
rect 562822 -3402 563004 -3166
rect 562404 -3486 563004 -3402
rect 562404 -3722 562586 -3486
rect 562822 -3722 563004 -3486
rect 562404 -3744 563004 -3722
rect 566004 -5046 566604 6000
rect 566004 -5282 566186 -5046
rect 566422 -5282 566604 -5046
rect 566004 -5366 566604 -5282
rect 566004 -5602 566186 -5366
rect 566422 -5602 566604 -5366
rect 566004 -5624 566604 -5602
rect 551604 -6222 551786 -5986
rect 552022 -6222 552204 -5986
rect 551604 -6306 552204 -6222
rect 551604 -6542 551786 -6306
rect 552022 -6542 552204 -6306
rect 551604 -7504 552204 -6542
rect 569604 -6926 570204 6000
rect 576804 5472 577404 6048
rect 576804 5408 576832 5472
rect 576896 5408 576912 5472
rect 576976 5408 576992 5472
rect 577056 5408 577072 5472
rect 577136 5408 577152 5472
rect 577216 5408 577232 5472
rect 577296 5408 577312 5472
rect 577376 5408 577404 5472
rect 576804 4384 577404 5408
rect 576804 4320 576832 4384
rect 576896 4320 576912 4384
rect 576976 4320 576992 4384
rect 577056 4320 577072 4384
rect 577136 4320 577152 4384
rect 577216 4320 577232 4384
rect 577296 4320 577312 4384
rect 577376 4320 577404 4384
rect 576804 3296 577404 4320
rect 576804 3232 576832 3296
rect 576896 3232 576912 3296
rect 576976 3232 576992 3296
rect 577056 3232 577072 3296
rect 577136 3232 577152 3296
rect 577216 3232 577232 3296
rect 577296 3232 577312 3296
rect 577376 3232 577404 3296
rect 576804 2406 577404 3232
rect 576804 2208 576986 2406
rect 577222 2208 577404 2406
rect 576804 2144 576832 2208
rect 576896 2144 576912 2208
rect 576976 2170 576986 2208
rect 577222 2170 577232 2208
rect 576976 2144 576992 2170
rect 577056 2144 577072 2170
rect 577136 2144 577152 2170
rect 577216 2144 577232 2170
rect 577296 2144 577312 2208
rect 577376 2144 577404 2208
rect 576804 2086 577404 2144
rect 576804 1850 576986 2086
rect 577222 1850 577404 2086
rect 576804 -346 577404 1850
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1864 577404 -902
rect 580404 5818 580586 6054
rect 580822 5818 581004 6054
rect 580404 5734 581004 5818
rect 580404 5498 580586 5734
rect 580822 5498 581004 5734
rect 580404 -2226 581004 5498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686406 585920 704282
rect 585320 686170 585502 686406
rect 585738 686170 585920 686406
rect 585320 686086 585920 686170
rect 585320 685850 585502 686086
rect 585738 685850 585920 686086
rect 585320 650406 585920 685850
rect 585320 650170 585502 650406
rect 585738 650170 585920 650406
rect 585320 650086 585920 650170
rect 585320 649850 585502 650086
rect 585738 649850 585920 650086
rect 585320 614406 585920 649850
rect 585320 614170 585502 614406
rect 585738 614170 585920 614406
rect 585320 614086 585920 614170
rect 585320 613850 585502 614086
rect 585738 613850 585920 614086
rect 585320 578406 585920 613850
rect 585320 578170 585502 578406
rect 585738 578170 585920 578406
rect 585320 578086 585920 578170
rect 585320 577850 585502 578086
rect 585738 577850 585920 578086
rect 585320 542406 585920 577850
rect 585320 542170 585502 542406
rect 585738 542170 585920 542406
rect 585320 542086 585920 542170
rect 585320 541850 585502 542086
rect 585738 541850 585920 542086
rect 585320 506406 585920 541850
rect 585320 506170 585502 506406
rect 585738 506170 585920 506406
rect 585320 506086 585920 506170
rect 585320 505850 585502 506086
rect 585738 505850 585920 506086
rect 585320 470406 585920 505850
rect 585320 470170 585502 470406
rect 585738 470170 585920 470406
rect 585320 470086 585920 470170
rect 585320 469850 585502 470086
rect 585738 469850 585920 470086
rect 585320 434406 585920 469850
rect 585320 434170 585502 434406
rect 585738 434170 585920 434406
rect 585320 434086 585920 434170
rect 585320 433850 585502 434086
rect 585738 433850 585920 434086
rect 585320 398406 585920 433850
rect 585320 398170 585502 398406
rect 585738 398170 585920 398406
rect 585320 398086 585920 398170
rect 585320 397850 585502 398086
rect 585738 397850 585920 398086
rect 585320 362406 585920 397850
rect 585320 362170 585502 362406
rect 585738 362170 585920 362406
rect 585320 362086 585920 362170
rect 585320 361850 585502 362086
rect 585738 361850 585920 362086
rect 585320 326406 585920 361850
rect 585320 326170 585502 326406
rect 585738 326170 585920 326406
rect 585320 326086 585920 326170
rect 585320 325850 585502 326086
rect 585738 325850 585920 326086
rect 585320 290406 585920 325850
rect 585320 290170 585502 290406
rect 585738 290170 585920 290406
rect 585320 290086 585920 290170
rect 585320 289850 585502 290086
rect 585738 289850 585920 290086
rect 585320 254406 585920 289850
rect 585320 254170 585502 254406
rect 585738 254170 585920 254406
rect 585320 254086 585920 254170
rect 585320 253850 585502 254086
rect 585738 253850 585920 254086
rect 585320 218406 585920 253850
rect 585320 218170 585502 218406
rect 585738 218170 585920 218406
rect 585320 218086 585920 218170
rect 585320 217850 585502 218086
rect 585738 217850 585920 218086
rect 585320 182406 585920 217850
rect 585320 182170 585502 182406
rect 585738 182170 585920 182406
rect 585320 182086 585920 182170
rect 585320 181850 585502 182086
rect 585738 181850 585920 182086
rect 585320 146406 585920 181850
rect 585320 146170 585502 146406
rect 585738 146170 585920 146406
rect 585320 146086 585920 146170
rect 585320 145850 585502 146086
rect 585738 145850 585920 146086
rect 585320 110406 585920 145850
rect 585320 110170 585502 110406
rect 585738 110170 585920 110406
rect 585320 110086 585920 110170
rect 585320 109850 585502 110086
rect 585738 109850 585920 110086
rect 585320 74406 585920 109850
rect 585320 74170 585502 74406
rect 585738 74170 585920 74406
rect 585320 74086 585920 74170
rect 585320 73850 585502 74086
rect 585738 73850 585920 74086
rect 585320 38406 585920 73850
rect 585320 38170 585502 38406
rect 585738 38170 585920 38406
rect 585320 38086 585920 38170
rect 585320 37850 585502 38086
rect 585738 37850 585920 38086
rect 585320 2406 585920 37850
rect 585320 2170 585502 2406
rect 585738 2170 585920 2406
rect 585320 2086 585920 2170
rect 585320 1850 585502 2086
rect 585738 1850 585920 2086
rect 585320 -346 585920 1850
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586260 668406 586860 705222
rect 586260 668170 586442 668406
rect 586678 668170 586860 668406
rect 586260 668086 586860 668170
rect 586260 667850 586442 668086
rect 586678 667850 586860 668086
rect 586260 632406 586860 667850
rect 586260 632170 586442 632406
rect 586678 632170 586860 632406
rect 586260 632086 586860 632170
rect 586260 631850 586442 632086
rect 586678 631850 586860 632086
rect 586260 596406 586860 631850
rect 586260 596170 586442 596406
rect 586678 596170 586860 596406
rect 586260 596086 586860 596170
rect 586260 595850 586442 596086
rect 586678 595850 586860 596086
rect 586260 560406 586860 595850
rect 586260 560170 586442 560406
rect 586678 560170 586860 560406
rect 586260 560086 586860 560170
rect 586260 559850 586442 560086
rect 586678 559850 586860 560086
rect 586260 524406 586860 559850
rect 586260 524170 586442 524406
rect 586678 524170 586860 524406
rect 586260 524086 586860 524170
rect 586260 523850 586442 524086
rect 586678 523850 586860 524086
rect 586260 488406 586860 523850
rect 586260 488170 586442 488406
rect 586678 488170 586860 488406
rect 586260 488086 586860 488170
rect 586260 487850 586442 488086
rect 586678 487850 586860 488086
rect 586260 452406 586860 487850
rect 586260 452170 586442 452406
rect 586678 452170 586860 452406
rect 586260 452086 586860 452170
rect 586260 451850 586442 452086
rect 586678 451850 586860 452086
rect 586260 416406 586860 451850
rect 586260 416170 586442 416406
rect 586678 416170 586860 416406
rect 586260 416086 586860 416170
rect 586260 415850 586442 416086
rect 586678 415850 586860 416086
rect 586260 380406 586860 415850
rect 586260 380170 586442 380406
rect 586678 380170 586860 380406
rect 586260 380086 586860 380170
rect 586260 379850 586442 380086
rect 586678 379850 586860 380086
rect 586260 344406 586860 379850
rect 586260 344170 586442 344406
rect 586678 344170 586860 344406
rect 586260 344086 586860 344170
rect 586260 343850 586442 344086
rect 586678 343850 586860 344086
rect 586260 308406 586860 343850
rect 586260 308170 586442 308406
rect 586678 308170 586860 308406
rect 586260 308086 586860 308170
rect 586260 307850 586442 308086
rect 586678 307850 586860 308086
rect 586260 272406 586860 307850
rect 586260 272170 586442 272406
rect 586678 272170 586860 272406
rect 586260 272086 586860 272170
rect 586260 271850 586442 272086
rect 586678 271850 586860 272086
rect 586260 236406 586860 271850
rect 586260 236170 586442 236406
rect 586678 236170 586860 236406
rect 586260 236086 586860 236170
rect 586260 235850 586442 236086
rect 586678 235850 586860 236086
rect 586260 200406 586860 235850
rect 586260 200170 586442 200406
rect 586678 200170 586860 200406
rect 586260 200086 586860 200170
rect 586260 199850 586442 200086
rect 586678 199850 586860 200086
rect 586260 164406 586860 199850
rect 586260 164170 586442 164406
rect 586678 164170 586860 164406
rect 586260 164086 586860 164170
rect 586260 163850 586442 164086
rect 586678 163850 586860 164086
rect 586260 128406 586860 163850
rect 586260 128170 586442 128406
rect 586678 128170 586860 128406
rect 586260 128086 586860 128170
rect 586260 127850 586442 128086
rect 586678 127850 586860 128086
rect 586260 92406 586860 127850
rect 586260 92170 586442 92406
rect 586678 92170 586860 92406
rect 586260 92086 586860 92170
rect 586260 91850 586442 92086
rect 586678 91850 586860 92086
rect 586260 56406 586860 91850
rect 586260 56170 586442 56406
rect 586678 56170 586860 56406
rect 586260 56086 586860 56170
rect 586260 55850 586442 56086
rect 586678 55850 586860 56086
rect 586260 20406 586860 55850
rect 586260 20170 586442 20406
rect 586678 20170 586860 20406
rect 586260 20086 586860 20170
rect 586260 19850 586442 20086
rect 586678 19850 586860 20086
rect 586260 -1286 586860 19850
rect 586260 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect 586260 -1606 586860 -1522
rect 586260 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect 586260 -1864 586860 -1842
rect 587200 690054 587800 706162
rect 587200 689818 587382 690054
rect 587618 689818 587800 690054
rect 587200 689734 587800 689818
rect 587200 689498 587382 689734
rect 587618 689498 587800 689734
rect 587200 654054 587800 689498
rect 587200 653818 587382 654054
rect 587618 653818 587800 654054
rect 587200 653734 587800 653818
rect 587200 653498 587382 653734
rect 587618 653498 587800 653734
rect 587200 618054 587800 653498
rect 587200 617818 587382 618054
rect 587618 617818 587800 618054
rect 587200 617734 587800 617818
rect 587200 617498 587382 617734
rect 587618 617498 587800 617734
rect 587200 582054 587800 617498
rect 587200 581818 587382 582054
rect 587618 581818 587800 582054
rect 587200 581734 587800 581818
rect 587200 581498 587382 581734
rect 587618 581498 587800 581734
rect 587200 546054 587800 581498
rect 587200 545818 587382 546054
rect 587618 545818 587800 546054
rect 587200 545734 587800 545818
rect 587200 545498 587382 545734
rect 587618 545498 587800 545734
rect 587200 510054 587800 545498
rect 587200 509818 587382 510054
rect 587618 509818 587800 510054
rect 587200 509734 587800 509818
rect 587200 509498 587382 509734
rect 587618 509498 587800 509734
rect 587200 474054 587800 509498
rect 587200 473818 587382 474054
rect 587618 473818 587800 474054
rect 587200 473734 587800 473818
rect 587200 473498 587382 473734
rect 587618 473498 587800 473734
rect 587200 438054 587800 473498
rect 587200 437818 587382 438054
rect 587618 437818 587800 438054
rect 587200 437734 587800 437818
rect 587200 437498 587382 437734
rect 587618 437498 587800 437734
rect 587200 402054 587800 437498
rect 587200 401818 587382 402054
rect 587618 401818 587800 402054
rect 587200 401734 587800 401818
rect 587200 401498 587382 401734
rect 587618 401498 587800 401734
rect 587200 366054 587800 401498
rect 587200 365818 587382 366054
rect 587618 365818 587800 366054
rect 587200 365734 587800 365818
rect 587200 365498 587382 365734
rect 587618 365498 587800 365734
rect 587200 330054 587800 365498
rect 587200 329818 587382 330054
rect 587618 329818 587800 330054
rect 587200 329734 587800 329818
rect 587200 329498 587382 329734
rect 587618 329498 587800 329734
rect 587200 294054 587800 329498
rect 587200 293818 587382 294054
rect 587618 293818 587800 294054
rect 587200 293734 587800 293818
rect 587200 293498 587382 293734
rect 587618 293498 587800 293734
rect 587200 258054 587800 293498
rect 587200 257818 587382 258054
rect 587618 257818 587800 258054
rect 587200 257734 587800 257818
rect 587200 257498 587382 257734
rect 587618 257498 587800 257734
rect 587200 222054 587800 257498
rect 587200 221818 587382 222054
rect 587618 221818 587800 222054
rect 587200 221734 587800 221818
rect 587200 221498 587382 221734
rect 587618 221498 587800 221734
rect 587200 186054 587800 221498
rect 587200 185818 587382 186054
rect 587618 185818 587800 186054
rect 587200 185734 587800 185818
rect 587200 185498 587382 185734
rect 587618 185498 587800 185734
rect 587200 150054 587800 185498
rect 587200 149818 587382 150054
rect 587618 149818 587800 150054
rect 587200 149734 587800 149818
rect 587200 149498 587382 149734
rect 587618 149498 587800 149734
rect 587200 114054 587800 149498
rect 587200 113818 587382 114054
rect 587618 113818 587800 114054
rect 587200 113734 587800 113818
rect 587200 113498 587382 113734
rect 587618 113498 587800 113734
rect 587200 78054 587800 113498
rect 587200 77818 587382 78054
rect 587618 77818 587800 78054
rect 587200 77734 587800 77818
rect 587200 77498 587382 77734
rect 587618 77498 587800 77734
rect 587200 42054 587800 77498
rect 587200 41818 587382 42054
rect 587618 41818 587800 42054
rect 587200 41734 587800 41818
rect 587200 41498 587382 41734
rect 587618 41498 587800 41734
rect 587200 6054 587800 41498
rect 587200 5818 587382 6054
rect 587618 5818 587800 6054
rect 587200 5734 587800 5818
rect 587200 5498 587382 5734
rect 587618 5498 587800 5734
rect 580404 -2462 580586 -2226
rect 580822 -2462 581004 -2226
rect 580404 -2546 581004 -2462
rect 580404 -2782 580586 -2546
rect 580822 -2782 581004 -2546
rect 580404 -3744 581004 -2782
rect 587200 -2226 587800 5498
rect 587200 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect 587200 -2546 587800 -2462
rect 587200 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect 587200 -2804 587800 -2782
rect 588140 672054 588740 707102
rect 588140 671818 588322 672054
rect 588558 671818 588740 672054
rect 588140 671734 588740 671818
rect 588140 671498 588322 671734
rect 588558 671498 588740 671734
rect 588140 636054 588740 671498
rect 588140 635818 588322 636054
rect 588558 635818 588740 636054
rect 588140 635734 588740 635818
rect 588140 635498 588322 635734
rect 588558 635498 588740 635734
rect 588140 600054 588740 635498
rect 588140 599818 588322 600054
rect 588558 599818 588740 600054
rect 588140 599734 588740 599818
rect 588140 599498 588322 599734
rect 588558 599498 588740 599734
rect 588140 564054 588740 599498
rect 588140 563818 588322 564054
rect 588558 563818 588740 564054
rect 588140 563734 588740 563818
rect 588140 563498 588322 563734
rect 588558 563498 588740 563734
rect 588140 528054 588740 563498
rect 588140 527818 588322 528054
rect 588558 527818 588740 528054
rect 588140 527734 588740 527818
rect 588140 527498 588322 527734
rect 588558 527498 588740 527734
rect 588140 492054 588740 527498
rect 588140 491818 588322 492054
rect 588558 491818 588740 492054
rect 588140 491734 588740 491818
rect 588140 491498 588322 491734
rect 588558 491498 588740 491734
rect 588140 456054 588740 491498
rect 588140 455818 588322 456054
rect 588558 455818 588740 456054
rect 588140 455734 588740 455818
rect 588140 455498 588322 455734
rect 588558 455498 588740 455734
rect 588140 420054 588740 455498
rect 588140 419818 588322 420054
rect 588558 419818 588740 420054
rect 588140 419734 588740 419818
rect 588140 419498 588322 419734
rect 588558 419498 588740 419734
rect 588140 384054 588740 419498
rect 588140 383818 588322 384054
rect 588558 383818 588740 384054
rect 588140 383734 588740 383818
rect 588140 383498 588322 383734
rect 588558 383498 588740 383734
rect 588140 348054 588740 383498
rect 588140 347818 588322 348054
rect 588558 347818 588740 348054
rect 588140 347734 588740 347818
rect 588140 347498 588322 347734
rect 588558 347498 588740 347734
rect 588140 312054 588740 347498
rect 588140 311818 588322 312054
rect 588558 311818 588740 312054
rect 588140 311734 588740 311818
rect 588140 311498 588322 311734
rect 588558 311498 588740 311734
rect 588140 276054 588740 311498
rect 588140 275818 588322 276054
rect 588558 275818 588740 276054
rect 588140 275734 588740 275818
rect 588140 275498 588322 275734
rect 588558 275498 588740 275734
rect 588140 240054 588740 275498
rect 588140 239818 588322 240054
rect 588558 239818 588740 240054
rect 588140 239734 588740 239818
rect 588140 239498 588322 239734
rect 588558 239498 588740 239734
rect 588140 204054 588740 239498
rect 588140 203818 588322 204054
rect 588558 203818 588740 204054
rect 588140 203734 588740 203818
rect 588140 203498 588322 203734
rect 588558 203498 588740 203734
rect 588140 168054 588740 203498
rect 588140 167818 588322 168054
rect 588558 167818 588740 168054
rect 588140 167734 588740 167818
rect 588140 167498 588322 167734
rect 588558 167498 588740 167734
rect 588140 132054 588740 167498
rect 588140 131818 588322 132054
rect 588558 131818 588740 132054
rect 588140 131734 588740 131818
rect 588140 131498 588322 131734
rect 588558 131498 588740 131734
rect 588140 96054 588740 131498
rect 588140 95818 588322 96054
rect 588558 95818 588740 96054
rect 588140 95734 588740 95818
rect 588140 95498 588322 95734
rect 588558 95498 588740 95734
rect 588140 60054 588740 95498
rect 588140 59818 588322 60054
rect 588558 59818 588740 60054
rect 588140 59734 588740 59818
rect 588140 59498 588322 59734
rect 588558 59498 588740 59734
rect 588140 24054 588740 59498
rect 588140 23818 588322 24054
rect 588558 23818 588740 24054
rect 588140 23734 588740 23818
rect 588140 23498 588322 23734
rect 588558 23498 588740 23734
rect 588140 -3166 588740 23498
rect 588140 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect 588140 -3486 588740 -3402
rect 588140 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect 588140 -3744 588740 -3722
rect 589080 693654 589680 708042
rect 589080 693418 589262 693654
rect 589498 693418 589680 693654
rect 589080 693334 589680 693418
rect 589080 693098 589262 693334
rect 589498 693098 589680 693334
rect 589080 657654 589680 693098
rect 589080 657418 589262 657654
rect 589498 657418 589680 657654
rect 589080 657334 589680 657418
rect 589080 657098 589262 657334
rect 589498 657098 589680 657334
rect 589080 621654 589680 657098
rect 589080 621418 589262 621654
rect 589498 621418 589680 621654
rect 589080 621334 589680 621418
rect 589080 621098 589262 621334
rect 589498 621098 589680 621334
rect 589080 585654 589680 621098
rect 589080 585418 589262 585654
rect 589498 585418 589680 585654
rect 589080 585334 589680 585418
rect 589080 585098 589262 585334
rect 589498 585098 589680 585334
rect 589080 549654 589680 585098
rect 589080 549418 589262 549654
rect 589498 549418 589680 549654
rect 589080 549334 589680 549418
rect 589080 549098 589262 549334
rect 589498 549098 589680 549334
rect 589080 513654 589680 549098
rect 589080 513418 589262 513654
rect 589498 513418 589680 513654
rect 589080 513334 589680 513418
rect 589080 513098 589262 513334
rect 589498 513098 589680 513334
rect 589080 477654 589680 513098
rect 589080 477418 589262 477654
rect 589498 477418 589680 477654
rect 589080 477334 589680 477418
rect 589080 477098 589262 477334
rect 589498 477098 589680 477334
rect 589080 441654 589680 477098
rect 589080 441418 589262 441654
rect 589498 441418 589680 441654
rect 589080 441334 589680 441418
rect 589080 441098 589262 441334
rect 589498 441098 589680 441334
rect 589080 405654 589680 441098
rect 589080 405418 589262 405654
rect 589498 405418 589680 405654
rect 589080 405334 589680 405418
rect 589080 405098 589262 405334
rect 589498 405098 589680 405334
rect 589080 369654 589680 405098
rect 589080 369418 589262 369654
rect 589498 369418 589680 369654
rect 589080 369334 589680 369418
rect 589080 369098 589262 369334
rect 589498 369098 589680 369334
rect 589080 333654 589680 369098
rect 589080 333418 589262 333654
rect 589498 333418 589680 333654
rect 589080 333334 589680 333418
rect 589080 333098 589262 333334
rect 589498 333098 589680 333334
rect 589080 297654 589680 333098
rect 589080 297418 589262 297654
rect 589498 297418 589680 297654
rect 589080 297334 589680 297418
rect 589080 297098 589262 297334
rect 589498 297098 589680 297334
rect 589080 261654 589680 297098
rect 589080 261418 589262 261654
rect 589498 261418 589680 261654
rect 589080 261334 589680 261418
rect 589080 261098 589262 261334
rect 589498 261098 589680 261334
rect 589080 225654 589680 261098
rect 589080 225418 589262 225654
rect 589498 225418 589680 225654
rect 589080 225334 589680 225418
rect 589080 225098 589262 225334
rect 589498 225098 589680 225334
rect 589080 189654 589680 225098
rect 589080 189418 589262 189654
rect 589498 189418 589680 189654
rect 589080 189334 589680 189418
rect 589080 189098 589262 189334
rect 589498 189098 589680 189334
rect 589080 153654 589680 189098
rect 589080 153418 589262 153654
rect 589498 153418 589680 153654
rect 589080 153334 589680 153418
rect 589080 153098 589262 153334
rect 589498 153098 589680 153334
rect 589080 117654 589680 153098
rect 589080 117418 589262 117654
rect 589498 117418 589680 117654
rect 589080 117334 589680 117418
rect 589080 117098 589262 117334
rect 589498 117098 589680 117334
rect 589080 81654 589680 117098
rect 589080 81418 589262 81654
rect 589498 81418 589680 81654
rect 589080 81334 589680 81418
rect 589080 81098 589262 81334
rect 589498 81098 589680 81334
rect 589080 45654 589680 81098
rect 589080 45418 589262 45654
rect 589498 45418 589680 45654
rect 589080 45334 589680 45418
rect 589080 45098 589262 45334
rect 589498 45098 589680 45334
rect 589080 9654 589680 45098
rect 589080 9418 589262 9654
rect 589498 9418 589680 9654
rect 589080 9334 589680 9418
rect 589080 9098 589262 9334
rect 589498 9098 589680 9334
rect 589080 -4106 589680 9098
rect 589080 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect 589080 -4426 589680 -4342
rect 589080 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect 589080 -4684 589680 -4662
rect 590020 675654 590620 708982
rect 590020 675418 590202 675654
rect 590438 675418 590620 675654
rect 590020 675334 590620 675418
rect 590020 675098 590202 675334
rect 590438 675098 590620 675334
rect 590020 639654 590620 675098
rect 590020 639418 590202 639654
rect 590438 639418 590620 639654
rect 590020 639334 590620 639418
rect 590020 639098 590202 639334
rect 590438 639098 590620 639334
rect 590020 603654 590620 639098
rect 590020 603418 590202 603654
rect 590438 603418 590620 603654
rect 590020 603334 590620 603418
rect 590020 603098 590202 603334
rect 590438 603098 590620 603334
rect 590020 567654 590620 603098
rect 590020 567418 590202 567654
rect 590438 567418 590620 567654
rect 590020 567334 590620 567418
rect 590020 567098 590202 567334
rect 590438 567098 590620 567334
rect 590020 531654 590620 567098
rect 590020 531418 590202 531654
rect 590438 531418 590620 531654
rect 590020 531334 590620 531418
rect 590020 531098 590202 531334
rect 590438 531098 590620 531334
rect 590020 495654 590620 531098
rect 590020 495418 590202 495654
rect 590438 495418 590620 495654
rect 590020 495334 590620 495418
rect 590020 495098 590202 495334
rect 590438 495098 590620 495334
rect 590020 459654 590620 495098
rect 590020 459418 590202 459654
rect 590438 459418 590620 459654
rect 590020 459334 590620 459418
rect 590020 459098 590202 459334
rect 590438 459098 590620 459334
rect 590020 423654 590620 459098
rect 590020 423418 590202 423654
rect 590438 423418 590620 423654
rect 590020 423334 590620 423418
rect 590020 423098 590202 423334
rect 590438 423098 590620 423334
rect 590020 387654 590620 423098
rect 590020 387418 590202 387654
rect 590438 387418 590620 387654
rect 590020 387334 590620 387418
rect 590020 387098 590202 387334
rect 590438 387098 590620 387334
rect 590020 351654 590620 387098
rect 590020 351418 590202 351654
rect 590438 351418 590620 351654
rect 590020 351334 590620 351418
rect 590020 351098 590202 351334
rect 590438 351098 590620 351334
rect 590020 315654 590620 351098
rect 590020 315418 590202 315654
rect 590438 315418 590620 315654
rect 590020 315334 590620 315418
rect 590020 315098 590202 315334
rect 590438 315098 590620 315334
rect 590020 279654 590620 315098
rect 590020 279418 590202 279654
rect 590438 279418 590620 279654
rect 590020 279334 590620 279418
rect 590020 279098 590202 279334
rect 590438 279098 590620 279334
rect 590020 243654 590620 279098
rect 590020 243418 590202 243654
rect 590438 243418 590620 243654
rect 590020 243334 590620 243418
rect 590020 243098 590202 243334
rect 590438 243098 590620 243334
rect 590020 207654 590620 243098
rect 590020 207418 590202 207654
rect 590438 207418 590620 207654
rect 590020 207334 590620 207418
rect 590020 207098 590202 207334
rect 590438 207098 590620 207334
rect 590020 171654 590620 207098
rect 590020 171418 590202 171654
rect 590438 171418 590620 171654
rect 590020 171334 590620 171418
rect 590020 171098 590202 171334
rect 590438 171098 590620 171334
rect 590020 135654 590620 171098
rect 590020 135418 590202 135654
rect 590438 135418 590620 135654
rect 590020 135334 590620 135418
rect 590020 135098 590202 135334
rect 590438 135098 590620 135334
rect 590020 99654 590620 135098
rect 590020 99418 590202 99654
rect 590438 99418 590620 99654
rect 590020 99334 590620 99418
rect 590020 99098 590202 99334
rect 590438 99098 590620 99334
rect 590020 63654 590620 99098
rect 590020 63418 590202 63654
rect 590438 63418 590620 63654
rect 590020 63334 590620 63418
rect 590020 63098 590202 63334
rect 590438 63098 590620 63334
rect 590020 27654 590620 63098
rect 590020 27418 590202 27654
rect 590438 27418 590620 27654
rect 590020 27334 590620 27418
rect 590020 27098 590202 27334
rect 590438 27098 590620 27334
rect 590020 -5046 590620 27098
rect 590020 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect 590020 -5366 590620 -5282
rect 590020 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect 590020 -5624 590620 -5602
rect 590960 697254 591560 709922
rect 590960 697018 591142 697254
rect 591378 697018 591560 697254
rect 590960 696934 591560 697018
rect 590960 696698 591142 696934
rect 591378 696698 591560 696934
rect 590960 661254 591560 696698
rect 590960 661018 591142 661254
rect 591378 661018 591560 661254
rect 590960 660934 591560 661018
rect 590960 660698 591142 660934
rect 591378 660698 591560 660934
rect 590960 625254 591560 660698
rect 590960 625018 591142 625254
rect 591378 625018 591560 625254
rect 590960 624934 591560 625018
rect 590960 624698 591142 624934
rect 591378 624698 591560 624934
rect 590960 589254 591560 624698
rect 590960 589018 591142 589254
rect 591378 589018 591560 589254
rect 590960 588934 591560 589018
rect 590960 588698 591142 588934
rect 591378 588698 591560 588934
rect 590960 553254 591560 588698
rect 590960 553018 591142 553254
rect 591378 553018 591560 553254
rect 590960 552934 591560 553018
rect 590960 552698 591142 552934
rect 591378 552698 591560 552934
rect 590960 517254 591560 552698
rect 590960 517018 591142 517254
rect 591378 517018 591560 517254
rect 590960 516934 591560 517018
rect 590960 516698 591142 516934
rect 591378 516698 591560 516934
rect 590960 481254 591560 516698
rect 590960 481018 591142 481254
rect 591378 481018 591560 481254
rect 590960 480934 591560 481018
rect 590960 480698 591142 480934
rect 591378 480698 591560 480934
rect 590960 445254 591560 480698
rect 590960 445018 591142 445254
rect 591378 445018 591560 445254
rect 590960 444934 591560 445018
rect 590960 444698 591142 444934
rect 591378 444698 591560 444934
rect 590960 409254 591560 444698
rect 590960 409018 591142 409254
rect 591378 409018 591560 409254
rect 590960 408934 591560 409018
rect 590960 408698 591142 408934
rect 591378 408698 591560 408934
rect 590960 373254 591560 408698
rect 590960 373018 591142 373254
rect 591378 373018 591560 373254
rect 590960 372934 591560 373018
rect 590960 372698 591142 372934
rect 591378 372698 591560 372934
rect 590960 337254 591560 372698
rect 590960 337018 591142 337254
rect 591378 337018 591560 337254
rect 590960 336934 591560 337018
rect 590960 336698 591142 336934
rect 591378 336698 591560 336934
rect 590960 301254 591560 336698
rect 590960 301018 591142 301254
rect 591378 301018 591560 301254
rect 590960 300934 591560 301018
rect 590960 300698 591142 300934
rect 591378 300698 591560 300934
rect 590960 265254 591560 300698
rect 590960 265018 591142 265254
rect 591378 265018 591560 265254
rect 590960 264934 591560 265018
rect 590960 264698 591142 264934
rect 591378 264698 591560 264934
rect 590960 229254 591560 264698
rect 590960 229018 591142 229254
rect 591378 229018 591560 229254
rect 590960 228934 591560 229018
rect 590960 228698 591142 228934
rect 591378 228698 591560 228934
rect 590960 193254 591560 228698
rect 590960 193018 591142 193254
rect 591378 193018 591560 193254
rect 590960 192934 591560 193018
rect 590960 192698 591142 192934
rect 591378 192698 591560 192934
rect 590960 157254 591560 192698
rect 590960 157018 591142 157254
rect 591378 157018 591560 157254
rect 590960 156934 591560 157018
rect 590960 156698 591142 156934
rect 591378 156698 591560 156934
rect 590960 121254 591560 156698
rect 590960 121018 591142 121254
rect 591378 121018 591560 121254
rect 590960 120934 591560 121018
rect 590960 120698 591142 120934
rect 591378 120698 591560 120934
rect 590960 85254 591560 120698
rect 590960 85018 591142 85254
rect 591378 85018 591560 85254
rect 590960 84934 591560 85018
rect 590960 84698 591142 84934
rect 591378 84698 591560 84934
rect 590960 49254 591560 84698
rect 590960 49018 591142 49254
rect 591378 49018 591560 49254
rect 590960 48934 591560 49018
rect 590960 48698 591142 48934
rect 591378 48698 591560 48934
rect 590960 13254 591560 48698
rect 590960 13018 591142 13254
rect 591378 13018 591560 13254
rect 590960 12934 591560 13018
rect 590960 12698 591142 12934
rect 591378 12698 591560 12934
rect 590960 -5986 591560 12698
rect 590960 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect 590960 -6306 591560 -6222
rect 590960 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect 590960 -6564 591560 -6542
rect 591900 679254 592500 710862
rect 591900 679018 592082 679254
rect 592318 679018 592500 679254
rect 591900 678934 592500 679018
rect 591900 678698 592082 678934
rect 592318 678698 592500 678934
rect 591900 643254 592500 678698
rect 591900 643018 592082 643254
rect 592318 643018 592500 643254
rect 591900 642934 592500 643018
rect 591900 642698 592082 642934
rect 592318 642698 592500 642934
rect 591900 607254 592500 642698
rect 591900 607018 592082 607254
rect 592318 607018 592500 607254
rect 591900 606934 592500 607018
rect 591900 606698 592082 606934
rect 592318 606698 592500 606934
rect 591900 571254 592500 606698
rect 591900 571018 592082 571254
rect 592318 571018 592500 571254
rect 591900 570934 592500 571018
rect 591900 570698 592082 570934
rect 592318 570698 592500 570934
rect 591900 535254 592500 570698
rect 591900 535018 592082 535254
rect 592318 535018 592500 535254
rect 591900 534934 592500 535018
rect 591900 534698 592082 534934
rect 592318 534698 592500 534934
rect 591900 499254 592500 534698
rect 591900 499018 592082 499254
rect 592318 499018 592500 499254
rect 591900 498934 592500 499018
rect 591900 498698 592082 498934
rect 592318 498698 592500 498934
rect 591900 463254 592500 498698
rect 591900 463018 592082 463254
rect 592318 463018 592500 463254
rect 591900 462934 592500 463018
rect 591900 462698 592082 462934
rect 592318 462698 592500 462934
rect 591900 427254 592500 462698
rect 591900 427018 592082 427254
rect 592318 427018 592500 427254
rect 591900 426934 592500 427018
rect 591900 426698 592082 426934
rect 592318 426698 592500 426934
rect 591900 391254 592500 426698
rect 591900 391018 592082 391254
rect 592318 391018 592500 391254
rect 591900 390934 592500 391018
rect 591900 390698 592082 390934
rect 592318 390698 592500 390934
rect 591900 355254 592500 390698
rect 591900 355018 592082 355254
rect 592318 355018 592500 355254
rect 591900 354934 592500 355018
rect 591900 354698 592082 354934
rect 592318 354698 592500 354934
rect 591900 319254 592500 354698
rect 591900 319018 592082 319254
rect 592318 319018 592500 319254
rect 591900 318934 592500 319018
rect 591900 318698 592082 318934
rect 592318 318698 592500 318934
rect 591900 283254 592500 318698
rect 591900 283018 592082 283254
rect 592318 283018 592500 283254
rect 591900 282934 592500 283018
rect 591900 282698 592082 282934
rect 592318 282698 592500 282934
rect 591900 247254 592500 282698
rect 591900 247018 592082 247254
rect 592318 247018 592500 247254
rect 591900 246934 592500 247018
rect 591900 246698 592082 246934
rect 592318 246698 592500 246934
rect 591900 211254 592500 246698
rect 591900 211018 592082 211254
rect 592318 211018 592500 211254
rect 591900 210934 592500 211018
rect 591900 210698 592082 210934
rect 592318 210698 592500 210934
rect 591900 175254 592500 210698
rect 591900 175018 592082 175254
rect 592318 175018 592500 175254
rect 591900 174934 592500 175018
rect 591900 174698 592082 174934
rect 592318 174698 592500 174934
rect 591900 139254 592500 174698
rect 591900 139018 592082 139254
rect 592318 139018 592500 139254
rect 591900 138934 592500 139018
rect 591900 138698 592082 138934
rect 592318 138698 592500 138934
rect 591900 103254 592500 138698
rect 591900 103018 592082 103254
rect 592318 103018 592500 103254
rect 591900 102934 592500 103018
rect 591900 102698 592082 102934
rect 592318 102698 592500 102934
rect 591900 67254 592500 102698
rect 591900 67018 592082 67254
rect 592318 67018 592500 67254
rect 591900 66934 592500 67018
rect 591900 66698 592082 66934
rect 592318 66698 592500 66934
rect 591900 31254 592500 66698
rect 591900 31018 592082 31254
rect 592318 31018 592500 31254
rect 591900 30934 592500 31018
rect 591900 30698 592082 30934
rect 592318 30698 592500 30934
rect 569604 -7162 569786 -6926
rect 570022 -7162 570204 -6926
rect 569604 -7246 570204 -7162
rect 569604 -7482 569786 -7246
rect 570022 -7482 570204 -7246
rect 569604 -7504 570204 -7482
rect 591900 -6926 592500 30698
rect 591900 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect 591900 -7246 592500 -7162
rect 591900 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect 591900 -7504 592500 -7482
<< via4 >>
rect -8394 711182 -8158 711418
rect -8394 710862 -8158 711098
rect -8394 679018 -8158 679254
rect -8394 678698 -8158 678934
rect -8394 643018 -8158 643254
rect -8394 642698 -8158 642934
rect -8394 607018 -8158 607254
rect -8394 606698 -8158 606934
rect -8394 571018 -8158 571254
rect -8394 570698 -8158 570934
rect -8394 535018 -8158 535254
rect -8394 534698 -8158 534934
rect -8394 499018 -8158 499254
rect -8394 498698 -8158 498934
rect -8394 463018 -8158 463254
rect -8394 462698 -8158 462934
rect -8394 427018 -8158 427254
rect -8394 426698 -8158 426934
rect -8394 391018 -8158 391254
rect -8394 390698 -8158 390934
rect -8394 355018 -8158 355254
rect -8394 354698 -8158 354934
rect -8394 319018 -8158 319254
rect -8394 318698 -8158 318934
rect -8394 283018 -8158 283254
rect -8394 282698 -8158 282934
rect -8394 247018 -8158 247254
rect -8394 246698 -8158 246934
rect -8394 211018 -8158 211254
rect -8394 210698 -8158 210934
rect -8394 175018 -8158 175254
rect -8394 174698 -8158 174934
rect -8394 139018 -8158 139254
rect -8394 138698 -8158 138934
rect -8394 103018 -8158 103254
rect -8394 102698 -8158 102934
rect -8394 67018 -8158 67254
rect -8394 66698 -8158 66934
rect -8394 31018 -8158 31254
rect -8394 30698 -8158 30934
rect -7454 710242 -7218 710478
rect -7454 709922 -7218 710158
rect 11786 710242 12022 710478
rect 11786 709922 12022 710158
rect -7454 697018 -7218 697254
rect -7454 696698 -7218 696934
rect -7454 661018 -7218 661254
rect -7454 660698 -7218 660934
rect -7454 625018 -7218 625254
rect -7454 624698 -7218 624934
rect -7454 589018 -7218 589254
rect -7454 588698 -7218 588934
rect -7454 553018 -7218 553254
rect -7454 552698 -7218 552934
rect -7454 517018 -7218 517254
rect -7454 516698 -7218 516934
rect -7454 481018 -7218 481254
rect -7454 480698 -7218 480934
rect -7454 445018 -7218 445254
rect -7454 444698 -7218 444934
rect -7454 409018 -7218 409254
rect -7454 408698 -7218 408934
rect -7454 373018 -7218 373254
rect -7454 372698 -7218 372934
rect -7454 337018 -7218 337254
rect -7454 336698 -7218 336934
rect -7454 301018 -7218 301254
rect -7454 300698 -7218 300934
rect -7454 265018 -7218 265254
rect -7454 264698 -7218 264934
rect -7454 229018 -7218 229254
rect -7454 228698 -7218 228934
rect -7454 193018 -7218 193254
rect -7454 192698 -7218 192934
rect -7454 157018 -7218 157254
rect -7454 156698 -7218 156934
rect -7454 121018 -7218 121254
rect -7454 120698 -7218 120934
rect -7454 85018 -7218 85254
rect -7454 84698 -7218 84934
rect -7454 49018 -7218 49254
rect -7454 48698 -7218 48934
rect -7454 13018 -7218 13254
rect -7454 12698 -7218 12934
rect -6514 709302 -6278 709538
rect -6514 708982 -6278 709218
rect -6514 675418 -6278 675654
rect -6514 675098 -6278 675334
rect -6514 639418 -6278 639654
rect -6514 639098 -6278 639334
rect -6514 603418 -6278 603654
rect -6514 603098 -6278 603334
rect -6514 567418 -6278 567654
rect -6514 567098 -6278 567334
rect -6514 531418 -6278 531654
rect -6514 531098 -6278 531334
rect -6514 495418 -6278 495654
rect -6514 495098 -6278 495334
rect -6514 459418 -6278 459654
rect -6514 459098 -6278 459334
rect -6514 423418 -6278 423654
rect -6514 423098 -6278 423334
rect -6514 387418 -6278 387654
rect -6514 387098 -6278 387334
rect -6514 351418 -6278 351654
rect -6514 351098 -6278 351334
rect -6514 315418 -6278 315654
rect -6514 315098 -6278 315334
rect -6514 279418 -6278 279654
rect -6514 279098 -6278 279334
rect -6514 243418 -6278 243654
rect -6514 243098 -6278 243334
rect -6514 207418 -6278 207654
rect -6514 207098 -6278 207334
rect -6514 171418 -6278 171654
rect -6514 171098 -6278 171334
rect -6514 135418 -6278 135654
rect -6514 135098 -6278 135334
rect -6514 99418 -6278 99654
rect -6514 99098 -6278 99334
rect -6514 63418 -6278 63654
rect -6514 63098 -6278 63334
rect -6514 27418 -6278 27654
rect -6514 27098 -6278 27334
rect -5574 708362 -5338 708598
rect -5574 708042 -5338 708278
rect 8186 708362 8422 708598
rect 8186 708042 8422 708278
rect -5574 693418 -5338 693654
rect -5574 693098 -5338 693334
rect -5574 657418 -5338 657654
rect -5574 657098 -5338 657334
rect -5574 621418 -5338 621654
rect -5574 621098 -5338 621334
rect -5574 585418 -5338 585654
rect -5574 585098 -5338 585334
rect -5574 549418 -5338 549654
rect -5574 549098 -5338 549334
rect -5574 513418 -5338 513654
rect -5574 513098 -5338 513334
rect -5574 477418 -5338 477654
rect -5574 477098 -5338 477334
rect -5574 441418 -5338 441654
rect -5574 441098 -5338 441334
rect -5574 405418 -5338 405654
rect -5574 405098 -5338 405334
rect -5574 369418 -5338 369654
rect -5574 369098 -5338 369334
rect -5574 333418 -5338 333654
rect -5574 333098 -5338 333334
rect -5574 297418 -5338 297654
rect -5574 297098 -5338 297334
rect -5574 261418 -5338 261654
rect -5574 261098 -5338 261334
rect -5574 225418 -5338 225654
rect -5574 225098 -5338 225334
rect -5574 189418 -5338 189654
rect -5574 189098 -5338 189334
rect -5574 153418 -5338 153654
rect -5574 153098 -5338 153334
rect -5574 117418 -5338 117654
rect -5574 117098 -5338 117334
rect -5574 81418 -5338 81654
rect -5574 81098 -5338 81334
rect -5574 45418 -5338 45654
rect -5574 45098 -5338 45334
rect -5574 9418 -5338 9654
rect -5574 9098 -5338 9334
rect -4634 707422 -4398 707658
rect -4634 707102 -4398 707338
rect -4634 671818 -4398 672054
rect -4634 671498 -4398 671734
rect -4634 635818 -4398 636054
rect -4634 635498 -4398 635734
rect -4634 599818 -4398 600054
rect -4634 599498 -4398 599734
rect -4634 563818 -4398 564054
rect -4634 563498 -4398 563734
rect -4634 527818 -4398 528054
rect -4634 527498 -4398 527734
rect -4634 491818 -4398 492054
rect -4634 491498 -4398 491734
rect -4634 455818 -4398 456054
rect -4634 455498 -4398 455734
rect -4634 419818 -4398 420054
rect -4634 419498 -4398 419734
rect -4634 383818 -4398 384054
rect -4634 383498 -4398 383734
rect -4634 347818 -4398 348054
rect -4634 347498 -4398 347734
rect -4634 311818 -4398 312054
rect -4634 311498 -4398 311734
rect -4634 275818 -4398 276054
rect -4634 275498 -4398 275734
rect -4634 239818 -4398 240054
rect -4634 239498 -4398 239734
rect -4634 203818 -4398 204054
rect -4634 203498 -4398 203734
rect -4634 167818 -4398 168054
rect -4634 167498 -4398 167734
rect -4634 131818 -4398 132054
rect -4634 131498 -4398 131734
rect -4634 95818 -4398 96054
rect -4634 95498 -4398 95734
rect -4634 59818 -4398 60054
rect -4634 59498 -4398 59734
rect -4634 23818 -4398 24054
rect -4634 23498 -4398 23734
rect -3694 706482 -3458 706718
rect -3694 706162 -3458 706398
rect 4586 706482 4822 706718
rect 4586 706162 4822 706398
rect -3694 689818 -3458 690054
rect -3694 689498 -3458 689734
rect -3694 653818 -3458 654054
rect -3694 653498 -3458 653734
rect -3694 617818 -3458 618054
rect -3694 617498 -3458 617734
rect -3694 581818 -3458 582054
rect -3694 581498 -3458 581734
rect -3694 545818 -3458 546054
rect -3694 545498 -3458 545734
rect -3694 509818 -3458 510054
rect -3694 509498 -3458 509734
rect -3694 473818 -3458 474054
rect -3694 473498 -3458 473734
rect -3694 437818 -3458 438054
rect -3694 437498 -3458 437734
rect -3694 401818 -3458 402054
rect -3694 401498 -3458 401734
rect -3694 365818 -3458 366054
rect -3694 365498 -3458 365734
rect -3694 329818 -3458 330054
rect -3694 329498 -3458 329734
rect -3694 293818 -3458 294054
rect -3694 293498 -3458 293734
rect -3694 257818 -3458 258054
rect -3694 257498 -3458 257734
rect -3694 221818 -3458 222054
rect -3694 221498 -3458 221734
rect -3694 185818 -3458 186054
rect -3694 185498 -3458 185734
rect -3694 149818 -3458 150054
rect -3694 149498 -3458 149734
rect -3694 113818 -3458 114054
rect -3694 113498 -3458 113734
rect -3694 77818 -3458 78054
rect -3694 77498 -3458 77734
rect -3694 41818 -3458 42054
rect -3694 41498 -3458 41734
rect -3694 5818 -3458 6054
rect -3694 5498 -3458 5734
rect -2754 705542 -2518 705778
rect -2754 705222 -2518 705458
rect -2754 668170 -2518 668406
rect -2754 667850 -2518 668086
rect -2754 632170 -2518 632406
rect -2754 631850 -2518 632086
rect -2754 596170 -2518 596406
rect -2754 595850 -2518 596086
rect -2754 560170 -2518 560406
rect -2754 559850 -2518 560086
rect -2754 524170 -2518 524406
rect -2754 523850 -2518 524086
rect -2754 488170 -2518 488406
rect -2754 487850 -2518 488086
rect -2754 452170 -2518 452406
rect -2754 451850 -2518 452086
rect -2754 416170 -2518 416406
rect -2754 415850 -2518 416086
rect -2754 380170 -2518 380406
rect -2754 379850 -2518 380086
rect -2754 344170 -2518 344406
rect -2754 343850 -2518 344086
rect -2754 308170 -2518 308406
rect -2754 307850 -2518 308086
rect -2754 272170 -2518 272406
rect -2754 271850 -2518 272086
rect -2754 236170 -2518 236406
rect -2754 235850 -2518 236086
rect -2754 200170 -2518 200406
rect -2754 199850 -2518 200086
rect -2754 164170 -2518 164406
rect -2754 163850 -2518 164086
rect -2754 128170 -2518 128406
rect -2754 127850 -2518 128086
rect -2754 92170 -2518 92406
rect -2754 91850 -2518 92086
rect -2754 56170 -2518 56406
rect -2754 55850 -2518 56086
rect -2754 20170 -2518 20406
rect -2754 19850 -2518 20086
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686170 -1578 686406
rect -1814 685850 -1578 686086
rect -1814 650170 -1578 650406
rect -1814 649850 -1578 650086
rect -1814 614170 -1578 614406
rect -1814 613850 -1578 614086
rect -1814 578170 -1578 578406
rect -1814 577850 -1578 578086
rect -1814 542170 -1578 542406
rect -1814 541850 -1578 542086
rect -1814 506170 -1578 506406
rect -1814 505850 -1578 506086
rect -1814 470170 -1578 470406
rect -1814 469850 -1578 470086
rect -1814 434170 -1578 434406
rect -1814 433850 -1578 434086
rect -1814 398170 -1578 398406
rect -1814 397850 -1578 398086
rect -1814 362170 -1578 362406
rect -1814 361850 -1578 362086
rect -1814 326170 -1578 326406
rect -1814 325850 -1578 326086
rect -1814 290170 -1578 290406
rect -1814 289850 -1578 290086
rect -1814 254170 -1578 254406
rect -1814 253850 -1578 254086
rect -1814 218170 -1578 218406
rect -1814 217850 -1578 218086
rect -1814 182170 -1578 182406
rect -1814 181850 -1578 182086
rect -1814 146170 -1578 146406
rect -1814 145850 -1578 146086
rect -1814 110170 -1578 110406
rect -1814 109850 -1578 110086
rect -1814 74170 -1578 74406
rect -1814 73850 -1578 74086
rect -1814 38170 -1578 38406
rect -1814 37850 -1578 38086
rect -1814 2170 -1578 2406
rect -1814 1850 -1578 2086
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686170 1222 686406
rect 986 685850 1222 686086
rect 986 650170 1222 650406
rect 986 649850 1222 650086
rect 986 614170 1222 614406
rect 986 613850 1222 614086
rect 986 578170 1222 578406
rect 986 577850 1222 578086
rect 986 542170 1222 542406
rect 986 541850 1222 542086
rect 986 506170 1222 506406
rect 986 505850 1222 506086
rect 986 470170 1222 470406
rect 986 469850 1222 470086
rect 986 434170 1222 434406
rect 986 433850 1222 434086
rect 986 398170 1222 398406
rect 986 397850 1222 398086
rect 986 362170 1222 362406
rect 986 361850 1222 362086
rect 986 326170 1222 326406
rect 986 325850 1222 326086
rect 986 290170 1222 290406
rect 986 289850 1222 290086
rect 986 254170 1222 254406
rect 986 253850 1222 254086
rect 986 218170 1222 218406
rect 986 217850 1222 218086
rect 986 182170 1222 182406
rect 986 181850 1222 182086
rect 986 146170 1222 146406
rect 986 145850 1222 146086
rect 986 110170 1222 110406
rect 986 109850 1222 110086
rect 986 74170 1222 74406
rect 986 73850 1222 74086
rect 986 38170 1222 38406
rect 986 37850 1222 38086
rect 986 2170 1222 2406
rect 986 1850 1222 2086
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2754 -1522 -2518 -1286
rect -2754 -1842 -2518 -1606
rect 29786 711182 30022 711418
rect 29786 710862 30022 711098
rect 26186 709302 26422 709538
rect 26186 708982 26422 709218
rect 22586 707422 22822 707658
rect 22586 707102 22822 707338
rect 18986 705542 19222 705778
rect 18986 705222 19222 705458
rect 47786 710242 48022 710478
rect 47786 709922 48022 710158
rect 44186 708362 44422 708598
rect 44186 708042 44422 708278
rect 40586 706482 40822 706718
rect 40586 706162 40822 706398
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 65786 711182 66022 711418
rect 65786 710862 66022 711098
rect 62186 709302 62422 709538
rect 62186 708982 62422 709218
rect 58586 707422 58822 707658
rect 58586 707102 58822 707338
rect 54986 705542 55222 705778
rect 54986 705222 55222 705458
rect 83786 710242 84022 710478
rect 83786 709922 84022 710158
rect 80186 708362 80422 708598
rect 80186 708042 80422 708278
rect 76586 706482 76822 706718
rect 76586 706162 76822 706398
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 101786 711182 102022 711418
rect 101786 710862 102022 711098
rect 98186 709302 98422 709538
rect 98186 708982 98422 709218
rect 94586 707422 94822 707658
rect 94586 707102 94822 707338
rect 90986 705542 91222 705778
rect 90986 705222 91222 705458
rect 119786 710242 120022 710478
rect 119786 709922 120022 710158
rect 116186 708362 116422 708598
rect 116186 708042 116422 708278
rect 112586 706482 112822 706718
rect 112586 706162 112822 706398
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 137786 711182 138022 711418
rect 137786 710862 138022 711098
rect 134186 709302 134422 709538
rect 134186 708982 134422 709218
rect 130586 707422 130822 707658
rect 130586 707102 130822 707338
rect 126986 705542 127222 705778
rect 126986 705222 127222 705458
rect 155786 710242 156022 710478
rect 155786 709922 156022 710158
rect 152186 708362 152422 708598
rect 152186 708042 152422 708278
rect 148586 706482 148822 706718
rect 148586 706162 148822 706398
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 173786 711182 174022 711418
rect 173786 710862 174022 711098
rect 170186 709302 170422 709538
rect 170186 708982 170422 709218
rect 166586 707422 166822 707658
rect 166586 707102 166822 707338
rect 162986 705542 163222 705778
rect 162986 705222 163222 705458
rect 191786 710242 192022 710478
rect 191786 709922 192022 710158
rect 188186 708362 188422 708598
rect 188186 708042 188422 708278
rect 184586 706482 184822 706718
rect 184586 706162 184822 706398
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 209786 711182 210022 711418
rect 209786 710862 210022 711098
rect 206186 709302 206422 709538
rect 206186 708982 206422 709218
rect 202586 707422 202822 707658
rect 202586 707102 202822 707338
rect 198986 705542 199222 705778
rect 198986 705222 199222 705458
rect 227786 710242 228022 710478
rect 227786 709922 228022 710158
rect 224186 708362 224422 708598
rect 224186 708042 224422 708278
rect 220586 706482 220822 706718
rect 220586 706162 220822 706398
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 245786 711182 246022 711418
rect 245786 710862 246022 711098
rect 242186 709302 242422 709538
rect 242186 708982 242422 709218
rect 238586 707422 238822 707658
rect 238586 707102 238822 707338
rect 234986 705542 235222 705778
rect 234986 705222 235222 705458
rect 263786 710242 264022 710478
rect 263786 709922 264022 710158
rect 260186 708362 260422 708598
rect 260186 708042 260422 708278
rect 256586 706482 256822 706718
rect 256586 706162 256822 706398
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 281786 711182 282022 711418
rect 281786 710862 282022 711098
rect 278186 709302 278422 709538
rect 278186 708982 278422 709218
rect 274586 707422 274822 707658
rect 274586 707102 274822 707338
rect 270986 705542 271222 705778
rect 270986 705222 271222 705458
rect 299786 710242 300022 710478
rect 299786 709922 300022 710158
rect 296186 708362 296422 708598
rect 296186 708042 296422 708278
rect 292586 706482 292822 706718
rect 292586 706162 292822 706398
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 317786 711182 318022 711418
rect 317786 710862 318022 711098
rect 314186 709302 314422 709538
rect 314186 708982 314422 709218
rect 310586 707422 310822 707658
rect 310586 707102 310822 707338
rect 306986 705542 307222 705778
rect 306986 705222 307222 705458
rect 335786 710242 336022 710478
rect 335786 709922 336022 710158
rect 332186 708362 332422 708598
rect 332186 708042 332422 708278
rect 328586 706482 328822 706718
rect 328586 706162 328822 706398
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 353786 711182 354022 711418
rect 353786 710862 354022 711098
rect 350186 709302 350422 709538
rect 350186 708982 350422 709218
rect 346586 707422 346822 707658
rect 346586 707102 346822 707338
rect 342986 705542 343222 705778
rect 342986 705222 343222 705458
rect 371786 710242 372022 710478
rect 371786 709922 372022 710158
rect 368186 708362 368422 708598
rect 368186 708042 368422 708278
rect 364586 706482 364822 706718
rect 364586 706162 364822 706398
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 389786 711182 390022 711418
rect 389786 710862 390022 711098
rect 386186 709302 386422 709538
rect 386186 708982 386422 709218
rect 382586 707422 382822 707658
rect 382586 707102 382822 707338
rect 378986 705542 379222 705778
rect 378986 705222 379222 705458
rect 407786 710242 408022 710478
rect 407786 709922 408022 710158
rect 404186 708362 404422 708598
rect 404186 708042 404422 708278
rect 400586 706482 400822 706718
rect 400586 706162 400822 706398
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 425786 711182 426022 711418
rect 425786 710862 426022 711098
rect 422186 709302 422422 709538
rect 422186 708982 422422 709218
rect 418586 707422 418822 707658
rect 418586 707102 418822 707338
rect 414986 705542 415222 705778
rect 414986 705222 415222 705458
rect 443786 710242 444022 710478
rect 443786 709922 444022 710158
rect 440186 708362 440422 708598
rect 440186 708042 440422 708278
rect 436586 706482 436822 706718
rect 436586 706162 436822 706398
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 461786 711182 462022 711418
rect 461786 710862 462022 711098
rect 458186 709302 458422 709538
rect 458186 708982 458422 709218
rect 454586 707422 454822 707658
rect 454586 707102 454822 707338
rect 450986 705542 451222 705778
rect 450986 705222 451222 705458
rect 479786 710242 480022 710478
rect 479786 709922 480022 710158
rect 476186 708362 476422 708598
rect 476186 708042 476422 708278
rect 472586 706482 472822 706718
rect 472586 706162 472822 706398
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 497786 711182 498022 711418
rect 497786 710862 498022 711098
rect 494186 709302 494422 709538
rect 494186 708982 494422 709218
rect 490586 707422 490822 707658
rect 490586 707102 490822 707338
rect 486986 705542 487222 705778
rect 486986 705222 487222 705458
rect 515786 710242 516022 710478
rect 515786 709922 516022 710158
rect 512186 708362 512422 708598
rect 512186 708042 512422 708278
rect 508586 706482 508822 706718
rect 508586 706162 508822 706398
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 37142 692462 37378 692698
rect 46710 692462 46946 692698
rect 56462 692462 56698 692698
rect 66030 692462 66266 692698
rect 75782 692462 76018 692698
rect 84246 692462 84482 692698
rect 108718 692462 108954 692698
rect 114054 692462 114290 692698
rect 124174 692462 124410 692698
rect 133374 692462 133610 692698
rect 143678 692462 143914 692698
rect 152694 692462 152930 692698
rect 533786 711182 534022 711418
rect 533786 710862 534022 711098
rect 530186 709302 530422 709538
rect 530186 708982 530422 709218
rect 526586 707422 526822 707658
rect 526586 707102 526822 707338
rect 522986 705542 523222 705778
rect 522986 705222 523222 705458
rect 551786 710242 552022 710478
rect 551786 709922 552022 710158
rect 548186 708362 548422 708598
rect 548186 708042 548422 708278
rect 544586 706482 544822 706718
rect 544586 706162 544822 706398
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 569786 711182 570022 711418
rect 569786 710862 570022 711098
rect 566186 709302 566422 709538
rect 566186 708982 566422 709218
rect 562586 707422 562822 707658
rect 562586 707102 562822 707338
rect 558986 705542 559222 705778
rect 558986 705222 559222 705458
rect 592082 711182 592318 711418
rect 592082 710862 592318 711098
rect 591142 710242 591378 710478
rect 591142 709922 591378 710158
rect 590202 709302 590438 709538
rect 590202 708982 590438 709218
rect 589262 708362 589498 708598
rect 589262 708042 589498 708278
rect 588322 707422 588558 707658
rect 588322 707102 588558 707338
rect 580586 706482 580822 706718
rect 580586 706162 580822 706398
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 539462 692462 539698 692698
rect 549030 692462 549266 692698
rect 558782 692462 559018 692698
rect 565590 692462 565826 692698
rect 4586 689818 4822 690054
rect 4586 689498 4822 689734
rect 4586 653818 4822 654054
rect 4586 653498 4822 653734
rect 4586 617818 4822 618054
rect 4586 617498 4822 617734
rect 4586 581818 4822 582054
rect 4586 581498 4822 581734
rect 4586 545818 4822 546054
rect 4586 545498 4822 545734
rect 4586 509818 4822 510054
rect 4586 509498 4822 509734
rect 4586 473818 4822 474054
rect 4586 473498 4822 473734
rect 4586 437818 4822 438054
rect 4586 437498 4822 437734
rect 4586 401818 4822 402054
rect 4586 401498 4822 401734
rect 4586 365818 4822 366054
rect 4586 365498 4822 365734
rect 4586 329818 4822 330054
rect 4586 329498 4822 329734
rect 4586 293818 4822 294054
rect 4586 293498 4822 293734
rect 4586 257818 4822 258054
rect 4586 257498 4822 257734
rect 4586 221818 4822 222054
rect 4586 221498 4822 221734
rect 4586 185818 4822 186054
rect 4586 185498 4822 185734
rect 4586 149818 4822 150054
rect 4586 149498 4822 149734
rect 4586 113818 4822 114054
rect 4586 113498 4822 113734
rect 4586 77818 4822 78054
rect 4586 77498 4822 77734
rect 4586 41818 4822 42054
rect 4586 41498 4822 41734
rect 4586 5818 4822 6054
rect 587382 706482 587618 706718
rect 587382 706162 587618 706398
rect 586442 705542 586678 705778
rect 586442 705222 586678 705458
rect 580586 689818 580822 690054
rect 580586 689498 580822 689734
rect 580586 653818 580822 654054
rect 580586 653498 580822 653734
rect 580586 617818 580822 618054
rect 580586 617498 580822 617734
rect 580586 581818 580822 582054
rect 580586 581498 580822 581734
rect 580586 545818 580822 546054
rect 580586 545498 580822 545734
rect 580586 509818 580822 510054
rect 580586 509498 580822 509734
rect 580586 473818 580822 474054
rect 580586 473498 580822 473734
rect 580586 437818 580822 438054
rect 580586 437498 580822 437734
rect 580586 401818 580822 402054
rect 580586 401498 580822 401734
rect 580586 365818 580822 366054
rect 580586 365498 580822 365734
rect 580586 329818 580822 330054
rect 580586 329498 580822 329734
rect 580586 293818 580822 294054
rect 580586 293498 580822 293734
rect 580586 257818 580822 258054
rect 580586 257498 580822 257734
rect 580586 221818 580822 222054
rect 580586 221498 580822 221734
rect 580586 185818 580822 186054
rect 580586 185498 580822 185734
rect 580586 149818 580822 150054
rect 580586 149498 580822 149734
rect 580586 113818 580822 114054
rect 580586 113498 580822 113734
rect 580586 77818 580822 78054
rect 580586 77498 580822 77734
rect 580586 41818 580822 42054
rect 580586 41498 580822 41734
rect 4586 5498 4822 5734
rect -3694 -2462 -3458 -2226
rect -3694 -2782 -3458 -2546
rect 4586 -2462 4822 -2226
rect 4586 -2782 4822 -2546
rect -4634 -3402 -4398 -3166
rect -4634 -3722 -4398 -3486
rect -5574 -4342 -5338 -4106
rect -5574 -4662 -5338 -4426
rect 8186 -4342 8422 -4106
rect 8186 -4662 8422 -4426
rect -6514 -5282 -6278 -5046
rect -6514 -5602 -6278 -5366
rect -7454 -6222 -7218 -5986
rect -7454 -6542 -7218 -6306
rect 18986 -1522 19222 -1286
rect 18986 -1842 19222 -1606
rect 22586 -3402 22822 -3166
rect 22586 -3722 22822 -3486
rect 26186 -5282 26422 -5046
rect 26186 -5602 26422 -5366
rect 11786 -6222 12022 -5986
rect 11786 -6542 12022 -6306
rect -8394 -7162 -8158 -6926
rect -8394 -7482 -8158 -7246
rect 36986 2208 37222 2406
rect 36986 2170 36992 2208
rect 36992 2170 37056 2208
rect 37056 2170 37072 2208
rect 37072 2170 37136 2208
rect 37136 2170 37152 2208
rect 37152 2170 37216 2208
rect 37216 2170 37222 2208
rect 36986 1850 37222 2086
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 40586 -2462 40822 -2226
rect 40586 -2782 40822 -2546
rect 44186 -4342 44422 -4106
rect 44186 -4662 44422 -4426
rect 29786 -7162 30022 -6926
rect 29786 -7482 30022 -7246
rect 54986 -1522 55222 -1286
rect 54986 -1842 55222 -1606
rect 58586 -3402 58822 -3166
rect 58586 -3722 58822 -3486
rect 62186 -5282 62422 -5046
rect 62186 -5602 62422 -5366
rect 47786 -6222 48022 -5986
rect 47786 -6542 48022 -6306
rect 72986 2208 73222 2406
rect 72986 2170 72992 2208
rect 72992 2170 73056 2208
rect 73056 2170 73072 2208
rect 73072 2170 73136 2208
rect 73136 2170 73152 2208
rect 73152 2170 73216 2208
rect 73216 2170 73222 2208
rect 72986 1850 73222 2086
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76586 -2462 76822 -2226
rect 76586 -2782 76822 -2546
rect 80186 -4342 80422 -4106
rect 80186 -4662 80422 -4426
rect 65786 -7162 66022 -6926
rect 65786 -7482 66022 -7246
rect 90986 -1522 91222 -1286
rect 90986 -1842 91222 -1606
rect 94586 -3402 94822 -3166
rect 94586 -3722 94822 -3486
rect 98186 -5282 98422 -5046
rect 98186 -5602 98422 -5366
rect 83786 -6222 84022 -5986
rect 83786 -6542 84022 -6306
rect 108986 2208 109222 2406
rect 108986 2170 108992 2208
rect 108992 2170 109056 2208
rect 109056 2170 109072 2208
rect 109072 2170 109136 2208
rect 109136 2170 109152 2208
rect 109152 2170 109216 2208
rect 109216 2170 109222 2208
rect 108986 1850 109222 2086
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112586 -2462 112822 -2226
rect 112586 -2782 112822 -2546
rect 116186 -4342 116422 -4106
rect 116186 -4662 116422 -4426
rect 101786 -7162 102022 -6926
rect 101786 -7482 102022 -7246
rect 126986 -1522 127222 -1286
rect 126986 -1842 127222 -1606
rect 130586 -3402 130822 -3166
rect 130586 -3722 130822 -3486
rect 134186 -5282 134422 -5046
rect 134186 -5602 134422 -5366
rect 119786 -6222 120022 -5986
rect 119786 -6542 120022 -6306
rect 144986 2208 145222 2406
rect 144986 2170 144992 2208
rect 144992 2170 145056 2208
rect 145056 2170 145072 2208
rect 145072 2170 145136 2208
rect 145136 2170 145152 2208
rect 145152 2170 145216 2208
rect 145216 2170 145222 2208
rect 144986 1850 145222 2086
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148586 -2462 148822 -2226
rect 148586 -2782 148822 -2546
rect 152186 -4342 152422 -4106
rect 152186 -4662 152422 -4426
rect 137786 -7162 138022 -6926
rect 137786 -7482 138022 -7246
rect 162986 -1522 163222 -1286
rect 162986 -1842 163222 -1606
rect 166586 -3402 166822 -3166
rect 166586 -3722 166822 -3486
rect 170186 -5282 170422 -5046
rect 170186 -5602 170422 -5366
rect 155786 -6222 156022 -5986
rect 155786 -6542 156022 -6306
rect 180986 2208 181222 2406
rect 180986 2170 180992 2208
rect 180992 2170 181056 2208
rect 181056 2170 181072 2208
rect 181072 2170 181136 2208
rect 181136 2170 181152 2208
rect 181152 2170 181216 2208
rect 181216 2170 181222 2208
rect 180986 1850 181222 2086
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 -2462 184822 -2226
rect 184586 -2782 184822 -2546
rect 188186 -4342 188422 -4106
rect 188186 -4662 188422 -4426
rect 173786 -7162 174022 -6926
rect 173786 -7482 174022 -7246
rect 198986 -1522 199222 -1286
rect 198986 -1842 199222 -1606
rect 202586 -3402 202822 -3166
rect 202586 -3722 202822 -3486
rect 206186 -5282 206422 -5046
rect 206186 -5602 206422 -5366
rect 191786 -6222 192022 -5986
rect 191786 -6542 192022 -6306
rect 216986 2208 217222 2406
rect 216986 2170 216992 2208
rect 216992 2170 217056 2208
rect 217056 2170 217072 2208
rect 217072 2170 217136 2208
rect 217136 2170 217152 2208
rect 217152 2170 217216 2208
rect 217216 2170 217222 2208
rect 216986 1850 217222 2086
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 -2462 220822 -2226
rect 220586 -2782 220822 -2546
rect 224186 -4342 224422 -4106
rect 224186 -4662 224422 -4426
rect 209786 -7162 210022 -6926
rect 209786 -7482 210022 -7246
rect 234986 -1522 235222 -1286
rect 234986 -1842 235222 -1606
rect 238586 -3402 238822 -3166
rect 238586 -3722 238822 -3486
rect 242186 -5282 242422 -5046
rect 242186 -5602 242422 -5366
rect 227786 -6222 228022 -5986
rect 227786 -6542 228022 -6306
rect 252986 2208 253222 2406
rect 252986 2170 252992 2208
rect 252992 2170 253056 2208
rect 253056 2170 253072 2208
rect 253072 2170 253136 2208
rect 253136 2170 253152 2208
rect 253152 2170 253216 2208
rect 253216 2170 253222 2208
rect 252986 1850 253222 2086
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256586 -2462 256822 -2226
rect 256586 -2782 256822 -2546
rect 260186 -4342 260422 -4106
rect 260186 -4662 260422 -4426
rect 245786 -7162 246022 -6926
rect 245786 -7482 246022 -7246
rect 270986 -1522 271222 -1286
rect 270986 -1842 271222 -1606
rect 274586 -3402 274822 -3166
rect 274586 -3722 274822 -3486
rect 278186 -5282 278422 -5046
rect 278186 -5602 278422 -5366
rect 263786 -6222 264022 -5986
rect 263786 -6542 264022 -6306
rect 288986 2208 289222 2406
rect 288986 2170 288992 2208
rect 288992 2170 289056 2208
rect 289056 2170 289072 2208
rect 289072 2170 289136 2208
rect 289136 2170 289152 2208
rect 289152 2170 289216 2208
rect 289216 2170 289222 2208
rect 288986 1850 289222 2086
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 -2462 292822 -2226
rect 292586 -2782 292822 -2546
rect 296186 -4342 296422 -4106
rect 296186 -4662 296422 -4426
rect 281786 -7162 282022 -6926
rect 281786 -7482 282022 -7246
rect 306986 -1522 307222 -1286
rect 306986 -1842 307222 -1606
rect 310586 -3402 310822 -3166
rect 310586 -3722 310822 -3486
rect 314186 -5282 314422 -5046
rect 314186 -5602 314422 -5366
rect 299786 -6222 300022 -5986
rect 299786 -6542 300022 -6306
rect 324986 2208 325222 2406
rect 324986 2170 324992 2208
rect 324992 2170 325056 2208
rect 325056 2170 325072 2208
rect 325072 2170 325136 2208
rect 325136 2170 325152 2208
rect 325152 2170 325216 2208
rect 325216 2170 325222 2208
rect 324986 1850 325222 2086
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328586 -2462 328822 -2226
rect 328586 -2782 328822 -2546
rect 332186 -4342 332422 -4106
rect 332186 -4662 332422 -4426
rect 317786 -7162 318022 -6926
rect 317786 -7482 318022 -7246
rect 342986 -1522 343222 -1286
rect 342986 -1842 343222 -1606
rect 346586 -3402 346822 -3166
rect 346586 -3722 346822 -3486
rect 350186 -5282 350422 -5046
rect 350186 -5602 350422 -5366
rect 335786 -6222 336022 -5986
rect 335786 -6542 336022 -6306
rect 360986 2208 361222 2406
rect 360986 2170 360992 2208
rect 360992 2170 361056 2208
rect 361056 2170 361072 2208
rect 361072 2170 361136 2208
rect 361136 2170 361152 2208
rect 361152 2170 361216 2208
rect 361216 2170 361222 2208
rect 360986 1850 361222 2086
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 -2462 364822 -2226
rect 364586 -2782 364822 -2546
rect 368186 -4342 368422 -4106
rect 368186 -4662 368422 -4426
rect 353786 -7162 354022 -6926
rect 353786 -7482 354022 -7246
rect 378986 -1522 379222 -1286
rect 378986 -1842 379222 -1606
rect 382586 -3402 382822 -3166
rect 382586 -3722 382822 -3486
rect 386186 -5282 386422 -5046
rect 386186 -5602 386422 -5366
rect 371786 -6222 372022 -5986
rect 371786 -6542 372022 -6306
rect 396986 2208 397222 2406
rect 396986 2170 396992 2208
rect 396992 2170 397056 2208
rect 397056 2170 397072 2208
rect 397072 2170 397136 2208
rect 397136 2170 397152 2208
rect 397152 2170 397216 2208
rect 397216 2170 397222 2208
rect 396986 1850 397222 2086
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400586 -2462 400822 -2226
rect 400586 -2782 400822 -2546
rect 404186 -4342 404422 -4106
rect 404186 -4662 404422 -4426
rect 389786 -7162 390022 -6926
rect 389786 -7482 390022 -7246
rect 414986 -1522 415222 -1286
rect 414986 -1842 415222 -1606
rect 418586 -3402 418822 -3166
rect 418586 -3722 418822 -3486
rect 422186 -5282 422422 -5046
rect 422186 -5602 422422 -5366
rect 407786 -6222 408022 -5986
rect 407786 -6542 408022 -6306
rect 432986 2208 433222 2406
rect 432986 2170 432992 2208
rect 432992 2170 433056 2208
rect 433056 2170 433072 2208
rect 433072 2170 433136 2208
rect 433136 2170 433152 2208
rect 433152 2170 433216 2208
rect 433216 2170 433222 2208
rect 432986 1850 433222 2086
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436586 -2462 436822 -2226
rect 436586 -2782 436822 -2546
rect 440186 -4342 440422 -4106
rect 440186 -4662 440422 -4426
rect 425786 -7162 426022 -6926
rect 425786 -7482 426022 -7246
rect 450986 -1522 451222 -1286
rect 450986 -1842 451222 -1606
rect 454586 -3402 454822 -3166
rect 454586 -3722 454822 -3486
rect 458186 -5282 458422 -5046
rect 458186 -5602 458422 -5366
rect 443786 -6222 444022 -5986
rect 443786 -6542 444022 -6306
rect 468986 2208 469222 2406
rect 468986 2170 468992 2208
rect 468992 2170 469056 2208
rect 469056 2170 469072 2208
rect 469072 2170 469136 2208
rect 469136 2170 469152 2208
rect 469152 2170 469216 2208
rect 469216 2170 469222 2208
rect 468986 1850 469222 2086
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472586 -2462 472822 -2226
rect 472586 -2782 472822 -2546
rect 476186 -4342 476422 -4106
rect 476186 -4662 476422 -4426
rect 461786 -7162 462022 -6926
rect 461786 -7482 462022 -7246
rect 486986 -1522 487222 -1286
rect 486986 -1842 487222 -1606
rect 490586 -3402 490822 -3166
rect 490586 -3722 490822 -3486
rect 494186 -5282 494422 -5046
rect 494186 -5602 494422 -5366
rect 479786 -6222 480022 -5986
rect 479786 -6542 480022 -6306
rect 504986 2208 505222 2406
rect 504986 2170 504992 2208
rect 504992 2170 505056 2208
rect 505056 2170 505072 2208
rect 505072 2170 505136 2208
rect 505136 2170 505152 2208
rect 505152 2170 505216 2208
rect 505216 2170 505222 2208
rect 504986 1850 505222 2086
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508586 -2462 508822 -2226
rect 508586 -2782 508822 -2546
rect 512186 -4342 512422 -4106
rect 512186 -4662 512422 -4426
rect 497786 -7162 498022 -6926
rect 497786 -7482 498022 -7246
rect 522986 -1522 523222 -1286
rect 522986 -1842 523222 -1606
rect 526586 -3402 526822 -3166
rect 526586 -3722 526822 -3486
rect 530186 -5282 530422 -5046
rect 530186 -5602 530422 -5366
rect 515786 -6222 516022 -5986
rect 515786 -6542 516022 -6306
rect 540986 2208 541222 2406
rect 540986 2170 540992 2208
rect 540992 2170 541056 2208
rect 541056 2170 541072 2208
rect 541072 2170 541136 2208
rect 541136 2170 541152 2208
rect 541152 2170 541216 2208
rect 541216 2170 541222 2208
rect 540986 1850 541222 2086
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544586 -2462 544822 -2226
rect 544586 -2782 544822 -2546
rect 548186 -4342 548422 -4106
rect 548186 -4662 548422 -4426
rect 533786 -7162 534022 -6926
rect 533786 -7482 534022 -7246
rect 558986 -1522 559222 -1286
rect 558986 -1842 559222 -1606
rect 562586 -3402 562822 -3166
rect 562586 -3722 562822 -3486
rect 566186 -5282 566422 -5046
rect 566186 -5602 566422 -5366
rect 551786 -6222 552022 -5986
rect 551786 -6542 552022 -6306
rect 576986 2208 577222 2406
rect 576986 2170 576992 2208
rect 576992 2170 577056 2208
rect 577056 2170 577072 2208
rect 577072 2170 577136 2208
rect 577136 2170 577152 2208
rect 577152 2170 577216 2208
rect 577216 2170 577222 2208
rect 576986 1850 577222 2086
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 580586 5818 580822 6054
rect 580586 5498 580822 5734
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686170 585738 686406
rect 585502 685850 585738 686086
rect 585502 650170 585738 650406
rect 585502 649850 585738 650086
rect 585502 614170 585738 614406
rect 585502 613850 585738 614086
rect 585502 578170 585738 578406
rect 585502 577850 585738 578086
rect 585502 542170 585738 542406
rect 585502 541850 585738 542086
rect 585502 506170 585738 506406
rect 585502 505850 585738 506086
rect 585502 470170 585738 470406
rect 585502 469850 585738 470086
rect 585502 434170 585738 434406
rect 585502 433850 585738 434086
rect 585502 398170 585738 398406
rect 585502 397850 585738 398086
rect 585502 362170 585738 362406
rect 585502 361850 585738 362086
rect 585502 326170 585738 326406
rect 585502 325850 585738 326086
rect 585502 290170 585738 290406
rect 585502 289850 585738 290086
rect 585502 254170 585738 254406
rect 585502 253850 585738 254086
rect 585502 218170 585738 218406
rect 585502 217850 585738 218086
rect 585502 182170 585738 182406
rect 585502 181850 585738 182086
rect 585502 146170 585738 146406
rect 585502 145850 585738 146086
rect 585502 110170 585738 110406
rect 585502 109850 585738 110086
rect 585502 74170 585738 74406
rect 585502 73850 585738 74086
rect 585502 38170 585738 38406
rect 585502 37850 585738 38086
rect 585502 2170 585738 2406
rect 585502 1850 585738 2086
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586442 668170 586678 668406
rect 586442 667850 586678 668086
rect 586442 632170 586678 632406
rect 586442 631850 586678 632086
rect 586442 596170 586678 596406
rect 586442 595850 586678 596086
rect 586442 560170 586678 560406
rect 586442 559850 586678 560086
rect 586442 524170 586678 524406
rect 586442 523850 586678 524086
rect 586442 488170 586678 488406
rect 586442 487850 586678 488086
rect 586442 452170 586678 452406
rect 586442 451850 586678 452086
rect 586442 416170 586678 416406
rect 586442 415850 586678 416086
rect 586442 380170 586678 380406
rect 586442 379850 586678 380086
rect 586442 344170 586678 344406
rect 586442 343850 586678 344086
rect 586442 308170 586678 308406
rect 586442 307850 586678 308086
rect 586442 272170 586678 272406
rect 586442 271850 586678 272086
rect 586442 236170 586678 236406
rect 586442 235850 586678 236086
rect 586442 200170 586678 200406
rect 586442 199850 586678 200086
rect 586442 164170 586678 164406
rect 586442 163850 586678 164086
rect 586442 128170 586678 128406
rect 586442 127850 586678 128086
rect 586442 92170 586678 92406
rect 586442 91850 586678 92086
rect 586442 56170 586678 56406
rect 586442 55850 586678 56086
rect 586442 20170 586678 20406
rect 586442 19850 586678 20086
rect 586442 -1522 586678 -1286
rect 586442 -1842 586678 -1606
rect 587382 689818 587618 690054
rect 587382 689498 587618 689734
rect 587382 653818 587618 654054
rect 587382 653498 587618 653734
rect 587382 617818 587618 618054
rect 587382 617498 587618 617734
rect 587382 581818 587618 582054
rect 587382 581498 587618 581734
rect 587382 545818 587618 546054
rect 587382 545498 587618 545734
rect 587382 509818 587618 510054
rect 587382 509498 587618 509734
rect 587382 473818 587618 474054
rect 587382 473498 587618 473734
rect 587382 437818 587618 438054
rect 587382 437498 587618 437734
rect 587382 401818 587618 402054
rect 587382 401498 587618 401734
rect 587382 365818 587618 366054
rect 587382 365498 587618 365734
rect 587382 329818 587618 330054
rect 587382 329498 587618 329734
rect 587382 293818 587618 294054
rect 587382 293498 587618 293734
rect 587382 257818 587618 258054
rect 587382 257498 587618 257734
rect 587382 221818 587618 222054
rect 587382 221498 587618 221734
rect 587382 185818 587618 186054
rect 587382 185498 587618 185734
rect 587382 149818 587618 150054
rect 587382 149498 587618 149734
rect 587382 113818 587618 114054
rect 587382 113498 587618 113734
rect 587382 77818 587618 78054
rect 587382 77498 587618 77734
rect 587382 41818 587618 42054
rect 587382 41498 587618 41734
rect 587382 5818 587618 6054
rect 587382 5498 587618 5734
rect 580586 -2462 580822 -2226
rect 580586 -2782 580822 -2546
rect 587382 -2462 587618 -2226
rect 587382 -2782 587618 -2546
rect 588322 671818 588558 672054
rect 588322 671498 588558 671734
rect 588322 635818 588558 636054
rect 588322 635498 588558 635734
rect 588322 599818 588558 600054
rect 588322 599498 588558 599734
rect 588322 563818 588558 564054
rect 588322 563498 588558 563734
rect 588322 527818 588558 528054
rect 588322 527498 588558 527734
rect 588322 491818 588558 492054
rect 588322 491498 588558 491734
rect 588322 455818 588558 456054
rect 588322 455498 588558 455734
rect 588322 419818 588558 420054
rect 588322 419498 588558 419734
rect 588322 383818 588558 384054
rect 588322 383498 588558 383734
rect 588322 347818 588558 348054
rect 588322 347498 588558 347734
rect 588322 311818 588558 312054
rect 588322 311498 588558 311734
rect 588322 275818 588558 276054
rect 588322 275498 588558 275734
rect 588322 239818 588558 240054
rect 588322 239498 588558 239734
rect 588322 203818 588558 204054
rect 588322 203498 588558 203734
rect 588322 167818 588558 168054
rect 588322 167498 588558 167734
rect 588322 131818 588558 132054
rect 588322 131498 588558 131734
rect 588322 95818 588558 96054
rect 588322 95498 588558 95734
rect 588322 59818 588558 60054
rect 588322 59498 588558 59734
rect 588322 23818 588558 24054
rect 588322 23498 588558 23734
rect 588322 -3402 588558 -3166
rect 588322 -3722 588558 -3486
rect 589262 693418 589498 693654
rect 589262 693098 589498 693334
rect 589262 657418 589498 657654
rect 589262 657098 589498 657334
rect 589262 621418 589498 621654
rect 589262 621098 589498 621334
rect 589262 585418 589498 585654
rect 589262 585098 589498 585334
rect 589262 549418 589498 549654
rect 589262 549098 589498 549334
rect 589262 513418 589498 513654
rect 589262 513098 589498 513334
rect 589262 477418 589498 477654
rect 589262 477098 589498 477334
rect 589262 441418 589498 441654
rect 589262 441098 589498 441334
rect 589262 405418 589498 405654
rect 589262 405098 589498 405334
rect 589262 369418 589498 369654
rect 589262 369098 589498 369334
rect 589262 333418 589498 333654
rect 589262 333098 589498 333334
rect 589262 297418 589498 297654
rect 589262 297098 589498 297334
rect 589262 261418 589498 261654
rect 589262 261098 589498 261334
rect 589262 225418 589498 225654
rect 589262 225098 589498 225334
rect 589262 189418 589498 189654
rect 589262 189098 589498 189334
rect 589262 153418 589498 153654
rect 589262 153098 589498 153334
rect 589262 117418 589498 117654
rect 589262 117098 589498 117334
rect 589262 81418 589498 81654
rect 589262 81098 589498 81334
rect 589262 45418 589498 45654
rect 589262 45098 589498 45334
rect 589262 9418 589498 9654
rect 589262 9098 589498 9334
rect 589262 -4342 589498 -4106
rect 589262 -4662 589498 -4426
rect 590202 675418 590438 675654
rect 590202 675098 590438 675334
rect 590202 639418 590438 639654
rect 590202 639098 590438 639334
rect 590202 603418 590438 603654
rect 590202 603098 590438 603334
rect 590202 567418 590438 567654
rect 590202 567098 590438 567334
rect 590202 531418 590438 531654
rect 590202 531098 590438 531334
rect 590202 495418 590438 495654
rect 590202 495098 590438 495334
rect 590202 459418 590438 459654
rect 590202 459098 590438 459334
rect 590202 423418 590438 423654
rect 590202 423098 590438 423334
rect 590202 387418 590438 387654
rect 590202 387098 590438 387334
rect 590202 351418 590438 351654
rect 590202 351098 590438 351334
rect 590202 315418 590438 315654
rect 590202 315098 590438 315334
rect 590202 279418 590438 279654
rect 590202 279098 590438 279334
rect 590202 243418 590438 243654
rect 590202 243098 590438 243334
rect 590202 207418 590438 207654
rect 590202 207098 590438 207334
rect 590202 171418 590438 171654
rect 590202 171098 590438 171334
rect 590202 135418 590438 135654
rect 590202 135098 590438 135334
rect 590202 99418 590438 99654
rect 590202 99098 590438 99334
rect 590202 63418 590438 63654
rect 590202 63098 590438 63334
rect 590202 27418 590438 27654
rect 590202 27098 590438 27334
rect 590202 -5282 590438 -5046
rect 590202 -5602 590438 -5366
rect 591142 697018 591378 697254
rect 591142 696698 591378 696934
rect 591142 661018 591378 661254
rect 591142 660698 591378 660934
rect 591142 625018 591378 625254
rect 591142 624698 591378 624934
rect 591142 589018 591378 589254
rect 591142 588698 591378 588934
rect 591142 553018 591378 553254
rect 591142 552698 591378 552934
rect 591142 517018 591378 517254
rect 591142 516698 591378 516934
rect 591142 481018 591378 481254
rect 591142 480698 591378 480934
rect 591142 445018 591378 445254
rect 591142 444698 591378 444934
rect 591142 409018 591378 409254
rect 591142 408698 591378 408934
rect 591142 373018 591378 373254
rect 591142 372698 591378 372934
rect 591142 337018 591378 337254
rect 591142 336698 591378 336934
rect 591142 301018 591378 301254
rect 591142 300698 591378 300934
rect 591142 265018 591378 265254
rect 591142 264698 591378 264934
rect 591142 229018 591378 229254
rect 591142 228698 591378 228934
rect 591142 193018 591378 193254
rect 591142 192698 591378 192934
rect 591142 157018 591378 157254
rect 591142 156698 591378 156934
rect 591142 121018 591378 121254
rect 591142 120698 591378 120934
rect 591142 85018 591378 85254
rect 591142 84698 591378 84934
rect 591142 49018 591378 49254
rect 591142 48698 591378 48934
rect 591142 13018 591378 13254
rect 591142 12698 591378 12934
rect 591142 -6222 591378 -5986
rect 591142 -6542 591378 -6306
rect 592082 679018 592318 679254
rect 592082 678698 592318 678934
rect 592082 643018 592318 643254
rect 592082 642698 592318 642934
rect 592082 607018 592318 607254
rect 592082 606698 592318 606934
rect 592082 571018 592318 571254
rect 592082 570698 592318 570934
rect 592082 535018 592318 535254
rect 592082 534698 592318 534934
rect 592082 499018 592318 499254
rect 592082 498698 592318 498934
rect 592082 463018 592318 463254
rect 592082 462698 592318 462934
rect 592082 427018 592318 427254
rect 592082 426698 592318 426934
rect 592082 391018 592318 391254
rect 592082 390698 592318 390934
rect 592082 355018 592318 355254
rect 592082 354698 592318 354934
rect 592082 319018 592318 319254
rect 592082 318698 592318 318934
rect 592082 283018 592318 283254
rect 592082 282698 592318 282934
rect 592082 247018 592318 247254
rect 592082 246698 592318 246934
rect 592082 211018 592318 211254
rect 592082 210698 592318 210934
rect 592082 175018 592318 175254
rect 592082 174698 592318 174934
rect 592082 139018 592318 139254
rect 592082 138698 592318 138934
rect 592082 103018 592318 103254
rect 592082 102698 592318 102934
rect 592082 67018 592318 67254
rect 592082 66698 592318 66934
rect 592082 31018 592318 31254
rect 592082 30698 592318 30934
rect 569786 -7162 570022 -6926
rect 569786 -7482 570022 -7246
rect 592082 -7162 592318 -6926
rect 592082 -7482 592318 -7246
<< metal5 >>
rect -8576 711440 -7976 711442
rect 29604 711440 30204 711442
rect 65604 711440 66204 711442
rect 101604 711440 102204 711442
rect 137604 711440 138204 711442
rect 173604 711440 174204 711442
rect 209604 711440 210204 711442
rect 245604 711440 246204 711442
rect 281604 711440 282204 711442
rect 317604 711440 318204 711442
rect 353604 711440 354204 711442
rect 389604 711440 390204 711442
rect 425604 711440 426204 711442
rect 461604 711440 462204 711442
rect 497604 711440 498204 711442
rect 533604 711440 534204 711442
rect 569604 711440 570204 711442
rect 591900 711440 592500 711442
rect -8576 711418 592500 711440
rect -8576 711182 -8394 711418
rect -8158 711182 29786 711418
rect 30022 711182 65786 711418
rect 66022 711182 101786 711418
rect 102022 711182 137786 711418
rect 138022 711182 173786 711418
rect 174022 711182 209786 711418
rect 210022 711182 245786 711418
rect 246022 711182 281786 711418
rect 282022 711182 317786 711418
rect 318022 711182 353786 711418
rect 354022 711182 389786 711418
rect 390022 711182 425786 711418
rect 426022 711182 461786 711418
rect 462022 711182 497786 711418
rect 498022 711182 533786 711418
rect 534022 711182 569786 711418
rect 570022 711182 592082 711418
rect 592318 711182 592500 711418
rect -8576 711098 592500 711182
rect -8576 710862 -8394 711098
rect -8158 710862 29786 711098
rect 30022 710862 65786 711098
rect 66022 710862 101786 711098
rect 102022 710862 137786 711098
rect 138022 710862 173786 711098
rect 174022 710862 209786 711098
rect 210022 710862 245786 711098
rect 246022 710862 281786 711098
rect 282022 710862 317786 711098
rect 318022 710862 353786 711098
rect 354022 710862 389786 711098
rect 390022 710862 425786 711098
rect 426022 710862 461786 711098
rect 462022 710862 497786 711098
rect 498022 710862 533786 711098
rect 534022 710862 569786 711098
rect 570022 710862 592082 711098
rect 592318 710862 592500 711098
rect -8576 710840 592500 710862
rect -8576 710838 -7976 710840
rect 29604 710838 30204 710840
rect 65604 710838 66204 710840
rect 101604 710838 102204 710840
rect 137604 710838 138204 710840
rect 173604 710838 174204 710840
rect 209604 710838 210204 710840
rect 245604 710838 246204 710840
rect 281604 710838 282204 710840
rect 317604 710838 318204 710840
rect 353604 710838 354204 710840
rect 389604 710838 390204 710840
rect 425604 710838 426204 710840
rect 461604 710838 462204 710840
rect 497604 710838 498204 710840
rect 533604 710838 534204 710840
rect 569604 710838 570204 710840
rect 591900 710838 592500 710840
rect -7636 710500 -7036 710502
rect 11604 710500 12204 710502
rect 47604 710500 48204 710502
rect 83604 710500 84204 710502
rect 119604 710500 120204 710502
rect 155604 710500 156204 710502
rect 191604 710500 192204 710502
rect 227604 710500 228204 710502
rect 263604 710500 264204 710502
rect 299604 710500 300204 710502
rect 335604 710500 336204 710502
rect 371604 710500 372204 710502
rect 407604 710500 408204 710502
rect 443604 710500 444204 710502
rect 479604 710500 480204 710502
rect 515604 710500 516204 710502
rect 551604 710500 552204 710502
rect 590960 710500 591560 710502
rect -7636 710478 591560 710500
rect -7636 710242 -7454 710478
rect -7218 710242 11786 710478
rect 12022 710242 47786 710478
rect 48022 710242 83786 710478
rect 84022 710242 119786 710478
rect 120022 710242 155786 710478
rect 156022 710242 191786 710478
rect 192022 710242 227786 710478
rect 228022 710242 263786 710478
rect 264022 710242 299786 710478
rect 300022 710242 335786 710478
rect 336022 710242 371786 710478
rect 372022 710242 407786 710478
rect 408022 710242 443786 710478
rect 444022 710242 479786 710478
rect 480022 710242 515786 710478
rect 516022 710242 551786 710478
rect 552022 710242 591142 710478
rect 591378 710242 591560 710478
rect -7636 710158 591560 710242
rect -7636 709922 -7454 710158
rect -7218 709922 11786 710158
rect 12022 709922 47786 710158
rect 48022 709922 83786 710158
rect 84022 709922 119786 710158
rect 120022 709922 155786 710158
rect 156022 709922 191786 710158
rect 192022 709922 227786 710158
rect 228022 709922 263786 710158
rect 264022 709922 299786 710158
rect 300022 709922 335786 710158
rect 336022 709922 371786 710158
rect 372022 709922 407786 710158
rect 408022 709922 443786 710158
rect 444022 709922 479786 710158
rect 480022 709922 515786 710158
rect 516022 709922 551786 710158
rect 552022 709922 591142 710158
rect 591378 709922 591560 710158
rect -7636 709900 591560 709922
rect -7636 709898 -7036 709900
rect 11604 709898 12204 709900
rect 47604 709898 48204 709900
rect 83604 709898 84204 709900
rect 119604 709898 120204 709900
rect 155604 709898 156204 709900
rect 191604 709898 192204 709900
rect 227604 709898 228204 709900
rect 263604 709898 264204 709900
rect 299604 709898 300204 709900
rect 335604 709898 336204 709900
rect 371604 709898 372204 709900
rect 407604 709898 408204 709900
rect 443604 709898 444204 709900
rect 479604 709898 480204 709900
rect 515604 709898 516204 709900
rect 551604 709898 552204 709900
rect 590960 709898 591560 709900
rect -6696 709560 -6096 709562
rect 26004 709560 26604 709562
rect 62004 709560 62604 709562
rect 98004 709560 98604 709562
rect 134004 709560 134604 709562
rect 170004 709560 170604 709562
rect 206004 709560 206604 709562
rect 242004 709560 242604 709562
rect 278004 709560 278604 709562
rect 314004 709560 314604 709562
rect 350004 709560 350604 709562
rect 386004 709560 386604 709562
rect 422004 709560 422604 709562
rect 458004 709560 458604 709562
rect 494004 709560 494604 709562
rect 530004 709560 530604 709562
rect 566004 709560 566604 709562
rect 590020 709560 590620 709562
rect -6696 709538 590620 709560
rect -6696 709302 -6514 709538
rect -6278 709302 26186 709538
rect 26422 709302 62186 709538
rect 62422 709302 98186 709538
rect 98422 709302 134186 709538
rect 134422 709302 170186 709538
rect 170422 709302 206186 709538
rect 206422 709302 242186 709538
rect 242422 709302 278186 709538
rect 278422 709302 314186 709538
rect 314422 709302 350186 709538
rect 350422 709302 386186 709538
rect 386422 709302 422186 709538
rect 422422 709302 458186 709538
rect 458422 709302 494186 709538
rect 494422 709302 530186 709538
rect 530422 709302 566186 709538
rect 566422 709302 590202 709538
rect 590438 709302 590620 709538
rect -6696 709218 590620 709302
rect -6696 708982 -6514 709218
rect -6278 708982 26186 709218
rect 26422 708982 62186 709218
rect 62422 708982 98186 709218
rect 98422 708982 134186 709218
rect 134422 708982 170186 709218
rect 170422 708982 206186 709218
rect 206422 708982 242186 709218
rect 242422 708982 278186 709218
rect 278422 708982 314186 709218
rect 314422 708982 350186 709218
rect 350422 708982 386186 709218
rect 386422 708982 422186 709218
rect 422422 708982 458186 709218
rect 458422 708982 494186 709218
rect 494422 708982 530186 709218
rect 530422 708982 566186 709218
rect 566422 708982 590202 709218
rect 590438 708982 590620 709218
rect -6696 708960 590620 708982
rect -6696 708958 -6096 708960
rect 26004 708958 26604 708960
rect 62004 708958 62604 708960
rect 98004 708958 98604 708960
rect 134004 708958 134604 708960
rect 170004 708958 170604 708960
rect 206004 708958 206604 708960
rect 242004 708958 242604 708960
rect 278004 708958 278604 708960
rect 314004 708958 314604 708960
rect 350004 708958 350604 708960
rect 386004 708958 386604 708960
rect 422004 708958 422604 708960
rect 458004 708958 458604 708960
rect 494004 708958 494604 708960
rect 530004 708958 530604 708960
rect 566004 708958 566604 708960
rect 590020 708958 590620 708960
rect -5756 708620 -5156 708622
rect 8004 708620 8604 708622
rect 44004 708620 44604 708622
rect 80004 708620 80604 708622
rect 116004 708620 116604 708622
rect 152004 708620 152604 708622
rect 188004 708620 188604 708622
rect 224004 708620 224604 708622
rect 260004 708620 260604 708622
rect 296004 708620 296604 708622
rect 332004 708620 332604 708622
rect 368004 708620 368604 708622
rect 404004 708620 404604 708622
rect 440004 708620 440604 708622
rect 476004 708620 476604 708622
rect 512004 708620 512604 708622
rect 548004 708620 548604 708622
rect 589080 708620 589680 708622
rect -5756 708598 589680 708620
rect -5756 708362 -5574 708598
rect -5338 708362 8186 708598
rect 8422 708362 44186 708598
rect 44422 708362 80186 708598
rect 80422 708362 116186 708598
rect 116422 708362 152186 708598
rect 152422 708362 188186 708598
rect 188422 708362 224186 708598
rect 224422 708362 260186 708598
rect 260422 708362 296186 708598
rect 296422 708362 332186 708598
rect 332422 708362 368186 708598
rect 368422 708362 404186 708598
rect 404422 708362 440186 708598
rect 440422 708362 476186 708598
rect 476422 708362 512186 708598
rect 512422 708362 548186 708598
rect 548422 708362 589262 708598
rect 589498 708362 589680 708598
rect -5756 708278 589680 708362
rect -5756 708042 -5574 708278
rect -5338 708042 8186 708278
rect 8422 708042 44186 708278
rect 44422 708042 80186 708278
rect 80422 708042 116186 708278
rect 116422 708042 152186 708278
rect 152422 708042 188186 708278
rect 188422 708042 224186 708278
rect 224422 708042 260186 708278
rect 260422 708042 296186 708278
rect 296422 708042 332186 708278
rect 332422 708042 368186 708278
rect 368422 708042 404186 708278
rect 404422 708042 440186 708278
rect 440422 708042 476186 708278
rect 476422 708042 512186 708278
rect 512422 708042 548186 708278
rect 548422 708042 589262 708278
rect 589498 708042 589680 708278
rect -5756 708020 589680 708042
rect -5756 708018 -5156 708020
rect 8004 708018 8604 708020
rect 44004 708018 44604 708020
rect 80004 708018 80604 708020
rect 116004 708018 116604 708020
rect 152004 708018 152604 708020
rect 188004 708018 188604 708020
rect 224004 708018 224604 708020
rect 260004 708018 260604 708020
rect 296004 708018 296604 708020
rect 332004 708018 332604 708020
rect 368004 708018 368604 708020
rect 404004 708018 404604 708020
rect 440004 708018 440604 708020
rect 476004 708018 476604 708020
rect 512004 708018 512604 708020
rect 548004 708018 548604 708020
rect 589080 708018 589680 708020
rect -4816 707680 -4216 707682
rect 22404 707680 23004 707682
rect 58404 707680 59004 707682
rect 94404 707680 95004 707682
rect 130404 707680 131004 707682
rect 166404 707680 167004 707682
rect 202404 707680 203004 707682
rect 238404 707680 239004 707682
rect 274404 707680 275004 707682
rect 310404 707680 311004 707682
rect 346404 707680 347004 707682
rect 382404 707680 383004 707682
rect 418404 707680 419004 707682
rect 454404 707680 455004 707682
rect 490404 707680 491004 707682
rect 526404 707680 527004 707682
rect 562404 707680 563004 707682
rect 588140 707680 588740 707682
rect -4816 707658 588740 707680
rect -4816 707422 -4634 707658
rect -4398 707422 22586 707658
rect 22822 707422 58586 707658
rect 58822 707422 94586 707658
rect 94822 707422 130586 707658
rect 130822 707422 166586 707658
rect 166822 707422 202586 707658
rect 202822 707422 238586 707658
rect 238822 707422 274586 707658
rect 274822 707422 310586 707658
rect 310822 707422 346586 707658
rect 346822 707422 382586 707658
rect 382822 707422 418586 707658
rect 418822 707422 454586 707658
rect 454822 707422 490586 707658
rect 490822 707422 526586 707658
rect 526822 707422 562586 707658
rect 562822 707422 588322 707658
rect 588558 707422 588740 707658
rect -4816 707338 588740 707422
rect -4816 707102 -4634 707338
rect -4398 707102 22586 707338
rect 22822 707102 58586 707338
rect 58822 707102 94586 707338
rect 94822 707102 130586 707338
rect 130822 707102 166586 707338
rect 166822 707102 202586 707338
rect 202822 707102 238586 707338
rect 238822 707102 274586 707338
rect 274822 707102 310586 707338
rect 310822 707102 346586 707338
rect 346822 707102 382586 707338
rect 382822 707102 418586 707338
rect 418822 707102 454586 707338
rect 454822 707102 490586 707338
rect 490822 707102 526586 707338
rect 526822 707102 562586 707338
rect 562822 707102 588322 707338
rect 588558 707102 588740 707338
rect -4816 707080 588740 707102
rect -4816 707078 -4216 707080
rect 22404 707078 23004 707080
rect 58404 707078 59004 707080
rect 94404 707078 95004 707080
rect 130404 707078 131004 707080
rect 166404 707078 167004 707080
rect 202404 707078 203004 707080
rect 238404 707078 239004 707080
rect 274404 707078 275004 707080
rect 310404 707078 311004 707080
rect 346404 707078 347004 707080
rect 382404 707078 383004 707080
rect 418404 707078 419004 707080
rect 454404 707078 455004 707080
rect 490404 707078 491004 707080
rect 526404 707078 527004 707080
rect 562404 707078 563004 707080
rect 588140 707078 588740 707080
rect -3876 706740 -3276 706742
rect 4404 706740 5004 706742
rect 40404 706740 41004 706742
rect 76404 706740 77004 706742
rect 112404 706740 113004 706742
rect 148404 706740 149004 706742
rect 184404 706740 185004 706742
rect 220404 706740 221004 706742
rect 256404 706740 257004 706742
rect 292404 706740 293004 706742
rect 328404 706740 329004 706742
rect 364404 706740 365004 706742
rect 400404 706740 401004 706742
rect 436404 706740 437004 706742
rect 472404 706740 473004 706742
rect 508404 706740 509004 706742
rect 544404 706740 545004 706742
rect 580404 706740 581004 706742
rect 587200 706740 587800 706742
rect -3876 706718 587800 706740
rect -3876 706482 -3694 706718
rect -3458 706482 4586 706718
rect 4822 706482 40586 706718
rect 40822 706482 76586 706718
rect 76822 706482 112586 706718
rect 112822 706482 148586 706718
rect 148822 706482 184586 706718
rect 184822 706482 220586 706718
rect 220822 706482 256586 706718
rect 256822 706482 292586 706718
rect 292822 706482 328586 706718
rect 328822 706482 364586 706718
rect 364822 706482 400586 706718
rect 400822 706482 436586 706718
rect 436822 706482 472586 706718
rect 472822 706482 508586 706718
rect 508822 706482 544586 706718
rect 544822 706482 580586 706718
rect 580822 706482 587382 706718
rect 587618 706482 587800 706718
rect -3876 706398 587800 706482
rect -3876 706162 -3694 706398
rect -3458 706162 4586 706398
rect 4822 706162 40586 706398
rect 40822 706162 76586 706398
rect 76822 706162 112586 706398
rect 112822 706162 148586 706398
rect 148822 706162 184586 706398
rect 184822 706162 220586 706398
rect 220822 706162 256586 706398
rect 256822 706162 292586 706398
rect 292822 706162 328586 706398
rect 328822 706162 364586 706398
rect 364822 706162 400586 706398
rect 400822 706162 436586 706398
rect 436822 706162 472586 706398
rect 472822 706162 508586 706398
rect 508822 706162 544586 706398
rect 544822 706162 580586 706398
rect 580822 706162 587382 706398
rect 587618 706162 587800 706398
rect -3876 706140 587800 706162
rect -3876 706138 -3276 706140
rect 4404 706138 5004 706140
rect 40404 706138 41004 706140
rect 76404 706138 77004 706140
rect 112404 706138 113004 706140
rect 148404 706138 149004 706140
rect 184404 706138 185004 706140
rect 220404 706138 221004 706140
rect 256404 706138 257004 706140
rect 292404 706138 293004 706140
rect 328404 706138 329004 706140
rect 364404 706138 365004 706140
rect 400404 706138 401004 706140
rect 436404 706138 437004 706140
rect 472404 706138 473004 706140
rect 508404 706138 509004 706140
rect 544404 706138 545004 706140
rect 580404 706138 581004 706140
rect 587200 706138 587800 706140
rect -2936 705800 -2336 705802
rect 18804 705800 19404 705802
rect 54804 705800 55404 705802
rect 90804 705800 91404 705802
rect 126804 705800 127404 705802
rect 162804 705800 163404 705802
rect 198804 705800 199404 705802
rect 234804 705800 235404 705802
rect 270804 705800 271404 705802
rect 306804 705800 307404 705802
rect 342804 705800 343404 705802
rect 378804 705800 379404 705802
rect 414804 705800 415404 705802
rect 450804 705800 451404 705802
rect 486804 705800 487404 705802
rect 522804 705800 523404 705802
rect 558804 705800 559404 705802
rect 586260 705800 586860 705802
rect -2936 705778 586860 705800
rect -2936 705542 -2754 705778
rect -2518 705542 18986 705778
rect 19222 705542 54986 705778
rect 55222 705542 90986 705778
rect 91222 705542 126986 705778
rect 127222 705542 162986 705778
rect 163222 705542 198986 705778
rect 199222 705542 234986 705778
rect 235222 705542 270986 705778
rect 271222 705542 306986 705778
rect 307222 705542 342986 705778
rect 343222 705542 378986 705778
rect 379222 705542 414986 705778
rect 415222 705542 450986 705778
rect 451222 705542 486986 705778
rect 487222 705542 522986 705778
rect 523222 705542 558986 705778
rect 559222 705542 586442 705778
rect 586678 705542 586860 705778
rect -2936 705458 586860 705542
rect -2936 705222 -2754 705458
rect -2518 705222 18986 705458
rect 19222 705222 54986 705458
rect 55222 705222 90986 705458
rect 91222 705222 126986 705458
rect 127222 705222 162986 705458
rect 163222 705222 198986 705458
rect 199222 705222 234986 705458
rect 235222 705222 270986 705458
rect 271222 705222 306986 705458
rect 307222 705222 342986 705458
rect 343222 705222 378986 705458
rect 379222 705222 414986 705458
rect 415222 705222 450986 705458
rect 451222 705222 486986 705458
rect 487222 705222 522986 705458
rect 523222 705222 558986 705458
rect 559222 705222 586442 705458
rect 586678 705222 586860 705458
rect -2936 705200 586860 705222
rect -2936 705198 -2336 705200
rect 18804 705198 19404 705200
rect 54804 705198 55404 705200
rect 90804 705198 91404 705200
rect 126804 705198 127404 705200
rect 162804 705198 163404 705200
rect 198804 705198 199404 705200
rect 234804 705198 235404 705200
rect 270804 705198 271404 705200
rect 306804 705198 307404 705200
rect 342804 705198 343404 705200
rect 378804 705198 379404 705200
rect 414804 705198 415404 705200
rect 450804 705198 451404 705200
rect 486804 705198 487404 705200
rect 522804 705198 523404 705200
rect 558804 705198 559404 705200
rect 586260 705198 586860 705200
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -7636 697276 -7036 697278
rect 590960 697276 591560 697278
rect -8576 697254 592500 697276
rect -8576 697018 -7454 697254
rect -7218 697018 591142 697254
rect 591378 697018 592500 697254
rect -8576 696934 592500 697018
rect -8576 696698 -7454 696934
rect -7218 696698 591142 696934
rect 591378 696698 592500 696934
rect -8576 696676 592500 696698
rect -7636 696674 -7036 696676
rect 590960 696674 591560 696676
rect -5756 693676 -5156 693678
rect 589080 693676 589680 693678
rect -6696 693654 590620 693676
rect -6696 693418 -5574 693654
rect -5338 693418 589262 693654
rect 589498 693418 590620 693654
rect -6696 693334 590620 693418
rect -6696 693098 -5574 693334
rect -5338 693098 589262 693334
rect 589498 693098 590620 693334
rect -6696 693076 590620 693098
rect -5756 693074 -5156 693076
rect 589080 693074 589680 693076
rect 37100 692698 46988 692740
rect 37100 692462 37142 692698
rect 37378 692462 46710 692698
rect 46946 692462 46988 692698
rect 37100 692420 46988 692462
rect 56420 692698 66308 692740
rect 56420 692462 56462 692698
rect 56698 692462 66030 692698
rect 66266 692462 66308 692698
rect 56420 692420 66308 692462
rect 75740 692698 84524 692740
rect 75740 692462 75782 692698
rect 76018 692462 84246 692698
rect 84482 692462 84524 692698
rect 75740 692420 84524 692462
rect 108676 692698 114332 692740
rect 108676 692462 108718 692698
rect 108954 692462 114054 692698
rect 114290 692462 114332 692698
rect 108676 692420 114332 692462
rect 124132 692698 133652 692740
rect 124132 692462 124174 692698
rect 124410 692462 133374 692698
rect 133610 692462 133652 692698
rect 124132 692420 133652 692462
rect 143636 692698 152972 692740
rect 143636 692462 143678 692698
rect 143914 692462 152694 692698
rect 152930 692462 152972 692698
rect 143636 692420 152972 692462
rect 539420 692698 549308 692740
rect 539420 692462 539462 692698
rect 539698 692462 549030 692698
rect 549266 692462 549308 692698
rect 539420 692420 549308 692462
rect 558740 692698 565868 692740
rect 558740 692462 558782 692698
rect 559018 692462 565590 692698
rect 565826 692462 565868 692698
rect 558740 692420 565868 692462
rect -3876 690076 -3276 690078
rect 4404 690076 5004 690078
rect 580404 690076 581004 690078
rect 587200 690076 587800 690078
rect -4816 690054 588740 690076
rect -4816 689818 -3694 690054
rect -3458 689818 4586 690054
rect 4822 689818 580586 690054
rect 580822 689818 587382 690054
rect 587618 689818 588740 690054
rect -4816 689734 588740 689818
rect -4816 689498 -3694 689734
rect -3458 689498 4586 689734
rect 4822 689498 580586 689734
rect 580822 689498 587382 689734
rect 587618 689498 588740 689734
rect -4816 689476 588740 689498
rect -3876 689474 -3276 689476
rect 4404 689474 5004 689476
rect 580404 689474 581004 689476
rect 587200 689474 587800 689476
rect -1996 686428 -1396 686430
rect 804 686428 1404 686430
rect 585320 686428 585920 686430
rect -2936 686406 586860 686428
rect -2936 686170 -1814 686406
rect -1578 686170 986 686406
rect 1222 686170 585502 686406
rect 585738 686170 586860 686406
rect -2936 686086 586860 686170
rect -2936 685850 -1814 686086
rect -1578 685850 986 686086
rect 1222 685850 585502 686086
rect 585738 685850 586860 686086
rect -2936 685828 586860 685850
rect -1996 685826 -1396 685828
rect 804 685826 1404 685828
rect 585320 685826 585920 685828
rect -8576 679276 -7976 679278
rect 591900 679276 592500 679278
rect -8576 679254 592500 679276
rect -8576 679018 -8394 679254
rect -8158 679018 592082 679254
rect 592318 679018 592500 679254
rect -8576 678934 592500 679018
rect -8576 678698 -8394 678934
rect -8158 678698 592082 678934
rect 592318 678698 592500 678934
rect -8576 678676 592500 678698
rect -8576 678674 -7976 678676
rect 591900 678674 592500 678676
rect -6696 675676 -6096 675678
rect 590020 675676 590620 675678
rect -6696 675654 590620 675676
rect -6696 675418 -6514 675654
rect -6278 675418 590202 675654
rect 590438 675418 590620 675654
rect -6696 675334 590620 675418
rect -6696 675098 -6514 675334
rect -6278 675098 590202 675334
rect 590438 675098 590620 675334
rect -6696 675076 590620 675098
rect -6696 675074 -6096 675076
rect 590020 675074 590620 675076
rect -4816 672076 -4216 672078
rect 588140 672076 588740 672078
rect -4816 672054 588740 672076
rect -4816 671818 -4634 672054
rect -4398 671818 588322 672054
rect 588558 671818 588740 672054
rect -4816 671734 588740 671818
rect -4816 671498 -4634 671734
rect -4398 671498 588322 671734
rect 588558 671498 588740 671734
rect -4816 671476 588740 671498
rect -4816 671474 -4216 671476
rect 588140 671474 588740 671476
rect -2936 668428 -2336 668430
rect 586260 668428 586860 668430
rect -2936 668406 586860 668428
rect -2936 668170 -2754 668406
rect -2518 668170 586442 668406
rect 586678 668170 586860 668406
rect -2936 668086 586860 668170
rect -2936 667850 -2754 668086
rect -2518 667850 586442 668086
rect 586678 667850 586860 668086
rect -2936 667828 586860 667850
rect -2936 667826 -2336 667828
rect 586260 667826 586860 667828
rect -7636 661276 -7036 661278
rect 590960 661276 591560 661278
rect -8576 661254 592500 661276
rect -8576 661018 -7454 661254
rect -7218 661018 591142 661254
rect 591378 661018 592500 661254
rect -8576 660934 592500 661018
rect -8576 660698 -7454 660934
rect -7218 660698 591142 660934
rect 591378 660698 592500 660934
rect -8576 660676 592500 660698
rect -7636 660674 -7036 660676
rect 590960 660674 591560 660676
rect -5756 657676 -5156 657678
rect 589080 657676 589680 657678
rect -6696 657654 590620 657676
rect -6696 657418 -5574 657654
rect -5338 657418 589262 657654
rect 589498 657418 590620 657654
rect -6696 657334 590620 657418
rect -6696 657098 -5574 657334
rect -5338 657098 589262 657334
rect 589498 657098 590620 657334
rect -6696 657076 590620 657098
rect -5756 657074 -5156 657076
rect 589080 657074 589680 657076
rect -3876 654076 -3276 654078
rect 4404 654076 5004 654078
rect 580404 654076 581004 654078
rect 587200 654076 587800 654078
rect -4816 654054 588740 654076
rect -4816 653818 -3694 654054
rect -3458 653818 4586 654054
rect 4822 653818 580586 654054
rect 580822 653818 587382 654054
rect 587618 653818 588740 654054
rect -4816 653734 588740 653818
rect -4816 653498 -3694 653734
rect -3458 653498 4586 653734
rect 4822 653498 580586 653734
rect 580822 653498 587382 653734
rect 587618 653498 588740 653734
rect -4816 653476 588740 653498
rect -3876 653474 -3276 653476
rect 4404 653474 5004 653476
rect 580404 653474 581004 653476
rect 587200 653474 587800 653476
rect -1996 650428 -1396 650430
rect 804 650428 1404 650430
rect 585320 650428 585920 650430
rect -2936 650406 586860 650428
rect -2936 650170 -1814 650406
rect -1578 650170 986 650406
rect 1222 650170 585502 650406
rect 585738 650170 586860 650406
rect -2936 650086 586860 650170
rect -2936 649850 -1814 650086
rect -1578 649850 986 650086
rect 1222 649850 585502 650086
rect 585738 649850 586860 650086
rect -2936 649828 586860 649850
rect -1996 649826 -1396 649828
rect 804 649826 1404 649828
rect 585320 649826 585920 649828
rect -8576 643276 -7976 643278
rect 591900 643276 592500 643278
rect -8576 643254 592500 643276
rect -8576 643018 -8394 643254
rect -8158 643018 592082 643254
rect 592318 643018 592500 643254
rect -8576 642934 592500 643018
rect -8576 642698 -8394 642934
rect -8158 642698 592082 642934
rect 592318 642698 592500 642934
rect -8576 642676 592500 642698
rect -8576 642674 -7976 642676
rect 591900 642674 592500 642676
rect -6696 639676 -6096 639678
rect 590020 639676 590620 639678
rect -6696 639654 590620 639676
rect -6696 639418 -6514 639654
rect -6278 639418 590202 639654
rect 590438 639418 590620 639654
rect -6696 639334 590620 639418
rect -6696 639098 -6514 639334
rect -6278 639098 590202 639334
rect 590438 639098 590620 639334
rect -6696 639076 590620 639098
rect -6696 639074 -6096 639076
rect 590020 639074 590620 639076
rect -4816 636076 -4216 636078
rect 588140 636076 588740 636078
rect -4816 636054 588740 636076
rect -4816 635818 -4634 636054
rect -4398 635818 588322 636054
rect 588558 635818 588740 636054
rect -4816 635734 588740 635818
rect -4816 635498 -4634 635734
rect -4398 635498 588322 635734
rect 588558 635498 588740 635734
rect -4816 635476 588740 635498
rect -4816 635474 -4216 635476
rect 588140 635474 588740 635476
rect -2936 632428 -2336 632430
rect 586260 632428 586860 632430
rect -2936 632406 586860 632428
rect -2936 632170 -2754 632406
rect -2518 632170 586442 632406
rect 586678 632170 586860 632406
rect -2936 632086 586860 632170
rect -2936 631850 -2754 632086
rect -2518 631850 586442 632086
rect 586678 631850 586860 632086
rect -2936 631828 586860 631850
rect -2936 631826 -2336 631828
rect 586260 631826 586860 631828
rect -7636 625276 -7036 625278
rect 590960 625276 591560 625278
rect -8576 625254 592500 625276
rect -8576 625018 -7454 625254
rect -7218 625018 591142 625254
rect 591378 625018 592500 625254
rect -8576 624934 592500 625018
rect -8576 624698 -7454 624934
rect -7218 624698 591142 624934
rect 591378 624698 592500 624934
rect -8576 624676 592500 624698
rect -7636 624674 -7036 624676
rect 590960 624674 591560 624676
rect -5756 621676 -5156 621678
rect 589080 621676 589680 621678
rect -6696 621654 590620 621676
rect -6696 621418 -5574 621654
rect -5338 621418 589262 621654
rect 589498 621418 590620 621654
rect -6696 621334 590620 621418
rect -6696 621098 -5574 621334
rect -5338 621098 589262 621334
rect 589498 621098 590620 621334
rect -6696 621076 590620 621098
rect -5756 621074 -5156 621076
rect 589080 621074 589680 621076
rect -3876 618076 -3276 618078
rect 4404 618076 5004 618078
rect 580404 618076 581004 618078
rect 587200 618076 587800 618078
rect -4816 618054 588740 618076
rect -4816 617818 -3694 618054
rect -3458 617818 4586 618054
rect 4822 617818 580586 618054
rect 580822 617818 587382 618054
rect 587618 617818 588740 618054
rect -4816 617734 588740 617818
rect -4816 617498 -3694 617734
rect -3458 617498 4586 617734
rect 4822 617498 580586 617734
rect 580822 617498 587382 617734
rect 587618 617498 588740 617734
rect -4816 617476 588740 617498
rect -3876 617474 -3276 617476
rect 4404 617474 5004 617476
rect 580404 617474 581004 617476
rect 587200 617474 587800 617476
rect -1996 614428 -1396 614430
rect 804 614428 1404 614430
rect 585320 614428 585920 614430
rect -2936 614406 586860 614428
rect -2936 614170 -1814 614406
rect -1578 614170 986 614406
rect 1222 614170 585502 614406
rect 585738 614170 586860 614406
rect -2936 614086 586860 614170
rect -2936 613850 -1814 614086
rect -1578 613850 986 614086
rect 1222 613850 585502 614086
rect 585738 613850 586860 614086
rect -2936 613828 586860 613850
rect -1996 613826 -1396 613828
rect 804 613826 1404 613828
rect 585320 613826 585920 613828
rect -8576 607276 -7976 607278
rect 591900 607276 592500 607278
rect -8576 607254 592500 607276
rect -8576 607018 -8394 607254
rect -8158 607018 592082 607254
rect 592318 607018 592500 607254
rect -8576 606934 592500 607018
rect -8576 606698 -8394 606934
rect -8158 606698 592082 606934
rect 592318 606698 592500 606934
rect -8576 606676 592500 606698
rect -8576 606674 -7976 606676
rect 591900 606674 592500 606676
rect -6696 603676 -6096 603678
rect 590020 603676 590620 603678
rect -6696 603654 590620 603676
rect -6696 603418 -6514 603654
rect -6278 603418 590202 603654
rect 590438 603418 590620 603654
rect -6696 603334 590620 603418
rect -6696 603098 -6514 603334
rect -6278 603098 590202 603334
rect 590438 603098 590620 603334
rect -6696 603076 590620 603098
rect -6696 603074 -6096 603076
rect 590020 603074 590620 603076
rect -4816 600076 -4216 600078
rect 588140 600076 588740 600078
rect -4816 600054 588740 600076
rect -4816 599818 -4634 600054
rect -4398 599818 588322 600054
rect 588558 599818 588740 600054
rect -4816 599734 588740 599818
rect -4816 599498 -4634 599734
rect -4398 599498 588322 599734
rect 588558 599498 588740 599734
rect -4816 599476 588740 599498
rect -4816 599474 -4216 599476
rect 588140 599474 588740 599476
rect -2936 596428 -2336 596430
rect 586260 596428 586860 596430
rect -2936 596406 586860 596428
rect -2936 596170 -2754 596406
rect -2518 596170 586442 596406
rect 586678 596170 586860 596406
rect -2936 596086 586860 596170
rect -2936 595850 -2754 596086
rect -2518 595850 586442 596086
rect 586678 595850 586860 596086
rect -2936 595828 586860 595850
rect -2936 595826 -2336 595828
rect 586260 595826 586860 595828
rect -7636 589276 -7036 589278
rect 590960 589276 591560 589278
rect -8576 589254 592500 589276
rect -8576 589018 -7454 589254
rect -7218 589018 591142 589254
rect 591378 589018 592500 589254
rect -8576 588934 592500 589018
rect -8576 588698 -7454 588934
rect -7218 588698 591142 588934
rect 591378 588698 592500 588934
rect -8576 588676 592500 588698
rect -7636 588674 -7036 588676
rect 590960 588674 591560 588676
rect -5756 585676 -5156 585678
rect 589080 585676 589680 585678
rect -6696 585654 590620 585676
rect -6696 585418 -5574 585654
rect -5338 585418 589262 585654
rect 589498 585418 590620 585654
rect -6696 585334 590620 585418
rect -6696 585098 -5574 585334
rect -5338 585098 589262 585334
rect 589498 585098 590620 585334
rect -6696 585076 590620 585098
rect -5756 585074 -5156 585076
rect 589080 585074 589680 585076
rect -3876 582076 -3276 582078
rect 4404 582076 5004 582078
rect 580404 582076 581004 582078
rect 587200 582076 587800 582078
rect -4816 582054 588740 582076
rect -4816 581818 -3694 582054
rect -3458 581818 4586 582054
rect 4822 581818 580586 582054
rect 580822 581818 587382 582054
rect 587618 581818 588740 582054
rect -4816 581734 588740 581818
rect -4816 581498 -3694 581734
rect -3458 581498 4586 581734
rect 4822 581498 580586 581734
rect 580822 581498 587382 581734
rect 587618 581498 588740 581734
rect -4816 581476 588740 581498
rect -3876 581474 -3276 581476
rect 4404 581474 5004 581476
rect 580404 581474 581004 581476
rect 587200 581474 587800 581476
rect -1996 578428 -1396 578430
rect 804 578428 1404 578430
rect 585320 578428 585920 578430
rect -2936 578406 586860 578428
rect -2936 578170 -1814 578406
rect -1578 578170 986 578406
rect 1222 578170 585502 578406
rect 585738 578170 586860 578406
rect -2936 578086 586860 578170
rect -2936 577850 -1814 578086
rect -1578 577850 986 578086
rect 1222 577850 585502 578086
rect 585738 577850 586860 578086
rect -2936 577828 586860 577850
rect -1996 577826 -1396 577828
rect 804 577826 1404 577828
rect 585320 577826 585920 577828
rect -8576 571276 -7976 571278
rect 591900 571276 592500 571278
rect -8576 571254 592500 571276
rect -8576 571018 -8394 571254
rect -8158 571018 592082 571254
rect 592318 571018 592500 571254
rect -8576 570934 592500 571018
rect -8576 570698 -8394 570934
rect -8158 570698 592082 570934
rect 592318 570698 592500 570934
rect -8576 570676 592500 570698
rect -8576 570674 -7976 570676
rect 591900 570674 592500 570676
rect -6696 567676 -6096 567678
rect 590020 567676 590620 567678
rect -6696 567654 590620 567676
rect -6696 567418 -6514 567654
rect -6278 567418 590202 567654
rect 590438 567418 590620 567654
rect -6696 567334 590620 567418
rect -6696 567098 -6514 567334
rect -6278 567098 590202 567334
rect 590438 567098 590620 567334
rect -6696 567076 590620 567098
rect -6696 567074 -6096 567076
rect 590020 567074 590620 567076
rect -4816 564076 -4216 564078
rect 588140 564076 588740 564078
rect -4816 564054 588740 564076
rect -4816 563818 -4634 564054
rect -4398 563818 588322 564054
rect 588558 563818 588740 564054
rect -4816 563734 588740 563818
rect -4816 563498 -4634 563734
rect -4398 563498 588322 563734
rect 588558 563498 588740 563734
rect -4816 563476 588740 563498
rect -4816 563474 -4216 563476
rect 588140 563474 588740 563476
rect -2936 560428 -2336 560430
rect 586260 560428 586860 560430
rect -2936 560406 586860 560428
rect -2936 560170 -2754 560406
rect -2518 560170 586442 560406
rect 586678 560170 586860 560406
rect -2936 560086 586860 560170
rect -2936 559850 -2754 560086
rect -2518 559850 586442 560086
rect 586678 559850 586860 560086
rect -2936 559828 586860 559850
rect -2936 559826 -2336 559828
rect 586260 559826 586860 559828
rect -7636 553276 -7036 553278
rect 590960 553276 591560 553278
rect -8576 553254 592500 553276
rect -8576 553018 -7454 553254
rect -7218 553018 591142 553254
rect 591378 553018 592500 553254
rect -8576 552934 592500 553018
rect -8576 552698 -7454 552934
rect -7218 552698 591142 552934
rect 591378 552698 592500 552934
rect -8576 552676 592500 552698
rect -7636 552674 -7036 552676
rect 590960 552674 591560 552676
rect -5756 549676 -5156 549678
rect 589080 549676 589680 549678
rect -6696 549654 590620 549676
rect -6696 549418 -5574 549654
rect -5338 549418 589262 549654
rect 589498 549418 590620 549654
rect -6696 549334 590620 549418
rect -6696 549098 -5574 549334
rect -5338 549098 589262 549334
rect 589498 549098 590620 549334
rect -6696 549076 590620 549098
rect -5756 549074 -5156 549076
rect 589080 549074 589680 549076
rect -3876 546076 -3276 546078
rect 4404 546076 5004 546078
rect 580404 546076 581004 546078
rect 587200 546076 587800 546078
rect -4816 546054 588740 546076
rect -4816 545818 -3694 546054
rect -3458 545818 4586 546054
rect 4822 545818 580586 546054
rect 580822 545818 587382 546054
rect 587618 545818 588740 546054
rect -4816 545734 588740 545818
rect -4816 545498 -3694 545734
rect -3458 545498 4586 545734
rect 4822 545498 580586 545734
rect 580822 545498 587382 545734
rect 587618 545498 588740 545734
rect -4816 545476 588740 545498
rect -3876 545474 -3276 545476
rect 4404 545474 5004 545476
rect 580404 545474 581004 545476
rect 587200 545474 587800 545476
rect -1996 542428 -1396 542430
rect 804 542428 1404 542430
rect 585320 542428 585920 542430
rect -2936 542406 586860 542428
rect -2936 542170 -1814 542406
rect -1578 542170 986 542406
rect 1222 542170 585502 542406
rect 585738 542170 586860 542406
rect -2936 542086 586860 542170
rect -2936 541850 -1814 542086
rect -1578 541850 986 542086
rect 1222 541850 585502 542086
rect 585738 541850 586860 542086
rect -2936 541828 586860 541850
rect -1996 541826 -1396 541828
rect 804 541826 1404 541828
rect 585320 541826 585920 541828
rect -8576 535276 -7976 535278
rect 591900 535276 592500 535278
rect -8576 535254 592500 535276
rect -8576 535018 -8394 535254
rect -8158 535018 592082 535254
rect 592318 535018 592500 535254
rect -8576 534934 592500 535018
rect -8576 534698 -8394 534934
rect -8158 534698 592082 534934
rect 592318 534698 592500 534934
rect -8576 534676 592500 534698
rect -8576 534674 -7976 534676
rect 591900 534674 592500 534676
rect -6696 531676 -6096 531678
rect 590020 531676 590620 531678
rect -6696 531654 590620 531676
rect -6696 531418 -6514 531654
rect -6278 531418 590202 531654
rect 590438 531418 590620 531654
rect -6696 531334 590620 531418
rect -6696 531098 -6514 531334
rect -6278 531098 590202 531334
rect 590438 531098 590620 531334
rect -6696 531076 590620 531098
rect -6696 531074 -6096 531076
rect 590020 531074 590620 531076
rect -4816 528076 -4216 528078
rect 588140 528076 588740 528078
rect -4816 528054 588740 528076
rect -4816 527818 -4634 528054
rect -4398 527818 588322 528054
rect 588558 527818 588740 528054
rect -4816 527734 588740 527818
rect -4816 527498 -4634 527734
rect -4398 527498 588322 527734
rect 588558 527498 588740 527734
rect -4816 527476 588740 527498
rect -4816 527474 -4216 527476
rect 588140 527474 588740 527476
rect -2936 524428 -2336 524430
rect 586260 524428 586860 524430
rect -2936 524406 586860 524428
rect -2936 524170 -2754 524406
rect -2518 524170 586442 524406
rect 586678 524170 586860 524406
rect -2936 524086 586860 524170
rect -2936 523850 -2754 524086
rect -2518 523850 586442 524086
rect 586678 523850 586860 524086
rect -2936 523828 586860 523850
rect -2936 523826 -2336 523828
rect 586260 523826 586860 523828
rect -7636 517276 -7036 517278
rect 590960 517276 591560 517278
rect -8576 517254 592500 517276
rect -8576 517018 -7454 517254
rect -7218 517018 591142 517254
rect 591378 517018 592500 517254
rect -8576 516934 592500 517018
rect -8576 516698 -7454 516934
rect -7218 516698 591142 516934
rect 591378 516698 592500 516934
rect -8576 516676 592500 516698
rect -7636 516674 -7036 516676
rect 590960 516674 591560 516676
rect -5756 513676 -5156 513678
rect 589080 513676 589680 513678
rect -6696 513654 590620 513676
rect -6696 513418 -5574 513654
rect -5338 513418 589262 513654
rect 589498 513418 590620 513654
rect -6696 513334 590620 513418
rect -6696 513098 -5574 513334
rect -5338 513098 589262 513334
rect 589498 513098 590620 513334
rect -6696 513076 590620 513098
rect -5756 513074 -5156 513076
rect 589080 513074 589680 513076
rect -3876 510076 -3276 510078
rect 4404 510076 5004 510078
rect 580404 510076 581004 510078
rect 587200 510076 587800 510078
rect -4816 510054 588740 510076
rect -4816 509818 -3694 510054
rect -3458 509818 4586 510054
rect 4822 509818 580586 510054
rect 580822 509818 587382 510054
rect 587618 509818 588740 510054
rect -4816 509734 588740 509818
rect -4816 509498 -3694 509734
rect -3458 509498 4586 509734
rect 4822 509498 580586 509734
rect 580822 509498 587382 509734
rect 587618 509498 588740 509734
rect -4816 509476 588740 509498
rect -3876 509474 -3276 509476
rect 4404 509474 5004 509476
rect 580404 509474 581004 509476
rect 587200 509474 587800 509476
rect -1996 506428 -1396 506430
rect 804 506428 1404 506430
rect 585320 506428 585920 506430
rect -2936 506406 586860 506428
rect -2936 506170 -1814 506406
rect -1578 506170 986 506406
rect 1222 506170 585502 506406
rect 585738 506170 586860 506406
rect -2936 506086 586860 506170
rect -2936 505850 -1814 506086
rect -1578 505850 986 506086
rect 1222 505850 585502 506086
rect 585738 505850 586860 506086
rect -2936 505828 586860 505850
rect -1996 505826 -1396 505828
rect 804 505826 1404 505828
rect 585320 505826 585920 505828
rect -8576 499276 -7976 499278
rect 591900 499276 592500 499278
rect -8576 499254 592500 499276
rect -8576 499018 -8394 499254
rect -8158 499018 592082 499254
rect 592318 499018 592500 499254
rect -8576 498934 592500 499018
rect -8576 498698 -8394 498934
rect -8158 498698 592082 498934
rect 592318 498698 592500 498934
rect -8576 498676 592500 498698
rect -8576 498674 -7976 498676
rect 591900 498674 592500 498676
rect -6696 495676 -6096 495678
rect 590020 495676 590620 495678
rect -6696 495654 590620 495676
rect -6696 495418 -6514 495654
rect -6278 495418 590202 495654
rect 590438 495418 590620 495654
rect -6696 495334 590620 495418
rect -6696 495098 -6514 495334
rect -6278 495098 590202 495334
rect 590438 495098 590620 495334
rect -6696 495076 590620 495098
rect -6696 495074 -6096 495076
rect 590020 495074 590620 495076
rect -4816 492076 -4216 492078
rect 588140 492076 588740 492078
rect -4816 492054 588740 492076
rect -4816 491818 -4634 492054
rect -4398 491818 588322 492054
rect 588558 491818 588740 492054
rect -4816 491734 588740 491818
rect -4816 491498 -4634 491734
rect -4398 491498 588322 491734
rect 588558 491498 588740 491734
rect -4816 491476 588740 491498
rect -4816 491474 -4216 491476
rect 588140 491474 588740 491476
rect -2936 488428 -2336 488430
rect 586260 488428 586860 488430
rect -2936 488406 586860 488428
rect -2936 488170 -2754 488406
rect -2518 488170 586442 488406
rect 586678 488170 586860 488406
rect -2936 488086 586860 488170
rect -2936 487850 -2754 488086
rect -2518 487850 586442 488086
rect 586678 487850 586860 488086
rect -2936 487828 586860 487850
rect -2936 487826 -2336 487828
rect 586260 487826 586860 487828
rect -7636 481276 -7036 481278
rect 590960 481276 591560 481278
rect -8576 481254 592500 481276
rect -8576 481018 -7454 481254
rect -7218 481018 591142 481254
rect 591378 481018 592500 481254
rect -8576 480934 592500 481018
rect -8576 480698 -7454 480934
rect -7218 480698 591142 480934
rect 591378 480698 592500 480934
rect -8576 480676 592500 480698
rect -7636 480674 -7036 480676
rect 590960 480674 591560 480676
rect -5756 477676 -5156 477678
rect 589080 477676 589680 477678
rect -6696 477654 590620 477676
rect -6696 477418 -5574 477654
rect -5338 477418 589262 477654
rect 589498 477418 590620 477654
rect -6696 477334 590620 477418
rect -6696 477098 -5574 477334
rect -5338 477098 589262 477334
rect 589498 477098 590620 477334
rect -6696 477076 590620 477098
rect -5756 477074 -5156 477076
rect 589080 477074 589680 477076
rect -3876 474076 -3276 474078
rect 4404 474076 5004 474078
rect 580404 474076 581004 474078
rect 587200 474076 587800 474078
rect -4816 474054 588740 474076
rect -4816 473818 -3694 474054
rect -3458 473818 4586 474054
rect 4822 473818 580586 474054
rect 580822 473818 587382 474054
rect 587618 473818 588740 474054
rect -4816 473734 588740 473818
rect -4816 473498 -3694 473734
rect -3458 473498 4586 473734
rect 4822 473498 580586 473734
rect 580822 473498 587382 473734
rect 587618 473498 588740 473734
rect -4816 473476 588740 473498
rect -3876 473474 -3276 473476
rect 4404 473474 5004 473476
rect 580404 473474 581004 473476
rect 587200 473474 587800 473476
rect -1996 470428 -1396 470430
rect 804 470428 1404 470430
rect 585320 470428 585920 470430
rect -2936 470406 586860 470428
rect -2936 470170 -1814 470406
rect -1578 470170 986 470406
rect 1222 470170 585502 470406
rect 585738 470170 586860 470406
rect -2936 470086 586860 470170
rect -2936 469850 -1814 470086
rect -1578 469850 986 470086
rect 1222 469850 585502 470086
rect 585738 469850 586860 470086
rect -2936 469828 586860 469850
rect -1996 469826 -1396 469828
rect 804 469826 1404 469828
rect 585320 469826 585920 469828
rect -8576 463276 -7976 463278
rect 591900 463276 592500 463278
rect -8576 463254 592500 463276
rect -8576 463018 -8394 463254
rect -8158 463018 592082 463254
rect 592318 463018 592500 463254
rect -8576 462934 592500 463018
rect -8576 462698 -8394 462934
rect -8158 462698 592082 462934
rect 592318 462698 592500 462934
rect -8576 462676 592500 462698
rect -8576 462674 -7976 462676
rect 591900 462674 592500 462676
rect -6696 459676 -6096 459678
rect 590020 459676 590620 459678
rect -6696 459654 590620 459676
rect -6696 459418 -6514 459654
rect -6278 459418 590202 459654
rect 590438 459418 590620 459654
rect -6696 459334 590620 459418
rect -6696 459098 -6514 459334
rect -6278 459098 590202 459334
rect 590438 459098 590620 459334
rect -6696 459076 590620 459098
rect -6696 459074 -6096 459076
rect 590020 459074 590620 459076
rect -4816 456076 -4216 456078
rect 588140 456076 588740 456078
rect -4816 456054 588740 456076
rect -4816 455818 -4634 456054
rect -4398 455818 588322 456054
rect 588558 455818 588740 456054
rect -4816 455734 588740 455818
rect -4816 455498 -4634 455734
rect -4398 455498 588322 455734
rect 588558 455498 588740 455734
rect -4816 455476 588740 455498
rect -4816 455474 -4216 455476
rect 588140 455474 588740 455476
rect -2936 452428 -2336 452430
rect 586260 452428 586860 452430
rect -2936 452406 586860 452428
rect -2936 452170 -2754 452406
rect -2518 452170 586442 452406
rect 586678 452170 586860 452406
rect -2936 452086 586860 452170
rect -2936 451850 -2754 452086
rect -2518 451850 586442 452086
rect 586678 451850 586860 452086
rect -2936 451828 586860 451850
rect -2936 451826 -2336 451828
rect 586260 451826 586860 451828
rect -7636 445276 -7036 445278
rect 590960 445276 591560 445278
rect -8576 445254 592500 445276
rect -8576 445018 -7454 445254
rect -7218 445018 591142 445254
rect 591378 445018 592500 445254
rect -8576 444934 592500 445018
rect -8576 444698 -7454 444934
rect -7218 444698 591142 444934
rect 591378 444698 592500 444934
rect -8576 444676 592500 444698
rect -7636 444674 -7036 444676
rect 590960 444674 591560 444676
rect -5756 441676 -5156 441678
rect 589080 441676 589680 441678
rect -6696 441654 590620 441676
rect -6696 441418 -5574 441654
rect -5338 441418 589262 441654
rect 589498 441418 590620 441654
rect -6696 441334 590620 441418
rect -6696 441098 -5574 441334
rect -5338 441098 589262 441334
rect 589498 441098 590620 441334
rect -6696 441076 590620 441098
rect -5756 441074 -5156 441076
rect 589080 441074 589680 441076
rect -3876 438076 -3276 438078
rect 4404 438076 5004 438078
rect 580404 438076 581004 438078
rect 587200 438076 587800 438078
rect -4816 438054 588740 438076
rect -4816 437818 -3694 438054
rect -3458 437818 4586 438054
rect 4822 437818 580586 438054
rect 580822 437818 587382 438054
rect 587618 437818 588740 438054
rect -4816 437734 588740 437818
rect -4816 437498 -3694 437734
rect -3458 437498 4586 437734
rect 4822 437498 580586 437734
rect 580822 437498 587382 437734
rect 587618 437498 588740 437734
rect -4816 437476 588740 437498
rect -3876 437474 -3276 437476
rect 4404 437474 5004 437476
rect 580404 437474 581004 437476
rect 587200 437474 587800 437476
rect -1996 434428 -1396 434430
rect 804 434428 1404 434430
rect 585320 434428 585920 434430
rect -2936 434406 586860 434428
rect -2936 434170 -1814 434406
rect -1578 434170 986 434406
rect 1222 434170 585502 434406
rect 585738 434170 586860 434406
rect -2936 434086 586860 434170
rect -2936 433850 -1814 434086
rect -1578 433850 986 434086
rect 1222 433850 585502 434086
rect 585738 433850 586860 434086
rect -2936 433828 586860 433850
rect -1996 433826 -1396 433828
rect 804 433826 1404 433828
rect 585320 433826 585920 433828
rect -8576 427276 -7976 427278
rect 591900 427276 592500 427278
rect -8576 427254 592500 427276
rect -8576 427018 -8394 427254
rect -8158 427018 592082 427254
rect 592318 427018 592500 427254
rect -8576 426934 592500 427018
rect -8576 426698 -8394 426934
rect -8158 426698 592082 426934
rect 592318 426698 592500 426934
rect -8576 426676 592500 426698
rect -8576 426674 -7976 426676
rect 591900 426674 592500 426676
rect -6696 423676 -6096 423678
rect 590020 423676 590620 423678
rect -6696 423654 590620 423676
rect -6696 423418 -6514 423654
rect -6278 423418 590202 423654
rect 590438 423418 590620 423654
rect -6696 423334 590620 423418
rect -6696 423098 -6514 423334
rect -6278 423098 590202 423334
rect 590438 423098 590620 423334
rect -6696 423076 590620 423098
rect -6696 423074 -6096 423076
rect 590020 423074 590620 423076
rect -4816 420076 -4216 420078
rect 588140 420076 588740 420078
rect -4816 420054 588740 420076
rect -4816 419818 -4634 420054
rect -4398 419818 588322 420054
rect 588558 419818 588740 420054
rect -4816 419734 588740 419818
rect -4816 419498 -4634 419734
rect -4398 419498 588322 419734
rect 588558 419498 588740 419734
rect -4816 419476 588740 419498
rect -4816 419474 -4216 419476
rect 588140 419474 588740 419476
rect -2936 416428 -2336 416430
rect 586260 416428 586860 416430
rect -2936 416406 586860 416428
rect -2936 416170 -2754 416406
rect -2518 416170 586442 416406
rect 586678 416170 586860 416406
rect -2936 416086 586860 416170
rect -2936 415850 -2754 416086
rect -2518 415850 586442 416086
rect 586678 415850 586860 416086
rect -2936 415828 586860 415850
rect -2936 415826 -2336 415828
rect 586260 415826 586860 415828
rect -7636 409276 -7036 409278
rect 590960 409276 591560 409278
rect -8576 409254 592500 409276
rect -8576 409018 -7454 409254
rect -7218 409018 591142 409254
rect 591378 409018 592500 409254
rect -8576 408934 592500 409018
rect -8576 408698 -7454 408934
rect -7218 408698 591142 408934
rect 591378 408698 592500 408934
rect -8576 408676 592500 408698
rect -7636 408674 -7036 408676
rect 590960 408674 591560 408676
rect -5756 405676 -5156 405678
rect 589080 405676 589680 405678
rect -6696 405654 590620 405676
rect -6696 405418 -5574 405654
rect -5338 405418 589262 405654
rect 589498 405418 590620 405654
rect -6696 405334 590620 405418
rect -6696 405098 -5574 405334
rect -5338 405098 589262 405334
rect 589498 405098 590620 405334
rect -6696 405076 590620 405098
rect -5756 405074 -5156 405076
rect 589080 405074 589680 405076
rect -3876 402076 -3276 402078
rect 4404 402076 5004 402078
rect 580404 402076 581004 402078
rect 587200 402076 587800 402078
rect -4816 402054 588740 402076
rect -4816 401818 -3694 402054
rect -3458 401818 4586 402054
rect 4822 401818 580586 402054
rect 580822 401818 587382 402054
rect 587618 401818 588740 402054
rect -4816 401734 588740 401818
rect -4816 401498 -3694 401734
rect -3458 401498 4586 401734
rect 4822 401498 580586 401734
rect 580822 401498 587382 401734
rect 587618 401498 588740 401734
rect -4816 401476 588740 401498
rect -3876 401474 -3276 401476
rect 4404 401474 5004 401476
rect 580404 401474 581004 401476
rect 587200 401474 587800 401476
rect -1996 398428 -1396 398430
rect 804 398428 1404 398430
rect 585320 398428 585920 398430
rect -2936 398406 586860 398428
rect -2936 398170 -1814 398406
rect -1578 398170 986 398406
rect 1222 398170 585502 398406
rect 585738 398170 586860 398406
rect -2936 398086 586860 398170
rect -2936 397850 -1814 398086
rect -1578 397850 986 398086
rect 1222 397850 585502 398086
rect 585738 397850 586860 398086
rect -2936 397828 586860 397850
rect -1996 397826 -1396 397828
rect 804 397826 1404 397828
rect 585320 397826 585920 397828
rect -8576 391276 -7976 391278
rect 591900 391276 592500 391278
rect -8576 391254 592500 391276
rect -8576 391018 -8394 391254
rect -8158 391018 592082 391254
rect 592318 391018 592500 391254
rect -8576 390934 592500 391018
rect -8576 390698 -8394 390934
rect -8158 390698 592082 390934
rect 592318 390698 592500 390934
rect -8576 390676 592500 390698
rect -8576 390674 -7976 390676
rect 591900 390674 592500 390676
rect -6696 387676 -6096 387678
rect 590020 387676 590620 387678
rect -6696 387654 590620 387676
rect -6696 387418 -6514 387654
rect -6278 387418 590202 387654
rect 590438 387418 590620 387654
rect -6696 387334 590620 387418
rect -6696 387098 -6514 387334
rect -6278 387098 590202 387334
rect 590438 387098 590620 387334
rect -6696 387076 590620 387098
rect -6696 387074 -6096 387076
rect 590020 387074 590620 387076
rect -4816 384076 -4216 384078
rect 588140 384076 588740 384078
rect -4816 384054 588740 384076
rect -4816 383818 -4634 384054
rect -4398 383818 588322 384054
rect 588558 383818 588740 384054
rect -4816 383734 588740 383818
rect -4816 383498 -4634 383734
rect -4398 383498 588322 383734
rect 588558 383498 588740 383734
rect -4816 383476 588740 383498
rect -4816 383474 -4216 383476
rect 588140 383474 588740 383476
rect -2936 380428 -2336 380430
rect 586260 380428 586860 380430
rect -2936 380406 586860 380428
rect -2936 380170 -2754 380406
rect -2518 380170 586442 380406
rect 586678 380170 586860 380406
rect -2936 380086 586860 380170
rect -2936 379850 -2754 380086
rect -2518 379850 586442 380086
rect 586678 379850 586860 380086
rect -2936 379828 586860 379850
rect -2936 379826 -2336 379828
rect 586260 379826 586860 379828
rect -7636 373276 -7036 373278
rect 590960 373276 591560 373278
rect -8576 373254 592500 373276
rect -8576 373018 -7454 373254
rect -7218 373018 591142 373254
rect 591378 373018 592500 373254
rect -8576 372934 592500 373018
rect -8576 372698 -7454 372934
rect -7218 372698 591142 372934
rect 591378 372698 592500 372934
rect -8576 372676 592500 372698
rect -7636 372674 -7036 372676
rect 590960 372674 591560 372676
rect -5756 369676 -5156 369678
rect 589080 369676 589680 369678
rect -6696 369654 590620 369676
rect -6696 369418 -5574 369654
rect -5338 369418 589262 369654
rect 589498 369418 590620 369654
rect -6696 369334 590620 369418
rect -6696 369098 -5574 369334
rect -5338 369098 589262 369334
rect 589498 369098 590620 369334
rect -6696 369076 590620 369098
rect -5756 369074 -5156 369076
rect 589080 369074 589680 369076
rect -3876 366076 -3276 366078
rect 4404 366076 5004 366078
rect 580404 366076 581004 366078
rect 587200 366076 587800 366078
rect -4816 366054 588740 366076
rect -4816 365818 -3694 366054
rect -3458 365818 4586 366054
rect 4822 365818 580586 366054
rect 580822 365818 587382 366054
rect 587618 365818 588740 366054
rect -4816 365734 588740 365818
rect -4816 365498 -3694 365734
rect -3458 365498 4586 365734
rect 4822 365498 580586 365734
rect 580822 365498 587382 365734
rect 587618 365498 588740 365734
rect -4816 365476 588740 365498
rect -3876 365474 -3276 365476
rect 4404 365474 5004 365476
rect 580404 365474 581004 365476
rect 587200 365474 587800 365476
rect -1996 362428 -1396 362430
rect 804 362428 1404 362430
rect 585320 362428 585920 362430
rect -2936 362406 586860 362428
rect -2936 362170 -1814 362406
rect -1578 362170 986 362406
rect 1222 362170 585502 362406
rect 585738 362170 586860 362406
rect -2936 362086 586860 362170
rect -2936 361850 -1814 362086
rect -1578 361850 986 362086
rect 1222 361850 585502 362086
rect 585738 361850 586860 362086
rect -2936 361828 586860 361850
rect -1996 361826 -1396 361828
rect 804 361826 1404 361828
rect 585320 361826 585920 361828
rect -8576 355276 -7976 355278
rect 591900 355276 592500 355278
rect -8576 355254 592500 355276
rect -8576 355018 -8394 355254
rect -8158 355018 592082 355254
rect 592318 355018 592500 355254
rect -8576 354934 592500 355018
rect -8576 354698 -8394 354934
rect -8158 354698 592082 354934
rect 592318 354698 592500 354934
rect -8576 354676 592500 354698
rect -8576 354674 -7976 354676
rect 591900 354674 592500 354676
rect -6696 351676 -6096 351678
rect 590020 351676 590620 351678
rect -6696 351654 590620 351676
rect -6696 351418 -6514 351654
rect -6278 351418 590202 351654
rect 590438 351418 590620 351654
rect -6696 351334 590620 351418
rect -6696 351098 -6514 351334
rect -6278 351098 590202 351334
rect 590438 351098 590620 351334
rect -6696 351076 590620 351098
rect -6696 351074 -6096 351076
rect 590020 351074 590620 351076
rect -4816 348076 -4216 348078
rect 588140 348076 588740 348078
rect -4816 348054 588740 348076
rect -4816 347818 -4634 348054
rect -4398 347818 588322 348054
rect 588558 347818 588740 348054
rect -4816 347734 588740 347818
rect -4816 347498 -4634 347734
rect -4398 347498 588322 347734
rect 588558 347498 588740 347734
rect -4816 347476 588740 347498
rect -4816 347474 -4216 347476
rect 588140 347474 588740 347476
rect -2936 344428 -2336 344430
rect 586260 344428 586860 344430
rect -2936 344406 586860 344428
rect -2936 344170 -2754 344406
rect -2518 344170 586442 344406
rect 586678 344170 586860 344406
rect -2936 344086 586860 344170
rect -2936 343850 -2754 344086
rect -2518 343850 586442 344086
rect 586678 343850 586860 344086
rect -2936 343828 586860 343850
rect -2936 343826 -2336 343828
rect 586260 343826 586860 343828
rect -7636 337276 -7036 337278
rect 590960 337276 591560 337278
rect -8576 337254 592500 337276
rect -8576 337018 -7454 337254
rect -7218 337018 591142 337254
rect 591378 337018 592500 337254
rect -8576 336934 592500 337018
rect -8576 336698 -7454 336934
rect -7218 336698 591142 336934
rect 591378 336698 592500 336934
rect -8576 336676 592500 336698
rect -7636 336674 -7036 336676
rect 590960 336674 591560 336676
rect -5756 333676 -5156 333678
rect 589080 333676 589680 333678
rect -6696 333654 590620 333676
rect -6696 333418 -5574 333654
rect -5338 333418 589262 333654
rect 589498 333418 590620 333654
rect -6696 333334 590620 333418
rect -6696 333098 -5574 333334
rect -5338 333098 589262 333334
rect 589498 333098 590620 333334
rect -6696 333076 590620 333098
rect -5756 333074 -5156 333076
rect 589080 333074 589680 333076
rect -3876 330076 -3276 330078
rect 4404 330076 5004 330078
rect 580404 330076 581004 330078
rect 587200 330076 587800 330078
rect -4816 330054 588740 330076
rect -4816 329818 -3694 330054
rect -3458 329818 4586 330054
rect 4822 329818 580586 330054
rect 580822 329818 587382 330054
rect 587618 329818 588740 330054
rect -4816 329734 588740 329818
rect -4816 329498 -3694 329734
rect -3458 329498 4586 329734
rect 4822 329498 580586 329734
rect 580822 329498 587382 329734
rect 587618 329498 588740 329734
rect -4816 329476 588740 329498
rect -3876 329474 -3276 329476
rect 4404 329474 5004 329476
rect 580404 329474 581004 329476
rect 587200 329474 587800 329476
rect -1996 326428 -1396 326430
rect 804 326428 1404 326430
rect 585320 326428 585920 326430
rect -2936 326406 586860 326428
rect -2936 326170 -1814 326406
rect -1578 326170 986 326406
rect 1222 326170 585502 326406
rect 585738 326170 586860 326406
rect -2936 326086 586860 326170
rect -2936 325850 -1814 326086
rect -1578 325850 986 326086
rect 1222 325850 585502 326086
rect 585738 325850 586860 326086
rect -2936 325828 586860 325850
rect -1996 325826 -1396 325828
rect 804 325826 1404 325828
rect 585320 325826 585920 325828
rect -8576 319276 -7976 319278
rect 591900 319276 592500 319278
rect -8576 319254 592500 319276
rect -8576 319018 -8394 319254
rect -8158 319018 592082 319254
rect 592318 319018 592500 319254
rect -8576 318934 592500 319018
rect -8576 318698 -8394 318934
rect -8158 318698 592082 318934
rect 592318 318698 592500 318934
rect -8576 318676 592500 318698
rect -8576 318674 -7976 318676
rect 591900 318674 592500 318676
rect -6696 315676 -6096 315678
rect 590020 315676 590620 315678
rect -6696 315654 590620 315676
rect -6696 315418 -6514 315654
rect -6278 315418 590202 315654
rect 590438 315418 590620 315654
rect -6696 315334 590620 315418
rect -6696 315098 -6514 315334
rect -6278 315098 590202 315334
rect 590438 315098 590620 315334
rect -6696 315076 590620 315098
rect -6696 315074 -6096 315076
rect 590020 315074 590620 315076
rect -4816 312076 -4216 312078
rect 588140 312076 588740 312078
rect -4816 312054 588740 312076
rect -4816 311818 -4634 312054
rect -4398 311818 588322 312054
rect 588558 311818 588740 312054
rect -4816 311734 588740 311818
rect -4816 311498 -4634 311734
rect -4398 311498 588322 311734
rect 588558 311498 588740 311734
rect -4816 311476 588740 311498
rect -4816 311474 -4216 311476
rect 588140 311474 588740 311476
rect -2936 308428 -2336 308430
rect 586260 308428 586860 308430
rect -2936 308406 586860 308428
rect -2936 308170 -2754 308406
rect -2518 308170 586442 308406
rect 586678 308170 586860 308406
rect -2936 308086 586860 308170
rect -2936 307850 -2754 308086
rect -2518 307850 586442 308086
rect 586678 307850 586860 308086
rect -2936 307828 586860 307850
rect -2936 307826 -2336 307828
rect 586260 307826 586860 307828
rect -7636 301276 -7036 301278
rect 590960 301276 591560 301278
rect -8576 301254 592500 301276
rect -8576 301018 -7454 301254
rect -7218 301018 591142 301254
rect 591378 301018 592500 301254
rect -8576 300934 592500 301018
rect -8576 300698 -7454 300934
rect -7218 300698 591142 300934
rect 591378 300698 592500 300934
rect -8576 300676 592500 300698
rect -7636 300674 -7036 300676
rect 590960 300674 591560 300676
rect -5756 297676 -5156 297678
rect 589080 297676 589680 297678
rect -6696 297654 590620 297676
rect -6696 297418 -5574 297654
rect -5338 297418 589262 297654
rect 589498 297418 590620 297654
rect -6696 297334 590620 297418
rect -6696 297098 -5574 297334
rect -5338 297098 589262 297334
rect 589498 297098 590620 297334
rect -6696 297076 590620 297098
rect -5756 297074 -5156 297076
rect 589080 297074 589680 297076
rect -3876 294076 -3276 294078
rect 4404 294076 5004 294078
rect 580404 294076 581004 294078
rect 587200 294076 587800 294078
rect -4816 294054 588740 294076
rect -4816 293818 -3694 294054
rect -3458 293818 4586 294054
rect 4822 293818 580586 294054
rect 580822 293818 587382 294054
rect 587618 293818 588740 294054
rect -4816 293734 588740 293818
rect -4816 293498 -3694 293734
rect -3458 293498 4586 293734
rect 4822 293498 580586 293734
rect 580822 293498 587382 293734
rect 587618 293498 588740 293734
rect -4816 293476 588740 293498
rect -3876 293474 -3276 293476
rect 4404 293474 5004 293476
rect 580404 293474 581004 293476
rect 587200 293474 587800 293476
rect -1996 290428 -1396 290430
rect 804 290428 1404 290430
rect 585320 290428 585920 290430
rect -2936 290406 586860 290428
rect -2936 290170 -1814 290406
rect -1578 290170 986 290406
rect 1222 290170 585502 290406
rect 585738 290170 586860 290406
rect -2936 290086 586860 290170
rect -2936 289850 -1814 290086
rect -1578 289850 986 290086
rect 1222 289850 585502 290086
rect 585738 289850 586860 290086
rect -2936 289828 586860 289850
rect -1996 289826 -1396 289828
rect 804 289826 1404 289828
rect 585320 289826 585920 289828
rect -8576 283276 -7976 283278
rect 591900 283276 592500 283278
rect -8576 283254 592500 283276
rect -8576 283018 -8394 283254
rect -8158 283018 592082 283254
rect 592318 283018 592500 283254
rect -8576 282934 592500 283018
rect -8576 282698 -8394 282934
rect -8158 282698 592082 282934
rect 592318 282698 592500 282934
rect -8576 282676 592500 282698
rect -8576 282674 -7976 282676
rect 591900 282674 592500 282676
rect -6696 279676 -6096 279678
rect 590020 279676 590620 279678
rect -6696 279654 590620 279676
rect -6696 279418 -6514 279654
rect -6278 279418 590202 279654
rect 590438 279418 590620 279654
rect -6696 279334 590620 279418
rect -6696 279098 -6514 279334
rect -6278 279098 590202 279334
rect 590438 279098 590620 279334
rect -6696 279076 590620 279098
rect -6696 279074 -6096 279076
rect 590020 279074 590620 279076
rect -4816 276076 -4216 276078
rect 588140 276076 588740 276078
rect -4816 276054 588740 276076
rect -4816 275818 -4634 276054
rect -4398 275818 588322 276054
rect 588558 275818 588740 276054
rect -4816 275734 588740 275818
rect -4816 275498 -4634 275734
rect -4398 275498 588322 275734
rect 588558 275498 588740 275734
rect -4816 275476 588740 275498
rect -4816 275474 -4216 275476
rect 588140 275474 588740 275476
rect -2936 272428 -2336 272430
rect 586260 272428 586860 272430
rect -2936 272406 586860 272428
rect -2936 272170 -2754 272406
rect -2518 272170 586442 272406
rect 586678 272170 586860 272406
rect -2936 272086 586860 272170
rect -2936 271850 -2754 272086
rect -2518 271850 586442 272086
rect 586678 271850 586860 272086
rect -2936 271828 586860 271850
rect -2936 271826 -2336 271828
rect 586260 271826 586860 271828
rect -7636 265276 -7036 265278
rect 590960 265276 591560 265278
rect -8576 265254 592500 265276
rect -8576 265018 -7454 265254
rect -7218 265018 591142 265254
rect 591378 265018 592500 265254
rect -8576 264934 592500 265018
rect -8576 264698 -7454 264934
rect -7218 264698 591142 264934
rect 591378 264698 592500 264934
rect -8576 264676 592500 264698
rect -7636 264674 -7036 264676
rect 590960 264674 591560 264676
rect -5756 261676 -5156 261678
rect 589080 261676 589680 261678
rect -6696 261654 590620 261676
rect -6696 261418 -5574 261654
rect -5338 261418 589262 261654
rect 589498 261418 590620 261654
rect -6696 261334 590620 261418
rect -6696 261098 -5574 261334
rect -5338 261098 589262 261334
rect 589498 261098 590620 261334
rect -6696 261076 590620 261098
rect -5756 261074 -5156 261076
rect 589080 261074 589680 261076
rect -3876 258076 -3276 258078
rect 4404 258076 5004 258078
rect 580404 258076 581004 258078
rect 587200 258076 587800 258078
rect -4816 258054 588740 258076
rect -4816 257818 -3694 258054
rect -3458 257818 4586 258054
rect 4822 257818 580586 258054
rect 580822 257818 587382 258054
rect 587618 257818 588740 258054
rect -4816 257734 588740 257818
rect -4816 257498 -3694 257734
rect -3458 257498 4586 257734
rect 4822 257498 580586 257734
rect 580822 257498 587382 257734
rect 587618 257498 588740 257734
rect -4816 257476 588740 257498
rect -3876 257474 -3276 257476
rect 4404 257474 5004 257476
rect 580404 257474 581004 257476
rect 587200 257474 587800 257476
rect -1996 254428 -1396 254430
rect 804 254428 1404 254430
rect 585320 254428 585920 254430
rect -2936 254406 586860 254428
rect -2936 254170 -1814 254406
rect -1578 254170 986 254406
rect 1222 254170 585502 254406
rect 585738 254170 586860 254406
rect -2936 254086 586860 254170
rect -2936 253850 -1814 254086
rect -1578 253850 986 254086
rect 1222 253850 585502 254086
rect 585738 253850 586860 254086
rect -2936 253828 586860 253850
rect -1996 253826 -1396 253828
rect 804 253826 1404 253828
rect 585320 253826 585920 253828
rect -8576 247276 -7976 247278
rect 591900 247276 592500 247278
rect -8576 247254 592500 247276
rect -8576 247018 -8394 247254
rect -8158 247018 592082 247254
rect 592318 247018 592500 247254
rect -8576 246934 592500 247018
rect -8576 246698 -8394 246934
rect -8158 246698 592082 246934
rect 592318 246698 592500 246934
rect -8576 246676 592500 246698
rect -8576 246674 -7976 246676
rect 591900 246674 592500 246676
rect -6696 243676 -6096 243678
rect 590020 243676 590620 243678
rect -6696 243654 590620 243676
rect -6696 243418 -6514 243654
rect -6278 243418 590202 243654
rect 590438 243418 590620 243654
rect -6696 243334 590620 243418
rect -6696 243098 -6514 243334
rect -6278 243098 590202 243334
rect 590438 243098 590620 243334
rect -6696 243076 590620 243098
rect -6696 243074 -6096 243076
rect 590020 243074 590620 243076
rect -4816 240076 -4216 240078
rect 588140 240076 588740 240078
rect -4816 240054 588740 240076
rect -4816 239818 -4634 240054
rect -4398 239818 588322 240054
rect 588558 239818 588740 240054
rect -4816 239734 588740 239818
rect -4816 239498 -4634 239734
rect -4398 239498 588322 239734
rect 588558 239498 588740 239734
rect -4816 239476 588740 239498
rect -4816 239474 -4216 239476
rect 588140 239474 588740 239476
rect -2936 236428 -2336 236430
rect 586260 236428 586860 236430
rect -2936 236406 586860 236428
rect -2936 236170 -2754 236406
rect -2518 236170 586442 236406
rect 586678 236170 586860 236406
rect -2936 236086 586860 236170
rect -2936 235850 -2754 236086
rect -2518 235850 586442 236086
rect 586678 235850 586860 236086
rect -2936 235828 586860 235850
rect -2936 235826 -2336 235828
rect 586260 235826 586860 235828
rect -7636 229276 -7036 229278
rect 590960 229276 591560 229278
rect -8576 229254 592500 229276
rect -8576 229018 -7454 229254
rect -7218 229018 591142 229254
rect 591378 229018 592500 229254
rect -8576 228934 592500 229018
rect -8576 228698 -7454 228934
rect -7218 228698 591142 228934
rect 591378 228698 592500 228934
rect -8576 228676 592500 228698
rect -7636 228674 -7036 228676
rect 590960 228674 591560 228676
rect -5756 225676 -5156 225678
rect 589080 225676 589680 225678
rect -6696 225654 590620 225676
rect -6696 225418 -5574 225654
rect -5338 225418 589262 225654
rect 589498 225418 590620 225654
rect -6696 225334 590620 225418
rect -6696 225098 -5574 225334
rect -5338 225098 589262 225334
rect 589498 225098 590620 225334
rect -6696 225076 590620 225098
rect -5756 225074 -5156 225076
rect 589080 225074 589680 225076
rect -3876 222076 -3276 222078
rect 4404 222076 5004 222078
rect 580404 222076 581004 222078
rect 587200 222076 587800 222078
rect -4816 222054 588740 222076
rect -4816 221818 -3694 222054
rect -3458 221818 4586 222054
rect 4822 221818 580586 222054
rect 580822 221818 587382 222054
rect 587618 221818 588740 222054
rect -4816 221734 588740 221818
rect -4816 221498 -3694 221734
rect -3458 221498 4586 221734
rect 4822 221498 580586 221734
rect 580822 221498 587382 221734
rect 587618 221498 588740 221734
rect -4816 221476 588740 221498
rect -3876 221474 -3276 221476
rect 4404 221474 5004 221476
rect 580404 221474 581004 221476
rect 587200 221474 587800 221476
rect -1996 218428 -1396 218430
rect 804 218428 1404 218430
rect 585320 218428 585920 218430
rect -2936 218406 586860 218428
rect -2936 218170 -1814 218406
rect -1578 218170 986 218406
rect 1222 218170 585502 218406
rect 585738 218170 586860 218406
rect -2936 218086 586860 218170
rect -2936 217850 -1814 218086
rect -1578 217850 986 218086
rect 1222 217850 585502 218086
rect 585738 217850 586860 218086
rect -2936 217828 586860 217850
rect -1996 217826 -1396 217828
rect 804 217826 1404 217828
rect 585320 217826 585920 217828
rect -8576 211276 -7976 211278
rect 591900 211276 592500 211278
rect -8576 211254 592500 211276
rect -8576 211018 -8394 211254
rect -8158 211018 592082 211254
rect 592318 211018 592500 211254
rect -8576 210934 592500 211018
rect -8576 210698 -8394 210934
rect -8158 210698 592082 210934
rect 592318 210698 592500 210934
rect -8576 210676 592500 210698
rect -8576 210674 -7976 210676
rect 591900 210674 592500 210676
rect -6696 207676 -6096 207678
rect 590020 207676 590620 207678
rect -6696 207654 590620 207676
rect -6696 207418 -6514 207654
rect -6278 207418 590202 207654
rect 590438 207418 590620 207654
rect -6696 207334 590620 207418
rect -6696 207098 -6514 207334
rect -6278 207098 590202 207334
rect 590438 207098 590620 207334
rect -6696 207076 590620 207098
rect -6696 207074 -6096 207076
rect 590020 207074 590620 207076
rect -4816 204076 -4216 204078
rect 588140 204076 588740 204078
rect -4816 204054 588740 204076
rect -4816 203818 -4634 204054
rect -4398 203818 588322 204054
rect 588558 203818 588740 204054
rect -4816 203734 588740 203818
rect -4816 203498 -4634 203734
rect -4398 203498 588322 203734
rect 588558 203498 588740 203734
rect -4816 203476 588740 203498
rect -4816 203474 -4216 203476
rect 588140 203474 588740 203476
rect -2936 200428 -2336 200430
rect 586260 200428 586860 200430
rect -2936 200406 586860 200428
rect -2936 200170 -2754 200406
rect -2518 200170 586442 200406
rect 586678 200170 586860 200406
rect -2936 200086 586860 200170
rect -2936 199850 -2754 200086
rect -2518 199850 586442 200086
rect 586678 199850 586860 200086
rect -2936 199828 586860 199850
rect -2936 199826 -2336 199828
rect 586260 199826 586860 199828
rect -7636 193276 -7036 193278
rect 590960 193276 591560 193278
rect -8576 193254 592500 193276
rect -8576 193018 -7454 193254
rect -7218 193018 591142 193254
rect 591378 193018 592500 193254
rect -8576 192934 592500 193018
rect -8576 192698 -7454 192934
rect -7218 192698 591142 192934
rect 591378 192698 592500 192934
rect -8576 192676 592500 192698
rect -7636 192674 -7036 192676
rect 590960 192674 591560 192676
rect -5756 189676 -5156 189678
rect 589080 189676 589680 189678
rect -6696 189654 590620 189676
rect -6696 189418 -5574 189654
rect -5338 189418 589262 189654
rect 589498 189418 590620 189654
rect -6696 189334 590620 189418
rect -6696 189098 -5574 189334
rect -5338 189098 589262 189334
rect 589498 189098 590620 189334
rect -6696 189076 590620 189098
rect -5756 189074 -5156 189076
rect 589080 189074 589680 189076
rect -3876 186076 -3276 186078
rect 4404 186076 5004 186078
rect 580404 186076 581004 186078
rect 587200 186076 587800 186078
rect -4816 186054 588740 186076
rect -4816 185818 -3694 186054
rect -3458 185818 4586 186054
rect 4822 185818 580586 186054
rect 580822 185818 587382 186054
rect 587618 185818 588740 186054
rect -4816 185734 588740 185818
rect -4816 185498 -3694 185734
rect -3458 185498 4586 185734
rect 4822 185498 580586 185734
rect 580822 185498 587382 185734
rect 587618 185498 588740 185734
rect -4816 185476 588740 185498
rect -3876 185474 -3276 185476
rect 4404 185474 5004 185476
rect 580404 185474 581004 185476
rect 587200 185474 587800 185476
rect -1996 182428 -1396 182430
rect 804 182428 1404 182430
rect 585320 182428 585920 182430
rect -2936 182406 586860 182428
rect -2936 182170 -1814 182406
rect -1578 182170 986 182406
rect 1222 182170 585502 182406
rect 585738 182170 586860 182406
rect -2936 182086 586860 182170
rect -2936 181850 -1814 182086
rect -1578 181850 986 182086
rect 1222 181850 585502 182086
rect 585738 181850 586860 182086
rect -2936 181828 586860 181850
rect -1996 181826 -1396 181828
rect 804 181826 1404 181828
rect 585320 181826 585920 181828
rect -8576 175276 -7976 175278
rect 591900 175276 592500 175278
rect -8576 175254 592500 175276
rect -8576 175018 -8394 175254
rect -8158 175018 592082 175254
rect 592318 175018 592500 175254
rect -8576 174934 592500 175018
rect -8576 174698 -8394 174934
rect -8158 174698 592082 174934
rect 592318 174698 592500 174934
rect -8576 174676 592500 174698
rect -8576 174674 -7976 174676
rect 591900 174674 592500 174676
rect -6696 171676 -6096 171678
rect 590020 171676 590620 171678
rect -6696 171654 590620 171676
rect -6696 171418 -6514 171654
rect -6278 171418 590202 171654
rect 590438 171418 590620 171654
rect -6696 171334 590620 171418
rect -6696 171098 -6514 171334
rect -6278 171098 590202 171334
rect 590438 171098 590620 171334
rect -6696 171076 590620 171098
rect -6696 171074 -6096 171076
rect 590020 171074 590620 171076
rect -4816 168076 -4216 168078
rect 588140 168076 588740 168078
rect -4816 168054 588740 168076
rect -4816 167818 -4634 168054
rect -4398 167818 588322 168054
rect 588558 167818 588740 168054
rect -4816 167734 588740 167818
rect -4816 167498 -4634 167734
rect -4398 167498 588322 167734
rect 588558 167498 588740 167734
rect -4816 167476 588740 167498
rect -4816 167474 -4216 167476
rect 588140 167474 588740 167476
rect -2936 164428 -2336 164430
rect 586260 164428 586860 164430
rect -2936 164406 586860 164428
rect -2936 164170 -2754 164406
rect -2518 164170 586442 164406
rect 586678 164170 586860 164406
rect -2936 164086 586860 164170
rect -2936 163850 -2754 164086
rect -2518 163850 586442 164086
rect 586678 163850 586860 164086
rect -2936 163828 586860 163850
rect -2936 163826 -2336 163828
rect 586260 163826 586860 163828
rect -7636 157276 -7036 157278
rect 590960 157276 591560 157278
rect -8576 157254 592500 157276
rect -8576 157018 -7454 157254
rect -7218 157018 591142 157254
rect 591378 157018 592500 157254
rect -8576 156934 592500 157018
rect -8576 156698 -7454 156934
rect -7218 156698 591142 156934
rect 591378 156698 592500 156934
rect -8576 156676 592500 156698
rect -7636 156674 -7036 156676
rect 590960 156674 591560 156676
rect -5756 153676 -5156 153678
rect 589080 153676 589680 153678
rect -6696 153654 590620 153676
rect -6696 153418 -5574 153654
rect -5338 153418 589262 153654
rect 589498 153418 590620 153654
rect -6696 153334 590620 153418
rect -6696 153098 -5574 153334
rect -5338 153098 589262 153334
rect 589498 153098 590620 153334
rect -6696 153076 590620 153098
rect -5756 153074 -5156 153076
rect 589080 153074 589680 153076
rect -3876 150076 -3276 150078
rect 4404 150076 5004 150078
rect 580404 150076 581004 150078
rect 587200 150076 587800 150078
rect -4816 150054 588740 150076
rect -4816 149818 -3694 150054
rect -3458 149818 4586 150054
rect 4822 149818 580586 150054
rect 580822 149818 587382 150054
rect 587618 149818 588740 150054
rect -4816 149734 588740 149818
rect -4816 149498 -3694 149734
rect -3458 149498 4586 149734
rect 4822 149498 580586 149734
rect 580822 149498 587382 149734
rect 587618 149498 588740 149734
rect -4816 149476 588740 149498
rect -3876 149474 -3276 149476
rect 4404 149474 5004 149476
rect 580404 149474 581004 149476
rect 587200 149474 587800 149476
rect -1996 146428 -1396 146430
rect 804 146428 1404 146430
rect 585320 146428 585920 146430
rect -2936 146406 586860 146428
rect -2936 146170 -1814 146406
rect -1578 146170 986 146406
rect 1222 146170 585502 146406
rect 585738 146170 586860 146406
rect -2936 146086 586860 146170
rect -2936 145850 -1814 146086
rect -1578 145850 986 146086
rect 1222 145850 585502 146086
rect 585738 145850 586860 146086
rect -2936 145828 586860 145850
rect -1996 145826 -1396 145828
rect 804 145826 1404 145828
rect 585320 145826 585920 145828
rect -8576 139276 -7976 139278
rect 591900 139276 592500 139278
rect -8576 139254 592500 139276
rect -8576 139018 -8394 139254
rect -8158 139018 592082 139254
rect 592318 139018 592500 139254
rect -8576 138934 592500 139018
rect -8576 138698 -8394 138934
rect -8158 138698 592082 138934
rect 592318 138698 592500 138934
rect -8576 138676 592500 138698
rect -8576 138674 -7976 138676
rect 591900 138674 592500 138676
rect -6696 135676 -6096 135678
rect 590020 135676 590620 135678
rect -6696 135654 590620 135676
rect -6696 135418 -6514 135654
rect -6278 135418 590202 135654
rect 590438 135418 590620 135654
rect -6696 135334 590620 135418
rect -6696 135098 -6514 135334
rect -6278 135098 590202 135334
rect 590438 135098 590620 135334
rect -6696 135076 590620 135098
rect -6696 135074 -6096 135076
rect 590020 135074 590620 135076
rect -4816 132076 -4216 132078
rect 588140 132076 588740 132078
rect -4816 132054 588740 132076
rect -4816 131818 -4634 132054
rect -4398 131818 588322 132054
rect 588558 131818 588740 132054
rect -4816 131734 588740 131818
rect -4816 131498 -4634 131734
rect -4398 131498 588322 131734
rect 588558 131498 588740 131734
rect -4816 131476 588740 131498
rect -4816 131474 -4216 131476
rect 588140 131474 588740 131476
rect -2936 128428 -2336 128430
rect 586260 128428 586860 128430
rect -2936 128406 586860 128428
rect -2936 128170 -2754 128406
rect -2518 128170 586442 128406
rect 586678 128170 586860 128406
rect -2936 128086 586860 128170
rect -2936 127850 -2754 128086
rect -2518 127850 586442 128086
rect 586678 127850 586860 128086
rect -2936 127828 586860 127850
rect -2936 127826 -2336 127828
rect 586260 127826 586860 127828
rect -7636 121276 -7036 121278
rect 590960 121276 591560 121278
rect -8576 121254 592500 121276
rect -8576 121018 -7454 121254
rect -7218 121018 591142 121254
rect 591378 121018 592500 121254
rect -8576 120934 592500 121018
rect -8576 120698 -7454 120934
rect -7218 120698 591142 120934
rect 591378 120698 592500 120934
rect -8576 120676 592500 120698
rect -7636 120674 -7036 120676
rect 590960 120674 591560 120676
rect -5756 117676 -5156 117678
rect 589080 117676 589680 117678
rect -6696 117654 590620 117676
rect -6696 117418 -5574 117654
rect -5338 117418 589262 117654
rect 589498 117418 590620 117654
rect -6696 117334 590620 117418
rect -6696 117098 -5574 117334
rect -5338 117098 589262 117334
rect 589498 117098 590620 117334
rect -6696 117076 590620 117098
rect -5756 117074 -5156 117076
rect 589080 117074 589680 117076
rect -3876 114076 -3276 114078
rect 4404 114076 5004 114078
rect 580404 114076 581004 114078
rect 587200 114076 587800 114078
rect -4816 114054 588740 114076
rect -4816 113818 -3694 114054
rect -3458 113818 4586 114054
rect 4822 113818 580586 114054
rect 580822 113818 587382 114054
rect 587618 113818 588740 114054
rect -4816 113734 588740 113818
rect -4816 113498 -3694 113734
rect -3458 113498 4586 113734
rect 4822 113498 580586 113734
rect 580822 113498 587382 113734
rect 587618 113498 588740 113734
rect -4816 113476 588740 113498
rect -3876 113474 -3276 113476
rect 4404 113474 5004 113476
rect 580404 113474 581004 113476
rect 587200 113474 587800 113476
rect -1996 110428 -1396 110430
rect 804 110428 1404 110430
rect 585320 110428 585920 110430
rect -2936 110406 586860 110428
rect -2936 110170 -1814 110406
rect -1578 110170 986 110406
rect 1222 110170 585502 110406
rect 585738 110170 586860 110406
rect -2936 110086 586860 110170
rect -2936 109850 -1814 110086
rect -1578 109850 986 110086
rect 1222 109850 585502 110086
rect 585738 109850 586860 110086
rect -2936 109828 586860 109850
rect -1996 109826 -1396 109828
rect 804 109826 1404 109828
rect 585320 109826 585920 109828
rect -8576 103276 -7976 103278
rect 591900 103276 592500 103278
rect -8576 103254 592500 103276
rect -8576 103018 -8394 103254
rect -8158 103018 592082 103254
rect 592318 103018 592500 103254
rect -8576 102934 592500 103018
rect -8576 102698 -8394 102934
rect -8158 102698 592082 102934
rect 592318 102698 592500 102934
rect -8576 102676 592500 102698
rect -8576 102674 -7976 102676
rect 591900 102674 592500 102676
rect -6696 99676 -6096 99678
rect 590020 99676 590620 99678
rect -6696 99654 590620 99676
rect -6696 99418 -6514 99654
rect -6278 99418 590202 99654
rect 590438 99418 590620 99654
rect -6696 99334 590620 99418
rect -6696 99098 -6514 99334
rect -6278 99098 590202 99334
rect 590438 99098 590620 99334
rect -6696 99076 590620 99098
rect -6696 99074 -6096 99076
rect 590020 99074 590620 99076
rect -4816 96076 -4216 96078
rect 588140 96076 588740 96078
rect -4816 96054 588740 96076
rect -4816 95818 -4634 96054
rect -4398 95818 588322 96054
rect 588558 95818 588740 96054
rect -4816 95734 588740 95818
rect -4816 95498 -4634 95734
rect -4398 95498 588322 95734
rect 588558 95498 588740 95734
rect -4816 95476 588740 95498
rect -4816 95474 -4216 95476
rect 588140 95474 588740 95476
rect -2936 92428 -2336 92430
rect 586260 92428 586860 92430
rect -2936 92406 586860 92428
rect -2936 92170 -2754 92406
rect -2518 92170 586442 92406
rect 586678 92170 586860 92406
rect -2936 92086 586860 92170
rect -2936 91850 -2754 92086
rect -2518 91850 586442 92086
rect 586678 91850 586860 92086
rect -2936 91828 586860 91850
rect -2936 91826 -2336 91828
rect 586260 91826 586860 91828
rect -7636 85276 -7036 85278
rect 590960 85276 591560 85278
rect -8576 85254 592500 85276
rect -8576 85018 -7454 85254
rect -7218 85018 591142 85254
rect 591378 85018 592500 85254
rect -8576 84934 592500 85018
rect -8576 84698 -7454 84934
rect -7218 84698 591142 84934
rect 591378 84698 592500 84934
rect -8576 84676 592500 84698
rect -7636 84674 -7036 84676
rect 590960 84674 591560 84676
rect -5756 81676 -5156 81678
rect 589080 81676 589680 81678
rect -6696 81654 590620 81676
rect -6696 81418 -5574 81654
rect -5338 81418 589262 81654
rect 589498 81418 590620 81654
rect -6696 81334 590620 81418
rect -6696 81098 -5574 81334
rect -5338 81098 589262 81334
rect 589498 81098 590620 81334
rect -6696 81076 590620 81098
rect -5756 81074 -5156 81076
rect 589080 81074 589680 81076
rect -3876 78076 -3276 78078
rect 4404 78076 5004 78078
rect 580404 78076 581004 78078
rect 587200 78076 587800 78078
rect -4816 78054 588740 78076
rect -4816 77818 -3694 78054
rect -3458 77818 4586 78054
rect 4822 77818 580586 78054
rect 580822 77818 587382 78054
rect 587618 77818 588740 78054
rect -4816 77734 588740 77818
rect -4816 77498 -3694 77734
rect -3458 77498 4586 77734
rect 4822 77498 580586 77734
rect 580822 77498 587382 77734
rect 587618 77498 588740 77734
rect -4816 77476 588740 77498
rect -3876 77474 -3276 77476
rect 4404 77474 5004 77476
rect 580404 77474 581004 77476
rect 587200 77474 587800 77476
rect -1996 74428 -1396 74430
rect 804 74428 1404 74430
rect 585320 74428 585920 74430
rect -2936 74406 586860 74428
rect -2936 74170 -1814 74406
rect -1578 74170 986 74406
rect 1222 74170 585502 74406
rect 585738 74170 586860 74406
rect -2936 74086 586860 74170
rect -2936 73850 -1814 74086
rect -1578 73850 986 74086
rect 1222 73850 585502 74086
rect 585738 73850 586860 74086
rect -2936 73828 586860 73850
rect -1996 73826 -1396 73828
rect 804 73826 1404 73828
rect 585320 73826 585920 73828
rect -8576 67276 -7976 67278
rect 591900 67276 592500 67278
rect -8576 67254 592500 67276
rect -8576 67018 -8394 67254
rect -8158 67018 592082 67254
rect 592318 67018 592500 67254
rect -8576 66934 592500 67018
rect -8576 66698 -8394 66934
rect -8158 66698 592082 66934
rect 592318 66698 592500 66934
rect -8576 66676 592500 66698
rect -8576 66674 -7976 66676
rect 591900 66674 592500 66676
rect -6696 63676 -6096 63678
rect 590020 63676 590620 63678
rect -6696 63654 590620 63676
rect -6696 63418 -6514 63654
rect -6278 63418 590202 63654
rect 590438 63418 590620 63654
rect -6696 63334 590620 63418
rect -6696 63098 -6514 63334
rect -6278 63098 590202 63334
rect 590438 63098 590620 63334
rect -6696 63076 590620 63098
rect -6696 63074 -6096 63076
rect 590020 63074 590620 63076
rect -4816 60076 -4216 60078
rect 588140 60076 588740 60078
rect -4816 60054 588740 60076
rect -4816 59818 -4634 60054
rect -4398 59818 588322 60054
rect 588558 59818 588740 60054
rect -4816 59734 588740 59818
rect -4816 59498 -4634 59734
rect -4398 59498 588322 59734
rect 588558 59498 588740 59734
rect -4816 59476 588740 59498
rect -4816 59474 -4216 59476
rect 588140 59474 588740 59476
rect -2936 56428 -2336 56430
rect 586260 56428 586860 56430
rect -2936 56406 586860 56428
rect -2936 56170 -2754 56406
rect -2518 56170 586442 56406
rect 586678 56170 586860 56406
rect -2936 56086 586860 56170
rect -2936 55850 -2754 56086
rect -2518 55850 586442 56086
rect 586678 55850 586860 56086
rect -2936 55828 586860 55850
rect -2936 55826 -2336 55828
rect 586260 55826 586860 55828
rect -7636 49276 -7036 49278
rect 590960 49276 591560 49278
rect -8576 49254 592500 49276
rect -8576 49018 -7454 49254
rect -7218 49018 591142 49254
rect 591378 49018 592500 49254
rect -8576 48934 592500 49018
rect -8576 48698 -7454 48934
rect -7218 48698 591142 48934
rect 591378 48698 592500 48934
rect -8576 48676 592500 48698
rect -7636 48674 -7036 48676
rect 590960 48674 591560 48676
rect -5756 45676 -5156 45678
rect 589080 45676 589680 45678
rect -6696 45654 590620 45676
rect -6696 45418 -5574 45654
rect -5338 45418 589262 45654
rect 589498 45418 590620 45654
rect -6696 45334 590620 45418
rect -6696 45098 -5574 45334
rect -5338 45098 589262 45334
rect 589498 45098 590620 45334
rect -6696 45076 590620 45098
rect -5756 45074 -5156 45076
rect 589080 45074 589680 45076
rect -3876 42076 -3276 42078
rect 4404 42076 5004 42078
rect 580404 42076 581004 42078
rect 587200 42076 587800 42078
rect -4816 42054 588740 42076
rect -4816 41818 -3694 42054
rect -3458 41818 4586 42054
rect 4822 41818 580586 42054
rect 580822 41818 587382 42054
rect 587618 41818 588740 42054
rect -4816 41734 588740 41818
rect -4816 41498 -3694 41734
rect -3458 41498 4586 41734
rect 4822 41498 580586 41734
rect 580822 41498 587382 41734
rect 587618 41498 588740 41734
rect -4816 41476 588740 41498
rect -3876 41474 -3276 41476
rect 4404 41474 5004 41476
rect 580404 41474 581004 41476
rect 587200 41474 587800 41476
rect -1996 38428 -1396 38430
rect 804 38428 1404 38430
rect 585320 38428 585920 38430
rect -2936 38406 586860 38428
rect -2936 38170 -1814 38406
rect -1578 38170 986 38406
rect 1222 38170 585502 38406
rect 585738 38170 586860 38406
rect -2936 38086 586860 38170
rect -2936 37850 -1814 38086
rect -1578 37850 986 38086
rect 1222 37850 585502 38086
rect 585738 37850 586860 38086
rect -2936 37828 586860 37850
rect -1996 37826 -1396 37828
rect 804 37826 1404 37828
rect 585320 37826 585920 37828
rect -8576 31276 -7976 31278
rect 591900 31276 592500 31278
rect -8576 31254 592500 31276
rect -8576 31018 -8394 31254
rect -8158 31018 592082 31254
rect 592318 31018 592500 31254
rect -8576 30934 592500 31018
rect -8576 30698 -8394 30934
rect -8158 30698 592082 30934
rect 592318 30698 592500 30934
rect -8576 30676 592500 30698
rect -8576 30674 -7976 30676
rect 591900 30674 592500 30676
rect -6696 27676 -6096 27678
rect 590020 27676 590620 27678
rect -6696 27654 590620 27676
rect -6696 27418 -6514 27654
rect -6278 27418 590202 27654
rect 590438 27418 590620 27654
rect -6696 27334 590620 27418
rect -6696 27098 -6514 27334
rect -6278 27098 590202 27334
rect 590438 27098 590620 27334
rect -6696 27076 590620 27098
rect -6696 27074 -6096 27076
rect 590020 27074 590620 27076
rect -4816 24076 -4216 24078
rect 588140 24076 588740 24078
rect -4816 24054 588740 24076
rect -4816 23818 -4634 24054
rect -4398 23818 588322 24054
rect 588558 23818 588740 24054
rect -4816 23734 588740 23818
rect -4816 23498 -4634 23734
rect -4398 23498 588322 23734
rect 588558 23498 588740 23734
rect -4816 23476 588740 23498
rect -4816 23474 -4216 23476
rect 588140 23474 588740 23476
rect -2936 20428 -2336 20430
rect 586260 20428 586860 20430
rect -2936 20406 586860 20428
rect -2936 20170 -2754 20406
rect -2518 20170 586442 20406
rect 586678 20170 586860 20406
rect -2936 20086 586860 20170
rect -2936 19850 -2754 20086
rect -2518 19850 586442 20086
rect 586678 19850 586860 20086
rect -2936 19828 586860 19850
rect -2936 19826 -2336 19828
rect 586260 19826 586860 19828
rect -7636 13276 -7036 13278
rect 590960 13276 591560 13278
rect -8576 13254 592500 13276
rect -8576 13018 -7454 13254
rect -7218 13018 591142 13254
rect 591378 13018 592500 13254
rect -8576 12934 592500 13018
rect -8576 12698 -7454 12934
rect -7218 12698 591142 12934
rect 591378 12698 592500 12934
rect -8576 12676 592500 12698
rect -7636 12674 -7036 12676
rect 590960 12674 591560 12676
rect -5756 9676 -5156 9678
rect 589080 9676 589680 9678
rect -6696 9654 590620 9676
rect -6696 9418 -5574 9654
rect -5338 9418 589262 9654
rect 589498 9418 590620 9654
rect -6696 9334 590620 9418
rect -6696 9098 -5574 9334
rect -5338 9098 589262 9334
rect 589498 9098 590620 9334
rect -6696 9076 590620 9098
rect -5756 9074 -5156 9076
rect 589080 9074 589680 9076
rect -3876 6076 -3276 6078
rect 4404 6076 5004 6078
rect 580404 6076 581004 6078
rect 587200 6076 587800 6078
rect -4816 6054 588740 6076
rect -4816 5818 -3694 6054
rect -3458 5818 4586 6054
rect 4822 5818 580586 6054
rect 580822 5818 587382 6054
rect 587618 5818 588740 6054
rect -4816 5734 588740 5818
rect -4816 5498 -3694 5734
rect -3458 5498 4586 5734
rect 4822 5498 580586 5734
rect 580822 5498 587382 5734
rect 587618 5498 588740 5734
rect -4816 5476 588740 5498
rect -3876 5474 -3276 5476
rect 4404 5474 5004 5476
rect 580404 5474 581004 5476
rect 587200 5474 587800 5476
rect -1996 2428 -1396 2430
rect 804 2428 1404 2430
rect 36804 2428 37404 2430
rect 72804 2428 73404 2430
rect 108804 2428 109404 2430
rect 144804 2428 145404 2430
rect 180804 2428 181404 2430
rect 216804 2428 217404 2430
rect 252804 2428 253404 2430
rect 288804 2428 289404 2430
rect 324804 2428 325404 2430
rect 360804 2428 361404 2430
rect 396804 2428 397404 2430
rect 432804 2428 433404 2430
rect 468804 2428 469404 2430
rect 504804 2428 505404 2430
rect 540804 2428 541404 2430
rect 576804 2428 577404 2430
rect 585320 2428 585920 2430
rect -2936 2406 586860 2428
rect -2936 2170 -1814 2406
rect -1578 2170 986 2406
rect 1222 2170 36986 2406
rect 37222 2170 72986 2406
rect 73222 2170 108986 2406
rect 109222 2170 144986 2406
rect 145222 2170 180986 2406
rect 181222 2170 216986 2406
rect 217222 2170 252986 2406
rect 253222 2170 288986 2406
rect 289222 2170 324986 2406
rect 325222 2170 360986 2406
rect 361222 2170 396986 2406
rect 397222 2170 432986 2406
rect 433222 2170 468986 2406
rect 469222 2170 504986 2406
rect 505222 2170 540986 2406
rect 541222 2170 576986 2406
rect 577222 2170 585502 2406
rect 585738 2170 586860 2406
rect -2936 2086 586860 2170
rect -2936 1850 -1814 2086
rect -1578 1850 986 2086
rect 1222 1850 36986 2086
rect 37222 1850 72986 2086
rect 73222 1850 108986 2086
rect 109222 1850 144986 2086
rect 145222 1850 180986 2086
rect 181222 1850 216986 2086
rect 217222 1850 252986 2086
rect 253222 1850 288986 2086
rect 289222 1850 324986 2086
rect 325222 1850 360986 2086
rect 361222 1850 396986 2086
rect 397222 1850 432986 2086
rect 433222 1850 468986 2086
rect 469222 1850 504986 2086
rect 505222 1850 540986 2086
rect 541222 1850 576986 2086
rect 577222 1850 585502 2086
rect 585738 1850 586860 2086
rect -2936 1828 586860 1850
rect -1996 1826 -1396 1828
rect 804 1826 1404 1828
rect 36804 1826 37404 1828
rect 72804 1826 73404 1828
rect 108804 1826 109404 1828
rect 144804 1826 145404 1828
rect 180804 1826 181404 1828
rect 216804 1826 217404 1828
rect 252804 1826 253404 1828
rect 288804 1826 289404 1828
rect 324804 1826 325404 1828
rect 360804 1826 361404 1828
rect 396804 1826 397404 1828
rect 432804 1826 433404 1828
rect 468804 1826 469404 1828
rect 504804 1826 505404 1828
rect 540804 1826 541404 1828
rect 576804 1826 577404 1828
rect 585320 1826 585920 1828
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2936 -1264 -2336 -1262
rect 18804 -1264 19404 -1262
rect 54804 -1264 55404 -1262
rect 90804 -1264 91404 -1262
rect 126804 -1264 127404 -1262
rect 162804 -1264 163404 -1262
rect 198804 -1264 199404 -1262
rect 234804 -1264 235404 -1262
rect 270804 -1264 271404 -1262
rect 306804 -1264 307404 -1262
rect 342804 -1264 343404 -1262
rect 378804 -1264 379404 -1262
rect 414804 -1264 415404 -1262
rect 450804 -1264 451404 -1262
rect 486804 -1264 487404 -1262
rect 522804 -1264 523404 -1262
rect 558804 -1264 559404 -1262
rect 586260 -1264 586860 -1262
rect -2936 -1286 586860 -1264
rect -2936 -1522 -2754 -1286
rect -2518 -1522 18986 -1286
rect 19222 -1522 54986 -1286
rect 55222 -1522 90986 -1286
rect 91222 -1522 126986 -1286
rect 127222 -1522 162986 -1286
rect 163222 -1522 198986 -1286
rect 199222 -1522 234986 -1286
rect 235222 -1522 270986 -1286
rect 271222 -1522 306986 -1286
rect 307222 -1522 342986 -1286
rect 343222 -1522 378986 -1286
rect 379222 -1522 414986 -1286
rect 415222 -1522 450986 -1286
rect 451222 -1522 486986 -1286
rect 487222 -1522 522986 -1286
rect 523222 -1522 558986 -1286
rect 559222 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect -2936 -1606 586860 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 18986 -1606
rect 19222 -1842 54986 -1606
rect 55222 -1842 90986 -1606
rect 91222 -1842 126986 -1606
rect 127222 -1842 162986 -1606
rect 163222 -1842 198986 -1606
rect 199222 -1842 234986 -1606
rect 235222 -1842 270986 -1606
rect 271222 -1842 306986 -1606
rect 307222 -1842 342986 -1606
rect 343222 -1842 378986 -1606
rect 379222 -1842 414986 -1606
rect 415222 -1842 450986 -1606
rect 451222 -1842 486986 -1606
rect 487222 -1842 522986 -1606
rect 523222 -1842 558986 -1606
rect 559222 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect -2936 -1864 586860 -1842
rect -2936 -1866 -2336 -1864
rect 18804 -1866 19404 -1864
rect 54804 -1866 55404 -1864
rect 90804 -1866 91404 -1864
rect 126804 -1866 127404 -1864
rect 162804 -1866 163404 -1864
rect 198804 -1866 199404 -1864
rect 234804 -1866 235404 -1864
rect 270804 -1866 271404 -1864
rect 306804 -1866 307404 -1864
rect 342804 -1866 343404 -1864
rect 378804 -1866 379404 -1864
rect 414804 -1866 415404 -1864
rect 450804 -1866 451404 -1864
rect 486804 -1866 487404 -1864
rect 522804 -1866 523404 -1864
rect 558804 -1866 559404 -1864
rect 586260 -1866 586860 -1864
rect -3876 -2204 -3276 -2202
rect 4404 -2204 5004 -2202
rect 40404 -2204 41004 -2202
rect 76404 -2204 77004 -2202
rect 112404 -2204 113004 -2202
rect 148404 -2204 149004 -2202
rect 184404 -2204 185004 -2202
rect 220404 -2204 221004 -2202
rect 256404 -2204 257004 -2202
rect 292404 -2204 293004 -2202
rect 328404 -2204 329004 -2202
rect 364404 -2204 365004 -2202
rect 400404 -2204 401004 -2202
rect 436404 -2204 437004 -2202
rect 472404 -2204 473004 -2202
rect 508404 -2204 509004 -2202
rect 544404 -2204 545004 -2202
rect 580404 -2204 581004 -2202
rect 587200 -2204 587800 -2202
rect -3876 -2226 587800 -2204
rect -3876 -2462 -3694 -2226
rect -3458 -2462 4586 -2226
rect 4822 -2462 40586 -2226
rect 40822 -2462 76586 -2226
rect 76822 -2462 112586 -2226
rect 112822 -2462 148586 -2226
rect 148822 -2462 184586 -2226
rect 184822 -2462 220586 -2226
rect 220822 -2462 256586 -2226
rect 256822 -2462 292586 -2226
rect 292822 -2462 328586 -2226
rect 328822 -2462 364586 -2226
rect 364822 -2462 400586 -2226
rect 400822 -2462 436586 -2226
rect 436822 -2462 472586 -2226
rect 472822 -2462 508586 -2226
rect 508822 -2462 544586 -2226
rect 544822 -2462 580586 -2226
rect 580822 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect -3876 -2546 587800 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 4586 -2546
rect 4822 -2782 40586 -2546
rect 40822 -2782 76586 -2546
rect 76822 -2782 112586 -2546
rect 112822 -2782 148586 -2546
rect 148822 -2782 184586 -2546
rect 184822 -2782 220586 -2546
rect 220822 -2782 256586 -2546
rect 256822 -2782 292586 -2546
rect 292822 -2782 328586 -2546
rect 328822 -2782 364586 -2546
rect 364822 -2782 400586 -2546
rect 400822 -2782 436586 -2546
rect 436822 -2782 472586 -2546
rect 472822 -2782 508586 -2546
rect 508822 -2782 544586 -2546
rect 544822 -2782 580586 -2546
rect 580822 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect -3876 -2804 587800 -2782
rect -3876 -2806 -3276 -2804
rect 4404 -2806 5004 -2804
rect 40404 -2806 41004 -2804
rect 76404 -2806 77004 -2804
rect 112404 -2806 113004 -2804
rect 148404 -2806 149004 -2804
rect 184404 -2806 185004 -2804
rect 220404 -2806 221004 -2804
rect 256404 -2806 257004 -2804
rect 292404 -2806 293004 -2804
rect 328404 -2806 329004 -2804
rect 364404 -2806 365004 -2804
rect 400404 -2806 401004 -2804
rect 436404 -2806 437004 -2804
rect 472404 -2806 473004 -2804
rect 508404 -2806 509004 -2804
rect 544404 -2806 545004 -2804
rect 580404 -2806 581004 -2804
rect 587200 -2806 587800 -2804
rect -4816 -3144 -4216 -3142
rect 22404 -3144 23004 -3142
rect 58404 -3144 59004 -3142
rect 94404 -3144 95004 -3142
rect 130404 -3144 131004 -3142
rect 166404 -3144 167004 -3142
rect 202404 -3144 203004 -3142
rect 238404 -3144 239004 -3142
rect 274404 -3144 275004 -3142
rect 310404 -3144 311004 -3142
rect 346404 -3144 347004 -3142
rect 382404 -3144 383004 -3142
rect 418404 -3144 419004 -3142
rect 454404 -3144 455004 -3142
rect 490404 -3144 491004 -3142
rect 526404 -3144 527004 -3142
rect 562404 -3144 563004 -3142
rect 588140 -3144 588740 -3142
rect -4816 -3166 588740 -3144
rect -4816 -3402 -4634 -3166
rect -4398 -3402 22586 -3166
rect 22822 -3402 58586 -3166
rect 58822 -3402 94586 -3166
rect 94822 -3402 130586 -3166
rect 130822 -3402 166586 -3166
rect 166822 -3402 202586 -3166
rect 202822 -3402 238586 -3166
rect 238822 -3402 274586 -3166
rect 274822 -3402 310586 -3166
rect 310822 -3402 346586 -3166
rect 346822 -3402 382586 -3166
rect 382822 -3402 418586 -3166
rect 418822 -3402 454586 -3166
rect 454822 -3402 490586 -3166
rect 490822 -3402 526586 -3166
rect 526822 -3402 562586 -3166
rect 562822 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect -4816 -3486 588740 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 22586 -3486
rect 22822 -3722 58586 -3486
rect 58822 -3722 94586 -3486
rect 94822 -3722 130586 -3486
rect 130822 -3722 166586 -3486
rect 166822 -3722 202586 -3486
rect 202822 -3722 238586 -3486
rect 238822 -3722 274586 -3486
rect 274822 -3722 310586 -3486
rect 310822 -3722 346586 -3486
rect 346822 -3722 382586 -3486
rect 382822 -3722 418586 -3486
rect 418822 -3722 454586 -3486
rect 454822 -3722 490586 -3486
rect 490822 -3722 526586 -3486
rect 526822 -3722 562586 -3486
rect 562822 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect -4816 -3744 588740 -3722
rect -4816 -3746 -4216 -3744
rect 22404 -3746 23004 -3744
rect 58404 -3746 59004 -3744
rect 94404 -3746 95004 -3744
rect 130404 -3746 131004 -3744
rect 166404 -3746 167004 -3744
rect 202404 -3746 203004 -3744
rect 238404 -3746 239004 -3744
rect 274404 -3746 275004 -3744
rect 310404 -3746 311004 -3744
rect 346404 -3746 347004 -3744
rect 382404 -3746 383004 -3744
rect 418404 -3746 419004 -3744
rect 454404 -3746 455004 -3744
rect 490404 -3746 491004 -3744
rect 526404 -3746 527004 -3744
rect 562404 -3746 563004 -3744
rect 588140 -3746 588740 -3744
rect -5756 -4084 -5156 -4082
rect 8004 -4084 8604 -4082
rect 44004 -4084 44604 -4082
rect 80004 -4084 80604 -4082
rect 116004 -4084 116604 -4082
rect 152004 -4084 152604 -4082
rect 188004 -4084 188604 -4082
rect 224004 -4084 224604 -4082
rect 260004 -4084 260604 -4082
rect 296004 -4084 296604 -4082
rect 332004 -4084 332604 -4082
rect 368004 -4084 368604 -4082
rect 404004 -4084 404604 -4082
rect 440004 -4084 440604 -4082
rect 476004 -4084 476604 -4082
rect 512004 -4084 512604 -4082
rect 548004 -4084 548604 -4082
rect 589080 -4084 589680 -4082
rect -5756 -4106 589680 -4084
rect -5756 -4342 -5574 -4106
rect -5338 -4342 8186 -4106
rect 8422 -4342 44186 -4106
rect 44422 -4342 80186 -4106
rect 80422 -4342 116186 -4106
rect 116422 -4342 152186 -4106
rect 152422 -4342 188186 -4106
rect 188422 -4342 224186 -4106
rect 224422 -4342 260186 -4106
rect 260422 -4342 296186 -4106
rect 296422 -4342 332186 -4106
rect 332422 -4342 368186 -4106
rect 368422 -4342 404186 -4106
rect 404422 -4342 440186 -4106
rect 440422 -4342 476186 -4106
rect 476422 -4342 512186 -4106
rect 512422 -4342 548186 -4106
rect 548422 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect -5756 -4426 589680 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 8186 -4426
rect 8422 -4662 44186 -4426
rect 44422 -4662 80186 -4426
rect 80422 -4662 116186 -4426
rect 116422 -4662 152186 -4426
rect 152422 -4662 188186 -4426
rect 188422 -4662 224186 -4426
rect 224422 -4662 260186 -4426
rect 260422 -4662 296186 -4426
rect 296422 -4662 332186 -4426
rect 332422 -4662 368186 -4426
rect 368422 -4662 404186 -4426
rect 404422 -4662 440186 -4426
rect 440422 -4662 476186 -4426
rect 476422 -4662 512186 -4426
rect 512422 -4662 548186 -4426
rect 548422 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect -5756 -4684 589680 -4662
rect -5756 -4686 -5156 -4684
rect 8004 -4686 8604 -4684
rect 44004 -4686 44604 -4684
rect 80004 -4686 80604 -4684
rect 116004 -4686 116604 -4684
rect 152004 -4686 152604 -4684
rect 188004 -4686 188604 -4684
rect 224004 -4686 224604 -4684
rect 260004 -4686 260604 -4684
rect 296004 -4686 296604 -4684
rect 332004 -4686 332604 -4684
rect 368004 -4686 368604 -4684
rect 404004 -4686 404604 -4684
rect 440004 -4686 440604 -4684
rect 476004 -4686 476604 -4684
rect 512004 -4686 512604 -4684
rect 548004 -4686 548604 -4684
rect 589080 -4686 589680 -4684
rect -6696 -5024 -6096 -5022
rect 26004 -5024 26604 -5022
rect 62004 -5024 62604 -5022
rect 98004 -5024 98604 -5022
rect 134004 -5024 134604 -5022
rect 170004 -5024 170604 -5022
rect 206004 -5024 206604 -5022
rect 242004 -5024 242604 -5022
rect 278004 -5024 278604 -5022
rect 314004 -5024 314604 -5022
rect 350004 -5024 350604 -5022
rect 386004 -5024 386604 -5022
rect 422004 -5024 422604 -5022
rect 458004 -5024 458604 -5022
rect 494004 -5024 494604 -5022
rect 530004 -5024 530604 -5022
rect 566004 -5024 566604 -5022
rect 590020 -5024 590620 -5022
rect -6696 -5046 590620 -5024
rect -6696 -5282 -6514 -5046
rect -6278 -5282 26186 -5046
rect 26422 -5282 62186 -5046
rect 62422 -5282 98186 -5046
rect 98422 -5282 134186 -5046
rect 134422 -5282 170186 -5046
rect 170422 -5282 206186 -5046
rect 206422 -5282 242186 -5046
rect 242422 -5282 278186 -5046
rect 278422 -5282 314186 -5046
rect 314422 -5282 350186 -5046
rect 350422 -5282 386186 -5046
rect 386422 -5282 422186 -5046
rect 422422 -5282 458186 -5046
rect 458422 -5282 494186 -5046
rect 494422 -5282 530186 -5046
rect 530422 -5282 566186 -5046
rect 566422 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect -6696 -5366 590620 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 26186 -5366
rect 26422 -5602 62186 -5366
rect 62422 -5602 98186 -5366
rect 98422 -5602 134186 -5366
rect 134422 -5602 170186 -5366
rect 170422 -5602 206186 -5366
rect 206422 -5602 242186 -5366
rect 242422 -5602 278186 -5366
rect 278422 -5602 314186 -5366
rect 314422 -5602 350186 -5366
rect 350422 -5602 386186 -5366
rect 386422 -5602 422186 -5366
rect 422422 -5602 458186 -5366
rect 458422 -5602 494186 -5366
rect 494422 -5602 530186 -5366
rect 530422 -5602 566186 -5366
rect 566422 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect -6696 -5624 590620 -5602
rect -6696 -5626 -6096 -5624
rect 26004 -5626 26604 -5624
rect 62004 -5626 62604 -5624
rect 98004 -5626 98604 -5624
rect 134004 -5626 134604 -5624
rect 170004 -5626 170604 -5624
rect 206004 -5626 206604 -5624
rect 242004 -5626 242604 -5624
rect 278004 -5626 278604 -5624
rect 314004 -5626 314604 -5624
rect 350004 -5626 350604 -5624
rect 386004 -5626 386604 -5624
rect 422004 -5626 422604 -5624
rect 458004 -5626 458604 -5624
rect 494004 -5626 494604 -5624
rect 530004 -5626 530604 -5624
rect 566004 -5626 566604 -5624
rect 590020 -5626 590620 -5624
rect -7636 -5964 -7036 -5962
rect 11604 -5964 12204 -5962
rect 47604 -5964 48204 -5962
rect 83604 -5964 84204 -5962
rect 119604 -5964 120204 -5962
rect 155604 -5964 156204 -5962
rect 191604 -5964 192204 -5962
rect 227604 -5964 228204 -5962
rect 263604 -5964 264204 -5962
rect 299604 -5964 300204 -5962
rect 335604 -5964 336204 -5962
rect 371604 -5964 372204 -5962
rect 407604 -5964 408204 -5962
rect 443604 -5964 444204 -5962
rect 479604 -5964 480204 -5962
rect 515604 -5964 516204 -5962
rect 551604 -5964 552204 -5962
rect 590960 -5964 591560 -5962
rect -7636 -5986 591560 -5964
rect -7636 -6222 -7454 -5986
rect -7218 -6222 11786 -5986
rect 12022 -6222 47786 -5986
rect 48022 -6222 83786 -5986
rect 84022 -6222 119786 -5986
rect 120022 -6222 155786 -5986
rect 156022 -6222 191786 -5986
rect 192022 -6222 227786 -5986
rect 228022 -6222 263786 -5986
rect 264022 -6222 299786 -5986
rect 300022 -6222 335786 -5986
rect 336022 -6222 371786 -5986
rect 372022 -6222 407786 -5986
rect 408022 -6222 443786 -5986
rect 444022 -6222 479786 -5986
rect 480022 -6222 515786 -5986
rect 516022 -6222 551786 -5986
rect 552022 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect -7636 -6306 591560 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 11786 -6306
rect 12022 -6542 47786 -6306
rect 48022 -6542 83786 -6306
rect 84022 -6542 119786 -6306
rect 120022 -6542 155786 -6306
rect 156022 -6542 191786 -6306
rect 192022 -6542 227786 -6306
rect 228022 -6542 263786 -6306
rect 264022 -6542 299786 -6306
rect 300022 -6542 335786 -6306
rect 336022 -6542 371786 -6306
rect 372022 -6542 407786 -6306
rect 408022 -6542 443786 -6306
rect 444022 -6542 479786 -6306
rect 480022 -6542 515786 -6306
rect 516022 -6542 551786 -6306
rect 552022 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect -7636 -6564 591560 -6542
rect -7636 -6566 -7036 -6564
rect 11604 -6566 12204 -6564
rect 47604 -6566 48204 -6564
rect 83604 -6566 84204 -6564
rect 119604 -6566 120204 -6564
rect 155604 -6566 156204 -6564
rect 191604 -6566 192204 -6564
rect 227604 -6566 228204 -6564
rect 263604 -6566 264204 -6564
rect 299604 -6566 300204 -6564
rect 335604 -6566 336204 -6564
rect 371604 -6566 372204 -6564
rect 407604 -6566 408204 -6564
rect 443604 -6566 444204 -6564
rect 479604 -6566 480204 -6564
rect 515604 -6566 516204 -6564
rect 551604 -6566 552204 -6564
rect 590960 -6566 591560 -6564
rect -8576 -6904 -7976 -6902
rect 29604 -6904 30204 -6902
rect 65604 -6904 66204 -6902
rect 101604 -6904 102204 -6902
rect 137604 -6904 138204 -6902
rect 173604 -6904 174204 -6902
rect 209604 -6904 210204 -6902
rect 245604 -6904 246204 -6902
rect 281604 -6904 282204 -6902
rect 317604 -6904 318204 -6902
rect 353604 -6904 354204 -6902
rect 389604 -6904 390204 -6902
rect 425604 -6904 426204 -6902
rect 461604 -6904 462204 -6902
rect 497604 -6904 498204 -6902
rect 533604 -6904 534204 -6902
rect 569604 -6904 570204 -6902
rect 591900 -6904 592500 -6902
rect -8576 -6926 592500 -6904
rect -8576 -7162 -8394 -6926
rect -8158 -7162 29786 -6926
rect 30022 -7162 65786 -6926
rect 66022 -7162 101786 -6926
rect 102022 -7162 137786 -6926
rect 138022 -7162 173786 -6926
rect 174022 -7162 209786 -6926
rect 210022 -7162 245786 -6926
rect 246022 -7162 281786 -6926
rect 282022 -7162 317786 -6926
rect 318022 -7162 353786 -6926
rect 354022 -7162 389786 -6926
rect 390022 -7162 425786 -6926
rect 426022 -7162 461786 -6926
rect 462022 -7162 497786 -6926
rect 498022 -7162 533786 -6926
rect 534022 -7162 569786 -6926
rect 570022 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect -8576 -7246 592500 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 29786 -7246
rect 30022 -7482 65786 -7246
rect 66022 -7482 101786 -7246
rect 102022 -7482 137786 -7246
rect 138022 -7482 173786 -7246
rect 174022 -7482 209786 -7246
rect 210022 -7482 245786 -7246
rect 246022 -7482 281786 -7246
rect 282022 -7482 317786 -7246
rect 318022 -7482 353786 -7246
rect 354022 -7482 389786 -7246
rect 390022 -7482 425786 -7246
rect 426022 -7482 461786 -7246
rect 462022 -7482 497786 -7246
rect 498022 -7482 533786 -7246
rect 534022 -7482 569786 -7246
rect 570022 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect -8576 -7504 592500 -7482
rect -8576 -7506 -7976 -7504
rect 29604 -7506 30204 -7504
rect 65604 -7506 66204 -7504
rect 101604 -7506 102204 -7504
rect 137604 -7506 138204 -7504
rect 173604 -7506 174204 -7504
rect 209604 -7506 210204 -7504
rect 245604 -7506 246204 -7504
rect 281604 -7506 282204 -7504
rect 317604 -7506 318204 -7504
rect 353604 -7506 354204 -7504
rect 389604 -7506 390204 -7504
rect 425604 -7506 426204 -7504
rect 461604 -7506 462204 -7504
rect 497604 -7506 498204 -7504
rect 533604 -7506 534204 -7504
rect 569604 -7506 570204 -7504
rect 591900 -7506 592500 -7504
use user_proj_example  mprj
timestamp 1610260563
transform 1 0 8000 0 1 8000
box 0 0 568000 688000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew signal bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew signal bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew signal bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew signal bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew signal input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew signal input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew signal input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew signal input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew signal input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew signal input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew signal input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew signal input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew signal input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew signal input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew signal input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew signal input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew signal input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew signal input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew signal input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew signal input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew signal input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew signal input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew signal input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew signal input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew signal input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew signal input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew signal input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew signal input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew signal input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew signal input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew signal input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew signal input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew signal input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew signal tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew signal tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew signal tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew signal tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew signal tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew signal tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew signal tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew signal tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew signal tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew signal tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew signal tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew signal tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew signal tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew signal tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew signal tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew signal tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew signal tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew signal tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew signal tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew signal tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew signal tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew signal tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew signal tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew signal tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew signal tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew signal tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew signal tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew signal tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew signal tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew signal tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew signal tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew signal tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew signal tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew signal tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew signal tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew signal tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew signal tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew signal tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew signal tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew signal tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew signal tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew signal tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew signal tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew signal tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew signal tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew signal tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew signal tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew signal tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew signal tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew signal tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew signal tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew signal tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew signal tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew signal tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew signal tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew signal tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew signal tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew signal tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew signal input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew signal input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew signal input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew signal input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew signal input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew signal input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew signal input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew signal input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew signal input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew signal input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew signal input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew signal input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew signal input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew signal input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew signal input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew signal input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew signal input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew signal input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew signal input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew signal input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew signal input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew signal input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew signal input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew signal input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew signal input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew signal input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew signal input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew signal input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew signal input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew signal input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew signal input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew signal input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew signal input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew signal input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew signal input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew signal input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew signal input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew signal input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew signal input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew signal input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew signal input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew signal input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew signal input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew signal input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew signal input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew signal input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew signal input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew signal input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew signal input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew signal input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew signal input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew signal input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew signal input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew signal input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew signal input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew signal input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew signal input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew signal input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew signal input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew signal input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew signal input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew signal input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew signal input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew signal input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew signal input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew signal input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew signal input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew signal input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew signal input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew signal input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew signal input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew signal input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew signal input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew signal input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew signal input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew signal input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew signal input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew signal input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew signal input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew signal input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew signal input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew signal input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew signal input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew signal input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew signal input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew signal input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew signal input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew signal input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew signal input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew signal input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew signal input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew signal input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew signal input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew signal input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew signal input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew signal input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew signal input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew signal input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew signal input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew signal input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew signal input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew signal input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew signal input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew signal input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew signal input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew signal input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew signal input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew signal input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew signal input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew signal input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew signal input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew signal input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew signal input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew signal input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew signal input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew signal input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew signal input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew signal input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew signal input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew signal input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew signal input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew signal input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew signal tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew signal tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew signal tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew signal tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew signal tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew signal tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew signal tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew signal tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew signal tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew signal tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew signal tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew signal tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew signal tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew signal tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew signal tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew signal tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew signal tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew signal tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew signal tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew signal tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew signal tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew signal tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew signal tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew signal tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew signal tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew signal tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew signal tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew signal tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew signal tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew signal tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew signal tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew signal tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew signal tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew signal tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew signal tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew signal tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew signal tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew signal tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew signal tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew signal tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew signal tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew signal tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew signal tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew signal tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew signal tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew signal tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew signal tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew signal tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew signal tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew signal tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew signal tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew signal tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew signal tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew signal tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew signal tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew signal tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew signal tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew signal tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew signal tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew signal tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew signal tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew signal tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew signal tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew signal tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew signal tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew signal tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew signal tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew signal tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew signal tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew signal tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew signal tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew signal tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew signal tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew signal tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew signal tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew signal tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew signal tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew signal tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew signal tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew signal tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew signal tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew signal tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew signal tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew signal tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew signal tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew signal tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew signal tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew signal tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew signal tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew signal tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew signal tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew signal tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew signal tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew signal tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew signal tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew signal tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew signal tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew signal tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew signal tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew signal tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew signal tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew signal tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew signal tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew signal tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew signal tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew signal tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew signal tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew signal tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew signal tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew signal tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew signal tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew signal tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew signal tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew signal tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew signal tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew signal tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew signal tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew signal tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew signal tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew signal tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew signal tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew signal tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew signal tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew signal tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew signal tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew signal tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew signal tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew signal input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew signal input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew signal input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew signal input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew signal input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew signal input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew signal input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew signal input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew signal input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew signal input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew signal input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew signal input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew signal input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew signal input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew signal input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew signal input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew signal input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew signal input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew signal input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew signal input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew signal input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew signal input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew signal input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew signal input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew signal input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew signal input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew signal input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew signal input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew signal input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew signal input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew signal input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew signal input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew signal input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew signal input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew signal input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew signal input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew signal input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew signal input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew signal input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew signal input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew signal input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew signal input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew signal input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew signal input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew signal input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew signal input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew signal input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew signal input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew signal input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew signal input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew signal input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew signal input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew signal input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew signal input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew signal input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew signal input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew signal input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew signal input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew signal input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew signal input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew signal input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew signal input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew signal input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew signal input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew signal input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew signal input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew signal input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew signal input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew signal input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew signal input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew signal input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew signal input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew signal input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew signal input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew signal input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew signal input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew signal input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew signal input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew signal input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew signal input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew signal input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew signal input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew signal input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew signal input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew signal input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew signal input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew signal input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew signal input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew signal input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew signal input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew signal input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew signal input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew signal input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew signal input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew signal input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew signal input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew signal input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew signal input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew signal input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew signal input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew signal input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew signal input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew signal input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew signal input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew signal input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew signal input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew signal input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew signal input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew signal input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew signal input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew signal input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew signal input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew signal input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew signal input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew signal input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew signal input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew signal input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew signal input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew signal input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew signal input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew signal input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew signal input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew signal input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew signal input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew signal input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew signal input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew signal input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew signal input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew signal input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew signal input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew signal input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew signal input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew signal input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew signal input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew signal input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew signal input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew signal input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew signal input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew signal input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew signal input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew signal input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew signal input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew signal input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew signal input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew signal input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew signal input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew signal input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew signal input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew signal input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew signal input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew signal input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew signal input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew signal input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew signal input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew signal input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew signal input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew signal input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew signal input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew signal input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew signal input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew signal input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew signal input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew signal input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew signal input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew signal input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew signal input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew signal input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew signal input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew signal input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew signal input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew signal input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew signal input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew signal input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew signal input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew signal input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew signal input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew signal input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew signal input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew signal input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew signal input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew signal input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew signal input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew signal input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew signal input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew signal input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew signal input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew signal input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew signal input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew signal tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew signal tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew signal tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew signal tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew signal tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew signal tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew signal tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew signal tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew signal tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew signal tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew signal tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew signal tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew signal tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew signal tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew signal tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew signal tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew signal tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew signal tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew signal tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew signal tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew signal tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew signal tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew signal tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew signal tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew signal tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew signal tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew signal tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew signal tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew signal tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew signal tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew signal tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew signal tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew signal input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew signal input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew signal input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew signal input
rlabel metal4 s 576804 697952 577404 705800 6 vccd1
port 636 nsew power bidirectional
rlabel metal4 s 540804 697952 541404 705800 6 vccd1
port 637 nsew power bidirectional
rlabel metal4 s 504804 697952 505404 705800 6 vccd1
port 638 nsew power bidirectional
rlabel metal4 s 468804 697952 469404 705800 6 vccd1
port 639 nsew power bidirectional
rlabel metal4 s 432804 697952 433404 705800 6 vccd1
port 640 nsew power bidirectional
rlabel metal4 s 396804 697952 397404 705800 6 vccd1
port 641 nsew power bidirectional
rlabel metal4 s 360804 697952 361404 705800 6 vccd1
port 642 nsew power bidirectional
rlabel metal4 s 324804 697952 325404 705800 6 vccd1
port 643 nsew power bidirectional
rlabel metal4 s 288804 697952 289404 705800 6 vccd1
port 644 nsew power bidirectional
rlabel metal4 s 252804 697952 253404 705800 6 vccd1
port 645 nsew power bidirectional
rlabel metal4 s 216804 697952 217404 705800 6 vccd1
port 646 nsew power bidirectional
rlabel metal4 s 180804 697952 181404 705800 6 vccd1
port 647 nsew power bidirectional
rlabel metal4 s 144804 697952 145404 705800 6 vccd1
port 648 nsew power bidirectional
rlabel metal4 s 108804 697952 109404 705800 6 vccd1
port 649 nsew power bidirectional
rlabel metal4 s 72804 697952 73404 705800 6 vccd1
port 650 nsew power bidirectional
rlabel metal4 s 36804 697952 37404 705800 6 vccd1
port 651 nsew power bidirectional
rlabel metal4 s 804 -1864 1404 705800 6 vccd1
port 652 nsew power bidirectional
rlabel metal4 s 585320 -924 585920 704860 6 vccd1
port 653 nsew power bidirectional
rlabel metal4 s -1996 -924 -1396 704860 4 vccd1
port 654 nsew power bidirectional
rlabel metal4 s 576804 -1864 577404 6048 6 vccd1
port 655 nsew power bidirectional
rlabel metal4 s 540804 -1864 541404 6048 6 vccd1
port 656 nsew power bidirectional
rlabel metal4 s 504804 -1864 505404 6048 6 vccd1
port 657 nsew power bidirectional
rlabel metal4 s 468804 -1864 469404 6048 6 vccd1
port 658 nsew power bidirectional
rlabel metal4 s 432804 -1864 433404 6048 6 vccd1
port 659 nsew power bidirectional
rlabel metal4 s 396804 -1864 397404 6048 6 vccd1
port 660 nsew power bidirectional
rlabel metal4 s 360804 -1864 361404 6048 6 vccd1
port 661 nsew power bidirectional
rlabel metal4 s 324804 -1864 325404 6048 6 vccd1
port 662 nsew power bidirectional
rlabel metal4 s 288804 -1864 289404 6048 6 vccd1
port 663 nsew power bidirectional
rlabel metal4 s 252804 -1864 253404 6048 6 vccd1
port 664 nsew power bidirectional
rlabel metal4 s 216804 -1864 217404 6048 6 vccd1
port 665 nsew power bidirectional
rlabel metal4 s 180804 -1864 181404 6048 6 vccd1
port 666 nsew power bidirectional
rlabel metal4 s 144804 -1864 145404 6048 6 vccd1
port 667 nsew power bidirectional
rlabel metal4 s 108804 -1864 109404 6048 6 vccd1
port 668 nsew power bidirectional
rlabel metal4 s 72804 -1864 73404 6048 6 vccd1
port 669 nsew power bidirectional
rlabel metal4 s 36804 -1864 37404 6048 6 vccd1
port 670 nsew power bidirectional
rlabel metal5 s -1996 704260 585920 704860 6 vccd1
port 671 nsew power bidirectional
rlabel metal5 s -2936 685828 586860 686428 6 vccd1
port 672 nsew power bidirectional
rlabel metal5 s -2936 649828 586860 650428 6 vccd1
port 673 nsew power bidirectional
rlabel metal5 s -2936 613828 586860 614428 6 vccd1
port 674 nsew power bidirectional
rlabel metal5 s -2936 577828 586860 578428 6 vccd1
port 675 nsew power bidirectional
rlabel metal5 s -2936 541828 586860 542428 6 vccd1
port 676 nsew power bidirectional
rlabel metal5 s -2936 505828 586860 506428 6 vccd1
port 677 nsew power bidirectional
rlabel metal5 s -2936 469828 586860 470428 6 vccd1
port 678 nsew power bidirectional
rlabel metal5 s -2936 433828 586860 434428 6 vccd1
port 679 nsew power bidirectional
rlabel metal5 s -2936 397828 586860 398428 6 vccd1
port 680 nsew power bidirectional
rlabel metal5 s -2936 361828 586860 362428 6 vccd1
port 681 nsew power bidirectional
rlabel metal5 s -2936 325828 586860 326428 6 vccd1
port 682 nsew power bidirectional
rlabel metal5 s -2936 289828 586860 290428 6 vccd1
port 683 nsew power bidirectional
rlabel metal5 s -2936 253828 586860 254428 6 vccd1
port 684 nsew power bidirectional
rlabel metal5 s -2936 217828 586860 218428 6 vccd1
port 685 nsew power bidirectional
rlabel metal5 s -2936 181828 586860 182428 6 vccd1
port 686 nsew power bidirectional
rlabel metal5 s -2936 145828 586860 146428 6 vccd1
port 687 nsew power bidirectional
rlabel metal5 s -2936 109828 586860 110428 6 vccd1
port 688 nsew power bidirectional
rlabel metal5 s -2936 73828 586860 74428 6 vccd1
port 689 nsew power bidirectional
rlabel metal5 s -2936 37828 586860 38428 6 vccd1
port 690 nsew power bidirectional
rlabel metal5 s -2936 1828 586860 2428 6 vccd1
port 691 nsew power bidirectional
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 692 nsew power bidirectional
rlabel metal4 s 586260 -1864 586860 705800 6 vssd1
port 693 nsew ground bidirectional
rlabel metal4 s 558804 697952 559404 705800 6 vssd1
port 694 nsew ground bidirectional
rlabel metal4 s 522804 697952 523404 705800 6 vssd1
port 695 nsew ground bidirectional
rlabel metal4 s 486804 697952 487404 705800 6 vssd1
port 696 nsew ground bidirectional
rlabel metal4 s 450804 697952 451404 705800 6 vssd1
port 697 nsew ground bidirectional
rlabel metal4 s 414804 697952 415404 705800 6 vssd1
port 698 nsew ground bidirectional
rlabel metal4 s 378804 697952 379404 705800 6 vssd1
port 699 nsew ground bidirectional
rlabel metal4 s 342804 697952 343404 705800 6 vssd1
port 700 nsew ground bidirectional
rlabel metal4 s 306804 697952 307404 705800 6 vssd1
port 701 nsew ground bidirectional
rlabel metal4 s 270804 697952 271404 705800 6 vssd1
port 702 nsew ground bidirectional
rlabel metal4 s 234804 697952 235404 705800 6 vssd1
port 703 nsew ground bidirectional
rlabel metal4 s 198804 697952 199404 705800 6 vssd1
port 704 nsew ground bidirectional
rlabel metal4 s 162804 697952 163404 705800 6 vssd1
port 705 nsew ground bidirectional
rlabel metal4 s 126804 697952 127404 705800 6 vssd1
port 706 nsew ground bidirectional
rlabel metal4 s 90804 697952 91404 705800 6 vssd1
port 707 nsew ground bidirectional
rlabel metal4 s 54804 697952 55404 705800 6 vssd1
port 708 nsew ground bidirectional
rlabel metal4 s 18804 697952 19404 705800 6 vssd1
port 709 nsew ground bidirectional
rlabel metal4 s -2936 -1864 -2336 705800 4 vssd1
port 710 nsew ground bidirectional
rlabel metal4 s 558804 -1864 559404 6048 6 vssd1
port 711 nsew ground bidirectional
rlabel metal4 s 522804 -1864 523404 6048 6 vssd1
port 712 nsew ground bidirectional
rlabel metal4 s 486804 -1864 487404 6048 6 vssd1
port 713 nsew ground bidirectional
rlabel metal4 s 450804 -1864 451404 6048 6 vssd1
port 714 nsew ground bidirectional
rlabel metal4 s 414804 -1864 415404 6048 6 vssd1
port 715 nsew ground bidirectional
rlabel metal4 s 378804 -1864 379404 6048 6 vssd1
port 716 nsew ground bidirectional
rlabel metal4 s 342804 -1864 343404 6048 6 vssd1
port 717 nsew ground bidirectional
rlabel metal4 s 306804 -1864 307404 6048 6 vssd1
port 718 nsew ground bidirectional
rlabel metal4 s 270804 -1864 271404 6048 6 vssd1
port 719 nsew ground bidirectional
rlabel metal4 s 234804 -1864 235404 6048 6 vssd1
port 720 nsew ground bidirectional
rlabel metal4 s 198804 -1864 199404 6048 6 vssd1
port 721 nsew ground bidirectional
rlabel metal4 s 162804 -1864 163404 6048 6 vssd1
port 722 nsew ground bidirectional
rlabel metal4 s 126804 -1864 127404 6048 6 vssd1
port 723 nsew ground bidirectional
rlabel metal4 s 90804 -1864 91404 6048 6 vssd1
port 724 nsew ground bidirectional
rlabel metal4 s 54804 -1864 55404 6048 6 vssd1
port 725 nsew ground bidirectional
rlabel metal4 s 18804 -1864 19404 6048 6 vssd1
port 726 nsew ground bidirectional
rlabel metal5 s -2936 705200 586860 705800 6 vssd1
port 727 nsew ground bidirectional
rlabel metal5 s -2936 667828 586860 668428 6 vssd1
port 728 nsew ground bidirectional
rlabel metal5 s -2936 631828 586860 632428 6 vssd1
port 729 nsew ground bidirectional
rlabel metal5 s -2936 595828 586860 596428 6 vssd1
port 730 nsew ground bidirectional
rlabel metal5 s -2936 559828 586860 560428 6 vssd1
port 731 nsew ground bidirectional
rlabel metal5 s -2936 523828 586860 524428 6 vssd1
port 732 nsew ground bidirectional
rlabel metal5 s -2936 487828 586860 488428 6 vssd1
port 733 nsew ground bidirectional
rlabel metal5 s -2936 451828 586860 452428 6 vssd1
port 734 nsew ground bidirectional
rlabel metal5 s -2936 415828 586860 416428 6 vssd1
port 735 nsew ground bidirectional
rlabel metal5 s -2936 379828 586860 380428 6 vssd1
port 736 nsew ground bidirectional
rlabel metal5 s -2936 343828 586860 344428 6 vssd1
port 737 nsew ground bidirectional
rlabel metal5 s -2936 307828 586860 308428 6 vssd1
port 738 nsew ground bidirectional
rlabel metal5 s -2936 271828 586860 272428 6 vssd1
port 739 nsew ground bidirectional
rlabel metal5 s -2936 235828 586860 236428 6 vssd1
port 740 nsew ground bidirectional
rlabel metal5 s -2936 199828 586860 200428 6 vssd1
port 741 nsew ground bidirectional
rlabel metal5 s -2936 163828 586860 164428 6 vssd1
port 742 nsew ground bidirectional
rlabel metal5 s -2936 127828 586860 128428 6 vssd1
port 743 nsew ground bidirectional
rlabel metal5 s -2936 91828 586860 92428 6 vssd1
port 744 nsew ground bidirectional
rlabel metal5 s -2936 55828 586860 56428 6 vssd1
port 745 nsew ground bidirectional
rlabel metal5 s -2936 19828 586860 20428 6 vssd1
port 746 nsew ground bidirectional
rlabel metal5 s -2936 -1864 586860 -1264 8 vssd1
port 747 nsew ground bidirectional
rlabel metal4 s 580404 -3744 581004 707680 6 vccd2
port 748 nsew power bidirectional
rlabel metal4 s 544404 698000 545004 707680 6 vccd2
port 749 nsew power bidirectional
rlabel metal4 s 508404 698000 509004 707680 6 vccd2
port 750 nsew power bidirectional
rlabel metal4 s 472404 698000 473004 707680 6 vccd2
port 751 nsew power bidirectional
rlabel metal4 s 436404 698000 437004 707680 6 vccd2
port 752 nsew power bidirectional
rlabel metal4 s 400404 698000 401004 707680 6 vccd2
port 753 nsew power bidirectional
rlabel metal4 s 364404 698000 365004 707680 6 vccd2
port 754 nsew power bidirectional
rlabel metal4 s 328404 698000 329004 707680 6 vccd2
port 755 nsew power bidirectional
rlabel metal4 s 292404 698000 293004 707680 6 vccd2
port 756 nsew power bidirectional
rlabel metal4 s 256404 698000 257004 707680 6 vccd2
port 757 nsew power bidirectional
rlabel metal4 s 220404 698000 221004 707680 6 vccd2
port 758 nsew power bidirectional
rlabel metal4 s 184404 698000 185004 707680 6 vccd2
port 759 nsew power bidirectional
rlabel metal4 s 148404 698000 149004 707680 6 vccd2
port 760 nsew power bidirectional
rlabel metal4 s 112404 698000 113004 707680 6 vccd2
port 761 nsew power bidirectional
rlabel metal4 s 76404 698000 77004 707680 6 vccd2
port 762 nsew power bidirectional
rlabel metal4 s 40404 698000 41004 707680 6 vccd2
port 763 nsew power bidirectional
rlabel metal4 s 4404 -3744 5004 707680 6 vccd2
port 764 nsew power bidirectional
rlabel metal4 s 587200 -2804 587800 706740 6 vccd2
port 765 nsew power bidirectional
rlabel metal4 s -3876 -2804 -3276 706740 4 vccd2
port 766 nsew power bidirectional
rlabel metal4 s 544404 -3744 545004 6000 6 vccd2
port 767 nsew power bidirectional
rlabel metal4 s 508404 -3744 509004 6000 6 vccd2
port 768 nsew power bidirectional
rlabel metal4 s 472404 -3744 473004 6000 6 vccd2
port 769 nsew power bidirectional
rlabel metal4 s 436404 -3744 437004 6000 6 vccd2
port 770 nsew power bidirectional
rlabel metal4 s 400404 -3744 401004 6000 6 vccd2
port 771 nsew power bidirectional
rlabel metal4 s 364404 -3744 365004 6000 6 vccd2
port 772 nsew power bidirectional
rlabel metal4 s 328404 -3744 329004 6000 6 vccd2
port 773 nsew power bidirectional
rlabel metal4 s 292404 -3744 293004 6000 6 vccd2
port 774 nsew power bidirectional
rlabel metal4 s 256404 -3744 257004 6000 6 vccd2
port 775 nsew power bidirectional
rlabel metal4 s 220404 -3744 221004 6000 6 vccd2
port 776 nsew power bidirectional
rlabel metal4 s 184404 -3744 185004 6000 6 vccd2
port 777 nsew power bidirectional
rlabel metal4 s 148404 -3744 149004 6000 6 vccd2
port 778 nsew power bidirectional
rlabel metal4 s 112404 -3744 113004 6000 6 vccd2
port 779 nsew power bidirectional
rlabel metal4 s 76404 -3744 77004 6000 6 vccd2
port 780 nsew power bidirectional
rlabel metal4 s 40404 -3744 41004 6000 6 vccd2
port 781 nsew power bidirectional
rlabel metal5 s -3876 706140 587800 706740 6 vccd2
port 782 nsew power bidirectional
rlabel metal5 s -4816 689476 588740 690076 6 vccd2
port 783 nsew power bidirectional
rlabel metal5 s -4816 653476 588740 654076 6 vccd2
port 784 nsew power bidirectional
rlabel metal5 s -4816 617476 588740 618076 6 vccd2
port 785 nsew power bidirectional
rlabel metal5 s -4816 581476 588740 582076 6 vccd2
port 786 nsew power bidirectional
rlabel metal5 s -4816 545476 588740 546076 6 vccd2
port 787 nsew power bidirectional
rlabel metal5 s -4816 509476 588740 510076 6 vccd2
port 788 nsew power bidirectional
rlabel metal5 s -4816 473476 588740 474076 6 vccd2
port 789 nsew power bidirectional
rlabel metal5 s -4816 437476 588740 438076 6 vccd2
port 790 nsew power bidirectional
rlabel metal5 s -4816 401476 588740 402076 6 vccd2
port 791 nsew power bidirectional
rlabel metal5 s -4816 365476 588740 366076 6 vccd2
port 792 nsew power bidirectional
rlabel metal5 s -4816 329476 588740 330076 6 vccd2
port 793 nsew power bidirectional
rlabel metal5 s -4816 293476 588740 294076 6 vccd2
port 794 nsew power bidirectional
rlabel metal5 s -4816 257476 588740 258076 6 vccd2
port 795 nsew power bidirectional
rlabel metal5 s -4816 221476 588740 222076 6 vccd2
port 796 nsew power bidirectional
rlabel metal5 s -4816 185476 588740 186076 6 vccd2
port 797 nsew power bidirectional
rlabel metal5 s -4816 149476 588740 150076 6 vccd2
port 798 nsew power bidirectional
rlabel metal5 s -4816 113476 588740 114076 6 vccd2
port 799 nsew power bidirectional
rlabel metal5 s -4816 77476 588740 78076 6 vccd2
port 800 nsew power bidirectional
rlabel metal5 s -4816 41476 588740 42076 6 vccd2
port 801 nsew power bidirectional
rlabel metal5 s -4816 5476 588740 6076 6 vccd2
port 802 nsew power bidirectional
rlabel metal5 s -3876 -2804 587800 -2204 8 vccd2
port 803 nsew power bidirectional
rlabel metal4 s 588140 -3744 588740 707680 6 vssd2
port 804 nsew ground bidirectional
rlabel metal4 s 562404 698000 563004 707680 6 vssd2
port 805 nsew ground bidirectional
rlabel metal4 s 526404 698000 527004 707680 6 vssd2
port 806 nsew ground bidirectional
rlabel metal4 s 490404 698000 491004 707680 6 vssd2
port 807 nsew ground bidirectional
rlabel metal4 s 454404 698000 455004 707680 6 vssd2
port 808 nsew ground bidirectional
rlabel metal4 s 418404 698000 419004 707680 6 vssd2
port 809 nsew ground bidirectional
rlabel metal4 s 382404 698000 383004 707680 6 vssd2
port 810 nsew ground bidirectional
rlabel metal4 s 346404 698000 347004 707680 6 vssd2
port 811 nsew ground bidirectional
rlabel metal4 s 310404 698000 311004 707680 6 vssd2
port 812 nsew ground bidirectional
rlabel metal4 s 274404 698000 275004 707680 6 vssd2
port 813 nsew ground bidirectional
rlabel metal4 s 238404 698000 239004 707680 6 vssd2
port 814 nsew ground bidirectional
rlabel metal4 s 202404 698000 203004 707680 6 vssd2
port 815 nsew ground bidirectional
rlabel metal4 s 166404 698000 167004 707680 6 vssd2
port 816 nsew ground bidirectional
rlabel metal4 s 130404 698000 131004 707680 6 vssd2
port 817 nsew ground bidirectional
rlabel metal4 s 94404 698000 95004 707680 6 vssd2
port 818 nsew ground bidirectional
rlabel metal4 s 58404 698000 59004 707680 6 vssd2
port 819 nsew ground bidirectional
rlabel metal4 s 22404 698000 23004 707680 6 vssd2
port 820 nsew ground bidirectional
rlabel metal4 s -4816 -3744 -4216 707680 4 vssd2
port 821 nsew ground bidirectional
rlabel metal4 s 562404 -3744 563004 6000 6 vssd2
port 822 nsew ground bidirectional
rlabel metal4 s 526404 -3744 527004 6000 6 vssd2
port 823 nsew ground bidirectional
rlabel metal4 s 490404 -3744 491004 6000 6 vssd2
port 824 nsew ground bidirectional
rlabel metal4 s 454404 -3744 455004 6000 6 vssd2
port 825 nsew ground bidirectional
rlabel metal4 s 418404 -3744 419004 6000 6 vssd2
port 826 nsew ground bidirectional
rlabel metal4 s 382404 -3744 383004 6000 6 vssd2
port 827 nsew ground bidirectional
rlabel metal4 s 346404 -3744 347004 6000 6 vssd2
port 828 nsew ground bidirectional
rlabel metal4 s 310404 -3744 311004 6000 6 vssd2
port 829 nsew ground bidirectional
rlabel metal4 s 274404 -3744 275004 6000 6 vssd2
port 830 nsew ground bidirectional
rlabel metal4 s 238404 -3744 239004 6000 6 vssd2
port 831 nsew ground bidirectional
rlabel metal4 s 202404 -3744 203004 6000 6 vssd2
port 832 nsew ground bidirectional
rlabel metal4 s 166404 -3744 167004 6000 6 vssd2
port 833 nsew ground bidirectional
rlabel metal4 s 130404 -3744 131004 6000 6 vssd2
port 834 nsew ground bidirectional
rlabel metal4 s 94404 -3744 95004 6000 6 vssd2
port 835 nsew ground bidirectional
rlabel metal4 s 58404 -3744 59004 6000 6 vssd2
port 836 nsew ground bidirectional
rlabel metal4 s 22404 -3744 23004 6000 6 vssd2
port 837 nsew ground bidirectional
rlabel metal5 s -4816 707080 588740 707680 6 vssd2
port 838 nsew ground bidirectional
rlabel metal5 s -4816 671476 588740 672076 6 vssd2
port 839 nsew ground bidirectional
rlabel metal5 s -4816 635476 588740 636076 6 vssd2
port 840 nsew ground bidirectional
rlabel metal5 s -4816 599476 588740 600076 6 vssd2
port 841 nsew ground bidirectional
rlabel metal5 s -4816 563476 588740 564076 6 vssd2
port 842 nsew ground bidirectional
rlabel metal5 s -4816 527476 588740 528076 6 vssd2
port 843 nsew ground bidirectional
rlabel metal5 s -4816 491476 588740 492076 6 vssd2
port 844 nsew ground bidirectional
rlabel metal5 s -4816 455476 588740 456076 6 vssd2
port 845 nsew ground bidirectional
rlabel metal5 s -4816 419476 588740 420076 6 vssd2
port 846 nsew ground bidirectional
rlabel metal5 s -4816 383476 588740 384076 6 vssd2
port 847 nsew ground bidirectional
rlabel metal5 s -4816 347476 588740 348076 6 vssd2
port 848 nsew ground bidirectional
rlabel metal5 s -4816 311476 588740 312076 6 vssd2
port 849 nsew ground bidirectional
rlabel metal5 s -4816 275476 588740 276076 6 vssd2
port 850 nsew ground bidirectional
rlabel metal5 s -4816 239476 588740 240076 6 vssd2
port 851 nsew ground bidirectional
rlabel metal5 s -4816 203476 588740 204076 6 vssd2
port 852 nsew ground bidirectional
rlabel metal5 s -4816 167476 588740 168076 6 vssd2
port 853 nsew ground bidirectional
rlabel metal5 s -4816 131476 588740 132076 6 vssd2
port 854 nsew ground bidirectional
rlabel metal5 s -4816 95476 588740 96076 6 vssd2
port 855 nsew ground bidirectional
rlabel metal5 s -4816 59476 588740 60076 6 vssd2
port 856 nsew ground bidirectional
rlabel metal5 s -4816 23476 588740 24076 6 vssd2
port 857 nsew ground bidirectional
rlabel metal5 s -4816 -3744 588740 -3144 8 vssd2
port 858 nsew ground bidirectional
rlabel metal4 s 548004 698000 548604 709560 6 vdda1
port 859 nsew power bidirectional
rlabel metal4 s 512004 698000 512604 709560 6 vdda1
port 860 nsew power bidirectional
rlabel metal4 s 476004 698000 476604 709560 6 vdda1
port 861 nsew power bidirectional
rlabel metal4 s 440004 698000 440604 709560 6 vdda1
port 862 nsew power bidirectional
rlabel metal4 s 404004 698000 404604 709560 6 vdda1
port 863 nsew power bidirectional
rlabel metal4 s 368004 698000 368604 709560 6 vdda1
port 864 nsew power bidirectional
rlabel metal4 s 332004 698000 332604 709560 6 vdda1
port 865 nsew power bidirectional
rlabel metal4 s 296004 698000 296604 709560 6 vdda1
port 866 nsew power bidirectional
rlabel metal4 s 260004 698000 260604 709560 6 vdda1
port 867 nsew power bidirectional
rlabel metal4 s 224004 698000 224604 709560 6 vdda1
port 868 nsew power bidirectional
rlabel metal4 s 188004 698000 188604 709560 6 vdda1
port 869 nsew power bidirectional
rlabel metal4 s 152004 698000 152604 709560 6 vdda1
port 870 nsew power bidirectional
rlabel metal4 s 116004 698000 116604 709560 6 vdda1
port 871 nsew power bidirectional
rlabel metal4 s 80004 698000 80604 709560 6 vdda1
port 872 nsew power bidirectional
rlabel metal4 s 44004 698000 44604 709560 6 vdda1
port 873 nsew power bidirectional
rlabel metal4 s 8004 698000 8604 709560 6 vdda1
port 874 nsew power bidirectional
rlabel metal4 s 589080 -4684 589680 708620 6 vdda1
port 875 nsew power bidirectional
rlabel metal4 s -5756 -4684 -5156 708620 4 vdda1
port 876 nsew power bidirectional
rlabel metal4 s 548004 -5624 548604 6000 6 vdda1
port 877 nsew power bidirectional
rlabel metal4 s 512004 -5624 512604 6000 6 vdda1
port 878 nsew power bidirectional
rlabel metal4 s 476004 -5624 476604 6000 6 vdda1
port 879 nsew power bidirectional
rlabel metal4 s 440004 -5624 440604 6000 6 vdda1
port 880 nsew power bidirectional
rlabel metal4 s 404004 -5624 404604 6000 6 vdda1
port 881 nsew power bidirectional
rlabel metal4 s 368004 -5624 368604 6000 6 vdda1
port 882 nsew power bidirectional
rlabel metal4 s 332004 -5624 332604 6000 6 vdda1
port 883 nsew power bidirectional
rlabel metal4 s 296004 -5624 296604 6000 6 vdda1
port 884 nsew power bidirectional
rlabel metal4 s 260004 -5624 260604 6000 6 vdda1
port 885 nsew power bidirectional
rlabel metal4 s 224004 -5624 224604 6000 6 vdda1
port 886 nsew power bidirectional
rlabel metal4 s 188004 -5624 188604 6000 6 vdda1
port 887 nsew power bidirectional
rlabel metal4 s 152004 -5624 152604 6000 6 vdda1
port 888 nsew power bidirectional
rlabel metal4 s 116004 -5624 116604 6000 6 vdda1
port 889 nsew power bidirectional
rlabel metal4 s 80004 -5624 80604 6000 6 vdda1
port 890 nsew power bidirectional
rlabel metal4 s 44004 -5624 44604 6000 6 vdda1
port 891 nsew power bidirectional
rlabel metal4 s 8004 -5624 8604 6000 6 vdda1
port 892 nsew power bidirectional
rlabel metal5 s -5756 708020 589680 708620 6 vdda1
port 893 nsew power bidirectional
rlabel metal5 s -6696 693076 590620 693676 6 vdda1
port 894 nsew power bidirectional
rlabel metal5 s -6696 657076 590620 657676 6 vdda1
port 895 nsew power bidirectional
rlabel metal5 s -6696 621076 590620 621676 6 vdda1
port 896 nsew power bidirectional
rlabel metal5 s -6696 585076 590620 585676 6 vdda1
port 897 nsew power bidirectional
rlabel metal5 s -6696 549076 590620 549676 6 vdda1
port 898 nsew power bidirectional
rlabel metal5 s -6696 513076 590620 513676 6 vdda1
port 899 nsew power bidirectional
rlabel metal5 s -6696 477076 590620 477676 6 vdda1
port 900 nsew power bidirectional
rlabel metal5 s -6696 441076 590620 441676 6 vdda1
port 901 nsew power bidirectional
rlabel metal5 s -6696 405076 590620 405676 6 vdda1
port 902 nsew power bidirectional
rlabel metal5 s -6696 369076 590620 369676 6 vdda1
port 903 nsew power bidirectional
rlabel metal5 s -6696 333076 590620 333676 6 vdda1
port 904 nsew power bidirectional
rlabel metal5 s -6696 297076 590620 297676 6 vdda1
port 905 nsew power bidirectional
rlabel metal5 s -6696 261076 590620 261676 6 vdda1
port 906 nsew power bidirectional
rlabel metal5 s -6696 225076 590620 225676 6 vdda1
port 907 nsew power bidirectional
rlabel metal5 s -6696 189076 590620 189676 6 vdda1
port 908 nsew power bidirectional
rlabel metal5 s -6696 153076 590620 153676 6 vdda1
port 909 nsew power bidirectional
rlabel metal5 s -6696 117076 590620 117676 6 vdda1
port 910 nsew power bidirectional
rlabel metal5 s -6696 81076 590620 81676 6 vdda1
port 911 nsew power bidirectional
rlabel metal5 s -6696 45076 590620 45676 6 vdda1
port 912 nsew power bidirectional
rlabel metal5 s -6696 9076 590620 9676 6 vdda1
port 913 nsew power bidirectional
rlabel metal5 s -5756 -4684 589680 -4084 8 vdda1
port 914 nsew power bidirectional
rlabel metal4 s 590020 -5624 590620 709560 6 vssa1
port 915 nsew ground bidirectional
rlabel metal4 s 566004 698000 566604 709560 6 vssa1
port 916 nsew ground bidirectional
rlabel metal4 s 530004 698000 530604 709560 6 vssa1
port 917 nsew ground bidirectional
rlabel metal4 s 494004 698000 494604 709560 6 vssa1
port 918 nsew ground bidirectional
rlabel metal4 s 458004 698000 458604 709560 6 vssa1
port 919 nsew ground bidirectional
rlabel metal4 s 422004 698000 422604 709560 6 vssa1
port 920 nsew ground bidirectional
rlabel metal4 s 386004 698000 386604 709560 6 vssa1
port 921 nsew ground bidirectional
rlabel metal4 s 350004 698000 350604 709560 6 vssa1
port 922 nsew ground bidirectional
rlabel metal4 s 314004 698000 314604 709560 6 vssa1
port 923 nsew ground bidirectional
rlabel metal4 s 278004 698000 278604 709560 6 vssa1
port 924 nsew ground bidirectional
rlabel metal4 s 242004 698000 242604 709560 6 vssa1
port 925 nsew ground bidirectional
rlabel metal4 s 206004 698000 206604 709560 6 vssa1
port 926 nsew ground bidirectional
rlabel metal4 s 170004 698000 170604 709560 6 vssa1
port 927 nsew ground bidirectional
rlabel metal4 s 134004 698000 134604 709560 6 vssa1
port 928 nsew ground bidirectional
rlabel metal4 s 98004 698000 98604 709560 6 vssa1
port 929 nsew ground bidirectional
rlabel metal4 s 62004 698000 62604 709560 6 vssa1
port 930 nsew ground bidirectional
rlabel metal4 s 26004 698000 26604 709560 6 vssa1
port 931 nsew ground bidirectional
rlabel metal4 s -6696 -5624 -6096 709560 4 vssa1
port 932 nsew ground bidirectional
rlabel metal4 s 566004 -5624 566604 6000 6 vssa1
port 933 nsew ground bidirectional
rlabel metal4 s 530004 -5624 530604 6000 6 vssa1
port 934 nsew ground bidirectional
rlabel metal4 s 494004 -5624 494604 6000 6 vssa1
port 935 nsew ground bidirectional
rlabel metal4 s 458004 -5624 458604 6000 6 vssa1
port 936 nsew ground bidirectional
rlabel metal4 s 422004 -5624 422604 6000 6 vssa1
port 937 nsew ground bidirectional
rlabel metal4 s 386004 -5624 386604 6000 6 vssa1
port 938 nsew ground bidirectional
rlabel metal4 s 350004 -5624 350604 6000 6 vssa1
port 939 nsew ground bidirectional
rlabel metal4 s 314004 -5624 314604 6000 6 vssa1
port 940 nsew ground bidirectional
rlabel metal4 s 278004 -5624 278604 6000 6 vssa1
port 941 nsew ground bidirectional
rlabel metal4 s 242004 -5624 242604 6000 6 vssa1
port 942 nsew ground bidirectional
rlabel metal4 s 206004 -5624 206604 6000 6 vssa1
port 943 nsew ground bidirectional
rlabel metal4 s 170004 -5624 170604 6000 6 vssa1
port 944 nsew ground bidirectional
rlabel metal4 s 134004 -5624 134604 6000 6 vssa1
port 945 nsew ground bidirectional
rlabel metal4 s 98004 -5624 98604 6000 6 vssa1
port 946 nsew ground bidirectional
rlabel metal4 s 62004 -5624 62604 6000 6 vssa1
port 947 nsew ground bidirectional
rlabel metal4 s 26004 -5624 26604 6000 6 vssa1
port 948 nsew ground bidirectional
rlabel metal5 s -6696 708960 590620 709560 6 vssa1
port 949 nsew ground bidirectional
rlabel metal5 s -6696 675076 590620 675676 6 vssa1
port 950 nsew ground bidirectional
rlabel metal5 s -6696 639076 590620 639676 6 vssa1
port 951 nsew ground bidirectional
rlabel metal5 s -6696 603076 590620 603676 6 vssa1
port 952 nsew ground bidirectional
rlabel metal5 s -6696 567076 590620 567676 6 vssa1
port 953 nsew ground bidirectional
rlabel metal5 s -6696 531076 590620 531676 6 vssa1
port 954 nsew ground bidirectional
rlabel metal5 s -6696 495076 590620 495676 6 vssa1
port 955 nsew ground bidirectional
rlabel metal5 s -6696 459076 590620 459676 6 vssa1
port 956 nsew ground bidirectional
rlabel metal5 s -6696 423076 590620 423676 6 vssa1
port 957 nsew ground bidirectional
rlabel metal5 s -6696 387076 590620 387676 6 vssa1
port 958 nsew ground bidirectional
rlabel metal5 s -6696 351076 590620 351676 6 vssa1
port 959 nsew ground bidirectional
rlabel metal5 s -6696 315076 590620 315676 6 vssa1
port 960 nsew ground bidirectional
rlabel metal5 s -6696 279076 590620 279676 6 vssa1
port 961 nsew ground bidirectional
rlabel metal5 s -6696 243076 590620 243676 6 vssa1
port 962 nsew ground bidirectional
rlabel metal5 s -6696 207076 590620 207676 6 vssa1
port 963 nsew ground bidirectional
rlabel metal5 s -6696 171076 590620 171676 6 vssa1
port 964 nsew ground bidirectional
rlabel metal5 s -6696 135076 590620 135676 6 vssa1
port 965 nsew ground bidirectional
rlabel metal5 s -6696 99076 590620 99676 6 vssa1
port 966 nsew ground bidirectional
rlabel metal5 s -6696 63076 590620 63676 6 vssa1
port 967 nsew ground bidirectional
rlabel metal5 s -6696 27076 590620 27676 6 vssa1
port 968 nsew ground bidirectional
rlabel metal5 s -6696 -5624 590620 -5024 8 vssa1
port 969 nsew ground bidirectional
rlabel metal4 s 551604 698000 552204 711440 6 vdda2
port 970 nsew power bidirectional
rlabel metal4 s 515604 698000 516204 711440 6 vdda2
port 971 nsew power bidirectional
rlabel metal4 s 479604 698000 480204 711440 6 vdda2
port 972 nsew power bidirectional
rlabel metal4 s 443604 698000 444204 711440 6 vdda2
port 973 nsew power bidirectional
rlabel metal4 s 407604 698000 408204 711440 6 vdda2
port 974 nsew power bidirectional
rlabel metal4 s 371604 698000 372204 711440 6 vdda2
port 975 nsew power bidirectional
rlabel metal4 s 335604 698000 336204 711440 6 vdda2
port 976 nsew power bidirectional
rlabel metal4 s 299604 698000 300204 711440 6 vdda2
port 977 nsew power bidirectional
rlabel metal4 s 263604 698000 264204 711440 6 vdda2
port 978 nsew power bidirectional
rlabel metal4 s 227604 698000 228204 711440 6 vdda2
port 979 nsew power bidirectional
rlabel metal4 s 191604 698000 192204 711440 6 vdda2
port 980 nsew power bidirectional
rlabel metal4 s 155604 698000 156204 711440 6 vdda2
port 981 nsew power bidirectional
rlabel metal4 s 119604 698000 120204 711440 6 vdda2
port 982 nsew power bidirectional
rlabel metal4 s 83604 698000 84204 711440 6 vdda2
port 983 nsew power bidirectional
rlabel metal4 s 47604 698000 48204 711440 6 vdda2
port 984 nsew power bidirectional
rlabel metal4 s 11604 698000 12204 711440 6 vdda2
port 985 nsew power bidirectional
rlabel metal4 s 590960 -6564 591560 710500 6 vdda2
port 986 nsew power bidirectional
rlabel metal4 s -7636 -6564 -7036 710500 4 vdda2
port 987 nsew power bidirectional
rlabel metal4 s 551604 -7504 552204 6000 8 vdda2
port 988 nsew power bidirectional
rlabel metal4 s 515604 -7504 516204 6000 8 vdda2
port 989 nsew power bidirectional
rlabel metal4 s 479604 -7504 480204 6000 8 vdda2
port 990 nsew power bidirectional
rlabel metal4 s 443604 -7504 444204 6000 8 vdda2
port 991 nsew power bidirectional
rlabel metal4 s 407604 -7504 408204 6000 8 vdda2
port 992 nsew power bidirectional
rlabel metal4 s 371604 -7504 372204 6000 8 vdda2
port 993 nsew power bidirectional
rlabel metal4 s 335604 -7504 336204 6000 8 vdda2
port 994 nsew power bidirectional
rlabel metal4 s 299604 -7504 300204 6000 8 vdda2
port 995 nsew power bidirectional
rlabel metal4 s 263604 -7504 264204 6000 8 vdda2
port 996 nsew power bidirectional
rlabel metal4 s 227604 -7504 228204 6000 8 vdda2
port 997 nsew power bidirectional
rlabel metal4 s 191604 -7504 192204 6000 8 vdda2
port 998 nsew power bidirectional
rlabel metal4 s 155604 -7504 156204 6000 8 vdda2
port 999 nsew power bidirectional
rlabel metal4 s 119604 -7504 120204 6000 8 vdda2
port 1000 nsew power bidirectional
rlabel metal4 s 83604 -7504 84204 6000 8 vdda2
port 1001 nsew power bidirectional
rlabel metal4 s 47604 -7504 48204 6000 8 vdda2
port 1002 nsew power bidirectional
rlabel metal4 s 11604 -7504 12204 6000 8 vdda2
port 1003 nsew power bidirectional
rlabel metal5 s -7636 709900 591560 710500 6 vdda2
port 1004 nsew power bidirectional
rlabel metal5 s -8576 696676 592500 697276 6 vdda2
port 1005 nsew power bidirectional
rlabel metal5 s -8576 660676 592500 661276 6 vdda2
port 1006 nsew power bidirectional
rlabel metal5 s -8576 624676 592500 625276 6 vdda2
port 1007 nsew power bidirectional
rlabel metal5 s -8576 588676 592500 589276 6 vdda2
port 1008 nsew power bidirectional
rlabel metal5 s -8576 552676 592500 553276 6 vdda2
port 1009 nsew power bidirectional
rlabel metal5 s -8576 516676 592500 517276 6 vdda2
port 1010 nsew power bidirectional
rlabel metal5 s -8576 480676 592500 481276 6 vdda2
port 1011 nsew power bidirectional
rlabel metal5 s -8576 444676 592500 445276 6 vdda2
port 1012 nsew power bidirectional
rlabel metal5 s -8576 408676 592500 409276 6 vdda2
port 1013 nsew power bidirectional
rlabel metal5 s -8576 372676 592500 373276 6 vdda2
port 1014 nsew power bidirectional
rlabel metal5 s -8576 336676 592500 337276 6 vdda2
port 1015 nsew power bidirectional
rlabel metal5 s -8576 300676 592500 301276 6 vdda2
port 1016 nsew power bidirectional
rlabel metal5 s -8576 264676 592500 265276 6 vdda2
port 1017 nsew power bidirectional
rlabel metal5 s -8576 228676 592500 229276 6 vdda2
port 1018 nsew power bidirectional
rlabel metal5 s -8576 192676 592500 193276 6 vdda2
port 1019 nsew power bidirectional
rlabel metal5 s -8576 156676 592500 157276 6 vdda2
port 1020 nsew power bidirectional
rlabel metal5 s -8576 120676 592500 121276 6 vdda2
port 1021 nsew power bidirectional
rlabel metal5 s -8576 84676 592500 85276 6 vdda2
port 1022 nsew power bidirectional
rlabel metal5 s -8576 48676 592500 49276 6 vdda2
port 1023 nsew power bidirectional
rlabel metal5 s -8576 12676 592500 13276 6 vdda2
port 1024 nsew power bidirectional
rlabel metal5 s -7636 -6564 591560 -5964 8 vdda2
port 1025 nsew power bidirectional
rlabel metal4 s 591900 -7504 592500 711440 6 vssa2
port 1026 nsew ground bidirectional
rlabel metal4 s 569604 698000 570204 711440 6 vssa2
port 1027 nsew ground bidirectional
rlabel metal4 s 533604 698000 534204 711440 6 vssa2
port 1028 nsew ground bidirectional
rlabel metal4 s 497604 698000 498204 711440 6 vssa2
port 1029 nsew ground bidirectional
rlabel metal4 s 461604 698000 462204 711440 6 vssa2
port 1030 nsew ground bidirectional
rlabel metal4 s 425604 698000 426204 711440 6 vssa2
port 1031 nsew ground bidirectional
rlabel metal4 s 389604 698000 390204 711440 6 vssa2
port 1032 nsew ground bidirectional
rlabel metal4 s 353604 698000 354204 711440 6 vssa2
port 1033 nsew ground bidirectional
rlabel metal4 s 317604 698000 318204 711440 6 vssa2
port 1034 nsew ground bidirectional
rlabel metal4 s 281604 698000 282204 711440 6 vssa2
port 1035 nsew ground bidirectional
rlabel metal4 s 245604 698000 246204 711440 6 vssa2
port 1036 nsew ground bidirectional
rlabel metal4 s 209604 698000 210204 711440 6 vssa2
port 1037 nsew ground bidirectional
rlabel metal4 s 173604 698000 174204 711440 6 vssa2
port 1038 nsew ground bidirectional
rlabel metal4 s 137604 698000 138204 711440 6 vssa2
port 1039 nsew ground bidirectional
rlabel metal4 s 101604 698000 102204 711440 6 vssa2
port 1040 nsew ground bidirectional
rlabel metal4 s 65604 698000 66204 711440 6 vssa2
port 1041 nsew ground bidirectional
rlabel metal4 s 29604 698000 30204 711440 6 vssa2
port 1042 nsew ground bidirectional
rlabel metal4 s -8576 -7504 -7976 711440 4 vssa2
port 1043 nsew ground bidirectional
rlabel metal4 s 569604 -7504 570204 6000 8 vssa2
port 1044 nsew ground bidirectional
rlabel metal4 s 533604 -7504 534204 6000 8 vssa2
port 1045 nsew ground bidirectional
rlabel metal4 s 497604 -7504 498204 6000 8 vssa2
port 1046 nsew ground bidirectional
rlabel metal4 s 461604 -7504 462204 6000 8 vssa2
port 1047 nsew ground bidirectional
rlabel metal4 s 425604 -7504 426204 6000 8 vssa2
port 1048 nsew ground bidirectional
rlabel metal4 s 389604 -7504 390204 6000 8 vssa2
port 1049 nsew ground bidirectional
rlabel metal4 s 353604 -7504 354204 6000 8 vssa2
port 1050 nsew ground bidirectional
rlabel metal4 s 317604 -7504 318204 6000 8 vssa2
port 1051 nsew ground bidirectional
rlabel metal4 s 281604 -7504 282204 6000 8 vssa2
port 1052 nsew ground bidirectional
rlabel metal4 s 245604 -7504 246204 6000 8 vssa2
port 1053 nsew ground bidirectional
rlabel metal4 s 209604 -7504 210204 6000 8 vssa2
port 1054 nsew ground bidirectional
rlabel metal4 s 173604 -7504 174204 6000 8 vssa2
port 1055 nsew ground bidirectional
rlabel metal4 s 137604 -7504 138204 6000 8 vssa2
port 1056 nsew ground bidirectional
rlabel metal4 s 101604 -7504 102204 6000 8 vssa2
port 1057 nsew ground bidirectional
rlabel metal4 s 65604 -7504 66204 6000 8 vssa2
port 1058 nsew ground bidirectional
rlabel metal4 s 29604 -7504 30204 6000 8 vssa2
port 1059 nsew ground bidirectional
rlabel metal5 s -8576 710840 592500 711440 6 vssa2
port 1060 nsew ground bidirectional
rlabel metal5 s -8576 678676 592500 679276 6 vssa2
port 1061 nsew ground bidirectional
rlabel metal5 s -8576 642676 592500 643276 6 vssa2
port 1062 nsew ground bidirectional
rlabel metal5 s -8576 606676 592500 607276 6 vssa2
port 1063 nsew ground bidirectional
rlabel metal5 s -8576 570676 592500 571276 6 vssa2
port 1064 nsew ground bidirectional
rlabel metal5 s -8576 534676 592500 535276 6 vssa2
port 1065 nsew ground bidirectional
rlabel metal5 s -8576 498676 592500 499276 6 vssa2
port 1066 nsew ground bidirectional
rlabel metal5 s -8576 462676 592500 463276 6 vssa2
port 1067 nsew ground bidirectional
rlabel metal5 s -8576 426676 592500 427276 6 vssa2
port 1068 nsew ground bidirectional
rlabel metal5 s -8576 390676 592500 391276 6 vssa2
port 1069 nsew ground bidirectional
rlabel metal5 s -8576 354676 592500 355276 6 vssa2
port 1070 nsew ground bidirectional
rlabel metal5 s -8576 318676 592500 319276 6 vssa2
port 1071 nsew ground bidirectional
rlabel metal5 s -8576 282676 592500 283276 6 vssa2
port 1072 nsew ground bidirectional
rlabel metal5 s -8576 246676 592500 247276 6 vssa2
port 1073 nsew ground bidirectional
rlabel metal5 s -8576 210676 592500 211276 6 vssa2
port 1074 nsew ground bidirectional
rlabel metal5 s -8576 174676 592500 175276 6 vssa2
port 1075 nsew ground bidirectional
rlabel metal5 s -8576 138676 592500 139276 6 vssa2
port 1076 nsew ground bidirectional
rlabel metal5 s -8576 102676 592500 103276 6 vssa2
port 1077 nsew ground bidirectional
rlabel metal5 s -8576 66676 592500 67276 6 vssa2
port 1078 nsew ground bidirectional
rlabel metal5 s -8576 30676 592500 31276 6 vssa2
port 1079 nsew ground bidirectional
rlabel metal5 s -8576 -7504 592500 -6904 8 vssa2
port 1080 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>

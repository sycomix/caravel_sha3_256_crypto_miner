magic
tech sky130A
magscale 1 2
timestamp 1608503375
<< obsli1 >>
rect 1104 2159 566812 685457
<< obsm1 >>
rect 14 1096 566812 685488
<< metal2 >>
rect 2318 687200 2374 688000
rect 6918 687200 6974 688000
rect 11518 687200 11574 688000
rect 16118 687200 16174 688000
rect 20718 687200 20774 688000
rect 25318 687200 25374 688000
rect 30010 687200 30066 688000
rect 34610 687200 34666 688000
rect 39210 687200 39266 688000
rect 43810 687200 43866 688000
rect 48410 687200 48466 688000
rect 53102 687200 53158 688000
rect 57702 687200 57758 688000
rect 62302 687200 62358 688000
rect 66902 687200 66958 688000
rect 71502 687200 71558 688000
rect 76194 687200 76250 688000
rect 80794 687200 80850 688000
rect 85394 687200 85450 688000
rect 89994 687200 90050 688000
rect 94594 687200 94650 688000
rect 99286 687200 99342 688000
rect 103886 687200 103942 688000
rect 108486 687200 108542 688000
rect 113086 687200 113142 688000
rect 117686 687200 117742 688000
rect 122378 687200 122434 688000
rect 126978 687200 127034 688000
rect 131578 687200 131634 688000
rect 136178 687200 136234 688000
rect 140778 687200 140834 688000
rect 145470 687200 145526 688000
rect 150070 687200 150126 688000
rect 154670 687200 154726 688000
rect 159270 687200 159326 688000
rect 163870 687200 163926 688000
rect 168562 687200 168618 688000
rect 173162 687200 173218 688000
rect 177762 687200 177818 688000
rect 182362 687200 182418 688000
rect 186962 687200 187018 688000
rect 191654 687200 191710 688000
rect 196254 687200 196310 688000
rect 200854 687200 200910 688000
rect 205454 687200 205510 688000
rect 210054 687200 210110 688000
rect 214654 687200 214710 688000
rect 219346 687200 219402 688000
rect 223946 687200 224002 688000
rect 228546 687200 228602 688000
rect 233146 687200 233202 688000
rect 237746 687200 237802 688000
rect 242438 687200 242494 688000
rect 247038 687200 247094 688000
rect 251638 687200 251694 688000
rect 256238 687200 256294 688000
rect 260838 687200 260894 688000
rect 265530 687200 265586 688000
rect 270130 687200 270186 688000
rect 274730 687200 274786 688000
rect 279330 687200 279386 688000
rect 283930 687200 283986 688000
rect 288622 687200 288678 688000
rect 293222 687200 293278 688000
rect 297822 687200 297878 688000
rect 302422 687200 302478 688000
rect 307022 687200 307078 688000
rect 311714 687200 311770 688000
rect 316314 687200 316370 688000
rect 320914 687200 320970 688000
rect 325514 687200 325570 688000
rect 330114 687200 330170 688000
rect 334806 687200 334862 688000
rect 339406 687200 339462 688000
rect 344006 687200 344062 688000
rect 348606 687200 348662 688000
rect 353206 687200 353262 688000
rect 357898 687200 357954 688000
rect 362498 687200 362554 688000
rect 367098 687200 367154 688000
rect 371698 687200 371754 688000
rect 376298 687200 376354 688000
rect 380990 687200 381046 688000
rect 385590 687200 385646 688000
rect 390190 687200 390246 688000
rect 394790 687200 394846 688000
rect 399390 687200 399446 688000
rect 403990 687200 404046 688000
rect 408682 687200 408738 688000
rect 413282 687200 413338 688000
rect 417882 687200 417938 688000
rect 422482 687200 422538 688000
rect 427082 687200 427138 688000
rect 431774 687200 431830 688000
rect 436374 687200 436430 688000
rect 440974 687200 441030 688000
rect 445574 687200 445630 688000
rect 450174 687200 450230 688000
rect 454866 687200 454922 688000
rect 459466 687200 459522 688000
rect 464066 687200 464122 688000
rect 468666 687200 468722 688000
rect 473266 687200 473322 688000
rect 477958 687200 478014 688000
rect 482558 687200 482614 688000
rect 487158 687200 487214 688000
rect 491758 687200 491814 688000
rect 496358 687200 496414 688000
rect 501050 687200 501106 688000
rect 505650 687200 505706 688000
rect 510250 687200 510306 688000
rect 514850 687200 514906 688000
rect 519450 687200 519506 688000
rect 524142 687200 524198 688000
rect 528742 687200 528798 688000
rect 533342 687200 533398 688000
rect 537942 687200 537998 688000
rect 542542 687200 542598 688000
rect 547234 687200 547290 688000
rect 551834 687200 551890 688000
rect 556434 687200 556490 688000
rect 561034 687200 561090 688000
rect 565634 687200 565690 688000
rect 570 0 626 800
rect 1674 0 1730 800
rect 2778 0 2834 800
rect 3974 0 4030 800
rect 5078 0 5134 800
rect 6182 0 6238 800
rect 7378 0 7434 800
rect 8482 0 8538 800
rect 9586 0 9642 800
rect 10782 0 10838 800
rect 11886 0 11942 800
rect 12990 0 13046 800
rect 14186 0 14242 800
rect 15290 0 15346 800
rect 16394 0 16450 800
rect 17590 0 17646 800
rect 18694 0 18750 800
rect 19798 0 19854 800
rect 20994 0 21050 800
rect 22098 0 22154 800
rect 23202 0 23258 800
rect 24398 0 24454 800
rect 25502 0 25558 800
rect 26698 0 26754 800
rect 27802 0 27858 800
rect 28906 0 28962 800
rect 30102 0 30158 800
rect 31206 0 31262 800
rect 32310 0 32366 800
rect 33506 0 33562 800
rect 34610 0 34666 800
rect 35714 0 35770 800
rect 36910 0 36966 800
rect 38014 0 38070 800
rect 39118 0 39174 800
rect 40314 0 40370 800
rect 41418 0 41474 800
rect 42522 0 42578 800
rect 43718 0 43774 800
rect 44822 0 44878 800
rect 45926 0 45982 800
rect 47122 0 47178 800
rect 48226 0 48282 800
rect 49330 0 49386 800
rect 50526 0 50582 800
rect 51630 0 51686 800
rect 52826 0 52882 800
rect 53930 0 53986 800
rect 55034 0 55090 800
rect 56230 0 56286 800
rect 57334 0 57390 800
rect 58438 0 58494 800
rect 59634 0 59690 800
rect 60738 0 60794 800
rect 61842 0 61898 800
rect 63038 0 63094 800
rect 64142 0 64198 800
rect 65246 0 65302 800
rect 66442 0 66498 800
rect 67546 0 67602 800
rect 68650 0 68706 800
rect 69846 0 69902 800
rect 70950 0 71006 800
rect 72054 0 72110 800
rect 73250 0 73306 800
rect 74354 0 74410 800
rect 75458 0 75514 800
rect 76654 0 76710 800
rect 77758 0 77814 800
rect 78954 0 79010 800
rect 80058 0 80114 800
rect 81162 0 81218 800
rect 82358 0 82414 800
rect 83462 0 83518 800
rect 84566 0 84622 800
rect 85762 0 85818 800
rect 86866 0 86922 800
rect 87970 0 88026 800
rect 89166 0 89222 800
rect 90270 0 90326 800
rect 91374 0 91430 800
rect 92570 0 92626 800
rect 93674 0 93730 800
rect 94778 0 94834 800
rect 95974 0 96030 800
rect 97078 0 97134 800
rect 98182 0 98238 800
rect 99378 0 99434 800
rect 100482 0 100538 800
rect 101586 0 101642 800
rect 102782 0 102838 800
rect 103886 0 103942 800
rect 105082 0 105138 800
rect 106186 0 106242 800
rect 107290 0 107346 800
rect 108486 0 108542 800
rect 109590 0 109646 800
rect 110694 0 110750 800
rect 111890 0 111946 800
rect 112994 0 113050 800
rect 114098 0 114154 800
rect 115294 0 115350 800
rect 116398 0 116454 800
rect 117502 0 117558 800
rect 118698 0 118754 800
rect 119802 0 119858 800
rect 120906 0 120962 800
rect 122102 0 122158 800
rect 123206 0 123262 800
rect 124310 0 124366 800
rect 125506 0 125562 800
rect 126610 0 126666 800
rect 127714 0 127770 800
rect 128910 0 128966 800
rect 130014 0 130070 800
rect 131210 0 131266 800
rect 132314 0 132370 800
rect 133418 0 133474 800
rect 134614 0 134670 800
rect 135718 0 135774 800
rect 136822 0 136878 800
rect 138018 0 138074 800
rect 139122 0 139178 800
rect 140226 0 140282 800
rect 141422 0 141478 800
rect 142526 0 142582 800
rect 143630 0 143686 800
rect 144826 0 144882 800
rect 145930 0 145986 800
rect 147034 0 147090 800
rect 148230 0 148286 800
rect 149334 0 149390 800
rect 150438 0 150494 800
rect 151634 0 151690 800
rect 152738 0 152794 800
rect 153842 0 153898 800
rect 155038 0 155094 800
rect 156142 0 156198 800
rect 157338 0 157394 800
rect 158442 0 158498 800
rect 159546 0 159602 800
rect 160742 0 160798 800
rect 161846 0 161902 800
rect 162950 0 163006 800
rect 164146 0 164202 800
rect 165250 0 165306 800
rect 166354 0 166410 800
rect 167550 0 167606 800
rect 168654 0 168710 800
rect 169758 0 169814 800
rect 170954 0 171010 800
rect 172058 0 172114 800
rect 173162 0 173218 800
rect 174358 0 174414 800
rect 175462 0 175518 800
rect 176566 0 176622 800
rect 177762 0 177818 800
rect 178866 0 178922 800
rect 179970 0 180026 800
rect 181166 0 181222 800
rect 182270 0 182326 800
rect 183466 0 183522 800
rect 184570 0 184626 800
rect 185674 0 185730 800
rect 186870 0 186926 800
rect 187974 0 188030 800
rect 189078 0 189134 800
rect 190274 0 190330 800
rect 191378 0 191434 800
rect 192482 0 192538 800
rect 193678 0 193734 800
rect 194782 0 194838 800
rect 195886 0 195942 800
rect 197082 0 197138 800
rect 198186 0 198242 800
rect 199290 0 199346 800
rect 200486 0 200542 800
rect 201590 0 201646 800
rect 202694 0 202750 800
rect 203890 0 203946 800
rect 204994 0 205050 800
rect 206098 0 206154 800
rect 207294 0 207350 800
rect 208398 0 208454 800
rect 209594 0 209650 800
rect 210698 0 210754 800
rect 211802 0 211858 800
rect 212998 0 213054 800
rect 214102 0 214158 800
rect 215206 0 215262 800
rect 216402 0 216458 800
rect 217506 0 217562 800
rect 218610 0 218666 800
rect 219806 0 219862 800
rect 220910 0 220966 800
rect 222014 0 222070 800
rect 223210 0 223266 800
rect 224314 0 224370 800
rect 225418 0 225474 800
rect 226614 0 226670 800
rect 227718 0 227774 800
rect 228822 0 228878 800
rect 230018 0 230074 800
rect 231122 0 231178 800
rect 232226 0 232282 800
rect 233422 0 233478 800
rect 234526 0 234582 800
rect 235722 0 235778 800
rect 236826 0 236882 800
rect 237930 0 237986 800
rect 239126 0 239182 800
rect 240230 0 240286 800
rect 241334 0 241390 800
rect 242530 0 242586 800
rect 243634 0 243690 800
rect 244738 0 244794 800
rect 245934 0 245990 800
rect 247038 0 247094 800
rect 248142 0 248198 800
rect 249338 0 249394 800
rect 250442 0 250498 800
rect 251546 0 251602 800
rect 252742 0 252798 800
rect 253846 0 253902 800
rect 254950 0 255006 800
rect 256146 0 256202 800
rect 257250 0 257306 800
rect 258354 0 258410 800
rect 259550 0 259606 800
rect 260654 0 260710 800
rect 261850 0 261906 800
rect 262954 0 263010 800
rect 264058 0 264114 800
rect 265254 0 265310 800
rect 266358 0 266414 800
rect 267462 0 267518 800
rect 268658 0 268714 800
rect 269762 0 269818 800
rect 270866 0 270922 800
rect 272062 0 272118 800
rect 273166 0 273222 800
rect 274270 0 274326 800
rect 275466 0 275522 800
rect 276570 0 276626 800
rect 277674 0 277730 800
rect 278870 0 278926 800
rect 279974 0 280030 800
rect 281078 0 281134 800
rect 282274 0 282330 800
rect 283378 0 283434 800
rect 284574 0 284630 800
rect 285678 0 285734 800
rect 286782 0 286838 800
rect 287978 0 288034 800
rect 289082 0 289138 800
rect 290186 0 290242 800
rect 291382 0 291438 800
rect 292486 0 292542 800
rect 293590 0 293646 800
rect 294786 0 294842 800
rect 295890 0 295946 800
rect 296994 0 297050 800
rect 298190 0 298246 800
rect 299294 0 299350 800
rect 300398 0 300454 800
rect 301594 0 301650 800
rect 302698 0 302754 800
rect 303802 0 303858 800
rect 304998 0 305054 800
rect 306102 0 306158 800
rect 307206 0 307262 800
rect 308402 0 308458 800
rect 309506 0 309562 800
rect 310702 0 310758 800
rect 311806 0 311862 800
rect 312910 0 312966 800
rect 314106 0 314162 800
rect 315210 0 315266 800
rect 316314 0 316370 800
rect 317510 0 317566 800
rect 318614 0 318670 800
rect 319718 0 319774 800
rect 320914 0 320970 800
rect 322018 0 322074 800
rect 323122 0 323178 800
rect 324318 0 324374 800
rect 325422 0 325478 800
rect 326526 0 326582 800
rect 327722 0 327778 800
rect 328826 0 328882 800
rect 329930 0 329986 800
rect 331126 0 331182 800
rect 332230 0 332286 800
rect 333334 0 333390 800
rect 334530 0 334586 800
rect 335634 0 335690 800
rect 336830 0 336886 800
rect 337934 0 337990 800
rect 339038 0 339094 800
rect 340234 0 340290 800
rect 341338 0 341394 800
rect 342442 0 342498 800
rect 343638 0 343694 800
rect 344742 0 344798 800
rect 345846 0 345902 800
rect 347042 0 347098 800
rect 348146 0 348202 800
rect 349250 0 349306 800
rect 350446 0 350502 800
rect 351550 0 351606 800
rect 352654 0 352710 800
rect 353850 0 353906 800
rect 354954 0 355010 800
rect 356058 0 356114 800
rect 357254 0 357310 800
rect 358358 0 358414 800
rect 359462 0 359518 800
rect 360658 0 360714 800
rect 361762 0 361818 800
rect 362958 0 363014 800
rect 364062 0 364118 800
rect 365166 0 365222 800
rect 366362 0 366418 800
rect 367466 0 367522 800
rect 368570 0 368626 800
rect 369766 0 369822 800
rect 370870 0 370926 800
rect 371974 0 372030 800
rect 373170 0 373226 800
rect 374274 0 374330 800
rect 375378 0 375434 800
rect 376574 0 376630 800
rect 377678 0 377734 800
rect 378782 0 378838 800
rect 379978 0 380034 800
rect 381082 0 381138 800
rect 382186 0 382242 800
rect 383382 0 383438 800
rect 384486 0 384542 800
rect 385590 0 385646 800
rect 386786 0 386842 800
rect 387890 0 387946 800
rect 389086 0 389142 800
rect 390190 0 390246 800
rect 391294 0 391350 800
rect 392490 0 392546 800
rect 393594 0 393650 800
rect 394698 0 394754 800
rect 395894 0 395950 800
rect 396998 0 397054 800
rect 398102 0 398158 800
rect 399298 0 399354 800
rect 400402 0 400458 800
rect 401506 0 401562 800
rect 402702 0 402758 800
rect 403806 0 403862 800
rect 404910 0 404966 800
rect 406106 0 406162 800
rect 407210 0 407266 800
rect 408314 0 408370 800
rect 409510 0 409566 800
rect 410614 0 410670 800
rect 411718 0 411774 800
rect 412914 0 412970 800
rect 414018 0 414074 800
rect 415214 0 415270 800
rect 416318 0 416374 800
rect 417422 0 417478 800
rect 418618 0 418674 800
rect 419722 0 419778 800
rect 420826 0 420882 800
rect 422022 0 422078 800
rect 423126 0 423182 800
rect 424230 0 424286 800
rect 425426 0 425482 800
rect 426530 0 426586 800
rect 427634 0 427690 800
rect 428830 0 428886 800
rect 429934 0 429990 800
rect 431038 0 431094 800
rect 432234 0 432290 800
rect 433338 0 433394 800
rect 434442 0 434498 800
rect 435638 0 435694 800
rect 436742 0 436798 800
rect 437846 0 437902 800
rect 439042 0 439098 800
rect 440146 0 440202 800
rect 441342 0 441398 800
rect 442446 0 442502 800
rect 443550 0 443606 800
rect 444746 0 444802 800
rect 445850 0 445906 800
rect 446954 0 447010 800
rect 448150 0 448206 800
rect 449254 0 449310 800
rect 450358 0 450414 800
rect 451554 0 451610 800
rect 452658 0 452714 800
rect 453762 0 453818 800
rect 454958 0 455014 800
rect 456062 0 456118 800
rect 457166 0 457222 800
rect 458362 0 458418 800
rect 459466 0 459522 800
rect 460570 0 460626 800
rect 461766 0 461822 800
rect 462870 0 462926 800
rect 463974 0 464030 800
rect 465170 0 465226 800
rect 466274 0 466330 800
rect 467470 0 467526 800
rect 468574 0 468630 800
rect 469678 0 469734 800
rect 470874 0 470930 800
rect 471978 0 472034 800
rect 473082 0 473138 800
rect 474278 0 474334 800
rect 475382 0 475438 800
rect 476486 0 476542 800
rect 477682 0 477738 800
rect 478786 0 478842 800
rect 479890 0 479946 800
rect 481086 0 481142 800
rect 482190 0 482246 800
rect 483294 0 483350 800
rect 484490 0 484546 800
rect 485594 0 485650 800
rect 486698 0 486754 800
rect 487894 0 487950 800
rect 488998 0 489054 800
rect 490102 0 490158 800
rect 491298 0 491354 800
rect 492402 0 492458 800
rect 493598 0 493654 800
rect 494702 0 494758 800
rect 495806 0 495862 800
rect 497002 0 497058 800
rect 498106 0 498162 800
rect 499210 0 499266 800
rect 500406 0 500462 800
rect 501510 0 501566 800
rect 502614 0 502670 800
rect 503810 0 503866 800
rect 504914 0 504970 800
rect 506018 0 506074 800
rect 507214 0 507270 800
rect 508318 0 508374 800
rect 509422 0 509478 800
rect 510618 0 510674 800
rect 511722 0 511778 800
rect 512826 0 512882 800
rect 514022 0 514078 800
rect 515126 0 515182 800
rect 516230 0 516286 800
rect 517426 0 517482 800
rect 518530 0 518586 800
rect 519726 0 519782 800
rect 520830 0 520886 800
rect 521934 0 521990 800
rect 523130 0 523186 800
rect 524234 0 524290 800
rect 525338 0 525394 800
rect 526534 0 526590 800
rect 527638 0 527694 800
rect 528742 0 528798 800
rect 529938 0 529994 800
rect 531042 0 531098 800
rect 532146 0 532202 800
rect 533342 0 533398 800
rect 534446 0 534502 800
rect 535550 0 535606 800
rect 536746 0 536802 800
rect 537850 0 537906 800
rect 538954 0 539010 800
rect 540150 0 540206 800
rect 541254 0 541310 800
rect 542358 0 542414 800
rect 543554 0 543610 800
rect 544658 0 544714 800
rect 545854 0 545910 800
rect 546958 0 547014 800
rect 548062 0 548118 800
rect 549258 0 549314 800
rect 550362 0 550418 800
rect 551466 0 551522 800
rect 552662 0 552718 800
rect 553766 0 553822 800
rect 554870 0 554926 800
rect 556066 0 556122 800
rect 557170 0 557226 800
rect 558274 0 558330 800
rect 559470 0 559526 800
rect 560574 0 560630 800
rect 561678 0 561734 800
rect 562874 0 562930 800
rect 563978 0 564034 800
rect 565082 0 565138 800
rect 566278 0 566334 800
rect 567382 0 567438 800
<< obsm2 >>
rect 20 687144 2262 687200
rect 2430 687144 6862 687200
rect 7030 687144 11462 687200
rect 11630 687144 16062 687200
rect 16230 687144 20662 687200
rect 20830 687144 25262 687200
rect 25430 687144 29954 687200
rect 30122 687144 34554 687200
rect 34722 687144 39154 687200
rect 39322 687144 43754 687200
rect 43922 687144 48354 687200
rect 48522 687144 53046 687200
rect 53214 687144 57646 687200
rect 57814 687144 62246 687200
rect 62414 687144 66846 687200
rect 67014 687144 71446 687200
rect 71614 687144 76138 687200
rect 76306 687144 80738 687200
rect 80906 687144 85338 687200
rect 85506 687144 89938 687200
rect 90106 687144 94538 687200
rect 94706 687144 99230 687200
rect 99398 687144 103830 687200
rect 103998 687144 108430 687200
rect 108598 687144 113030 687200
rect 113198 687144 117630 687200
rect 117798 687144 122322 687200
rect 122490 687144 126922 687200
rect 127090 687144 131522 687200
rect 131690 687144 136122 687200
rect 136290 687144 140722 687200
rect 140890 687144 145414 687200
rect 145582 687144 150014 687200
rect 150182 687144 154614 687200
rect 154782 687144 159214 687200
rect 159382 687144 163814 687200
rect 163982 687144 168506 687200
rect 168674 687144 173106 687200
rect 173274 687144 177706 687200
rect 177874 687144 182306 687200
rect 182474 687144 186906 687200
rect 187074 687144 191598 687200
rect 191766 687144 196198 687200
rect 196366 687144 200798 687200
rect 200966 687144 205398 687200
rect 205566 687144 209998 687200
rect 210166 687144 214598 687200
rect 214766 687144 219290 687200
rect 219458 687144 223890 687200
rect 224058 687144 228490 687200
rect 228658 687144 233090 687200
rect 233258 687144 237690 687200
rect 237858 687144 242382 687200
rect 242550 687144 246982 687200
rect 247150 687144 251582 687200
rect 251750 687144 256182 687200
rect 256350 687144 260782 687200
rect 260950 687144 265474 687200
rect 265642 687144 270074 687200
rect 270242 687144 274674 687200
rect 274842 687144 279274 687200
rect 279442 687144 283874 687200
rect 284042 687144 288566 687200
rect 288734 687144 293166 687200
rect 293334 687144 297766 687200
rect 297934 687144 302366 687200
rect 302534 687144 306966 687200
rect 307134 687144 311658 687200
rect 311826 687144 316258 687200
rect 316426 687144 320858 687200
rect 321026 687144 325458 687200
rect 325626 687144 330058 687200
rect 330226 687144 334750 687200
rect 334918 687144 339350 687200
rect 339518 687144 343950 687200
rect 344118 687144 348550 687200
rect 348718 687144 353150 687200
rect 353318 687144 357842 687200
rect 358010 687144 362442 687200
rect 362610 687144 367042 687200
rect 367210 687144 371642 687200
rect 371810 687144 376242 687200
rect 376410 687144 380934 687200
rect 381102 687144 385534 687200
rect 385702 687144 390134 687200
rect 390302 687144 394734 687200
rect 394902 687144 399334 687200
rect 399502 687144 403934 687200
rect 404102 687144 408626 687200
rect 408794 687144 413226 687200
rect 413394 687144 417826 687200
rect 417994 687144 422426 687200
rect 422594 687144 427026 687200
rect 427194 687144 431718 687200
rect 431886 687144 436318 687200
rect 436486 687144 440918 687200
rect 441086 687144 445518 687200
rect 445686 687144 450118 687200
rect 450286 687144 454810 687200
rect 454978 687144 459410 687200
rect 459578 687144 464010 687200
rect 464178 687144 468610 687200
rect 468778 687144 473210 687200
rect 473378 687144 477902 687200
rect 478070 687144 482502 687200
rect 482670 687144 487102 687200
rect 487270 687144 491702 687200
rect 491870 687144 496302 687200
rect 496470 687144 500994 687200
rect 501162 687144 505594 687200
rect 505762 687144 510194 687200
rect 510362 687144 514794 687200
rect 514962 687144 519394 687200
rect 519562 687144 524086 687200
rect 524254 687144 528686 687200
rect 528854 687144 533286 687200
rect 533454 687144 537886 687200
rect 538054 687144 542486 687200
rect 542654 687144 547178 687200
rect 547346 687144 551778 687200
rect 551946 687144 556378 687200
rect 556546 687144 557476 687200
rect 20 856 557476 687144
rect 20 800 514 856
rect 682 800 1618 856
rect 1786 800 2722 856
rect 2890 800 3918 856
rect 4086 800 5022 856
rect 5190 800 6126 856
rect 6294 800 7322 856
rect 7490 800 8426 856
rect 8594 800 9530 856
rect 9698 800 10726 856
rect 10894 800 11830 856
rect 11998 800 12934 856
rect 13102 800 14130 856
rect 14298 800 15234 856
rect 15402 800 16338 856
rect 16506 800 17534 856
rect 17702 800 18638 856
rect 18806 800 19742 856
rect 19910 800 20938 856
rect 21106 800 22042 856
rect 22210 800 23146 856
rect 23314 800 24342 856
rect 24510 800 25446 856
rect 25614 800 26642 856
rect 26810 800 27746 856
rect 27914 800 28850 856
rect 29018 800 30046 856
rect 30214 800 31150 856
rect 31318 800 32254 856
rect 32422 800 33450 856
rect 33618 800 34554 856
rect 34722 800 35658 856
rect 35826 800 36854 856
rect 37022 800 37958 856
rect 38126 800 39062 856
rect 39230 800 40258 856
rect 40426 800 41362 856
rect 41530 800 42466 856
rect 42634 800 43662 856
rect 43830 800 44766 856
rect 44934 800 45870 856
rect 46038 800 47066 856
rect 47234 800 48170 856
rect 48338 800 49274 856
rect 49442 800 50470 856
rect 50638 800 51574 856
rect 51742 800 52770 856
rect 52938 800 53874 856
rect 54042 800 54978 856
rect 55146 800 56174 856
rect 56342 800 57278 856
rect 57446 800 58382 856
rect 58550 800 59578 856
rect 59746 800 60682 856
rect 60850 800 61786 856
rect 61954 800 62982 856
rect 63150 800 64086 856
rect 64254 800 65190 856
rect 65358 800 66386 856
rect 66554 800 67490 856
rect 67658 800 68594 856
rect 68762 800 69790 856
rect 69958 800 70894 856
rect 71062 800 71998 856
rect 72166 800 73194 856
rect 73362 800 74298 856
rect 74466 800 75402 856
rect 75570 800 76598 856
rect 76766 800 77702 856
rect 77870 800 78898 856
rect 79066 800 80002 856
rect 80170 800 81106 856
rect 81274 800 82302 856
rect 82470 800 83406 856
rect 83574 800 84510 856
rect 84678 800 85706 856
rect 85874 800 86810 856
rect 86978 800 87914 856
rect 88082 800 89110 856
rect 89278 800 90214 856
rect 90382 800 91318 856
rect 91486 800 92514 856
rect 92682 800 93618 856
rect 93786 800 94722 856
rect 94890 800 95918 856
rect 96086 800 97022 856
rect 97190 800 98126 856
rect 98294 800 99322 856
rect 99490 800 100426 856
rect 100594 800 101530 856
rect 101698 800 102726 856
rect 102894 800 103830 856
rect 103998 800 105026 856
rect 105194 800 106130 856
rect 106298 800 107234 856
rect 107402 800 108430 856
rect 108598 800 109534 856
rect 109702 800 110638 856
rect 110806 800 111834 856
rect 112002 800 112938 856
rect 113106 800 114042 856
rect 114210 800 115238 856
rect 115406 800 116342 856
rect 116510 800 117446 856
rect 117614 800 118642 856
rect 118810 800 119746 856
rect 119914 800 120850 856
rect 121018 800 122046 856
rect 122214 800 123150 856
rect 123318 800 124254 856
rect 124422 800 125450 856
rect 125618 800 126554 856
rect 126722 800 127658 856
rect 127826 800 128854 856
rect 129022 800 129958 856
rect 130126 800 131154 856
rect 131322 800 132258 856
rect 132426 800 133362 856
rect 133530 800 134558 856
rect 134726 800 135662 856
rect 135830 800 136766 856
rect 136934 800 137962 856
rect 138130 800 139066 856
rect 139234 800 140170 856
rect 140338 800 141366 856
rect 141534 800 142470 856
rect 142638 800 143574 856
rect 143742 800 144770 856
rect 144938 800 145874 856
rect 146042 800 146978 856
rect 147146 800 148174 856
rect 148342 800 149278 856
rect 149446 800 150382 856
rect 150550 800 151578 856
rect 151746 800 152682 856
rect 152850 800 153786 856
rect 153954 800 154982 856
rect 155150 800 156086 856
rect 156254 800 157282 856
rect 157450 800 158386 856
rect 158554 800 159490 856
rect 159658 800 160686 856
rect 160854 800 161790 856
rect 161958 800 162894 856
rect 163062 800 164090 856
rect 164258 800 165194 856
rect 165362 800 166298 856
rect 166466 800 167494 856
rect 167662 800 168598 856
rect 168766 800 169702 856
rect 169870 800 170898 856
rect 171066 800 172002 856
rect 172170 800 173106 856
rect 173274 800 174302 856
rect 174470 800 175406 856
rect 175574 800 176510 856
rect 176678 800 177706 856
rect 177874 800 178810 856
rect 178978 800 179914 856
rect 180082 800 181110 856
rect 181278 800 182214 856
rect 182382 800 183410 856
rect 183578 800 184514 856
rect 184682 800 185618 856
rect 185786 800 186814 856
rect 186982 800 187918 856
rect 188086 800 189022 856
rect 189190 800 190218 856
rect 190386 800 191322 856
rect 191490 800 192426 856
rect 192594 800 193622 856
rect 193790 800 194726 856
rect 194894 800 195830 856
rect 195998 800 197026 856
rect 197194 800 198130 856
rect 198298 800 199234 856
rect 199402 800 200430 856
rect 200598 800 201534 856
rect 201702 800 202638 856
rect 202806 800 203834 856
rect 204002 800 204938 856
rect 205106 800 206042 856
rect 206210 800 207238 856
rect 207406 800 208342 856
rect 208510 800 209538 856
rect 209706 800 210642 856
rect 210810 800 211746 856
rect 211914 800 212942 856
rect 213110 800 214046 856
rect 214214 800 215150 856
rect 215318 800 216346 856
rect 216514 800 217450 856
rect 217618 800 218554 856
rect 218722 800 219750 856
rect 219918 800 220854 856
rect 221022 800 221958 856
rect 222126 800 223154 856
rect 223322 800 224258 856
rect 224426 800 225362 856
rect 225530 800 226558 856
rect 226726 800 227662 856
rect 227830 800 228766 856
rect 228934 800 229962 856
rect 230130 800 231066 856
rect 231234 800 232170 856
rect 232338 800 233366 856
rect 233534 800 234470 856
rect 234638 800 235666 856
rect 235834 800 236770 856
rect 236938 800 237874 856
rect 238042 800 239070 856
rect 239238 800 240174 856
rect 240342 800 241278 856
rect 241446 800 242474 856
rect 242642 800 243578 856
rect 243746 800 244682 856
rect 244850 800 245878 856
rect 246046 800 246982 856
rect 247150 800 248086 856
rect 248254 800 249282 856
rect 249450 800 250386 856
rect 250554 800 251490 856
rect 251658 800 252686 856
rect 252854 800 253790 856
rect 253958 800 254894 856
rect 255062 800 256090 856
rect 256258 800 257194 856
rect 257362 800 258298 856
rect 258466 800 259494 856
rect 259662 800 260598 856
rect 260766 800 261794 856
rect 261962 800 262898 856
rect 263066 800 264002 856
rect 264170 800 265198 856
rect 265366 800 266302 856
rect 266470 800 267406 856
rect 267574 800 268602 856
rect 268770 800 269706 856
rect 269874 800 270810 856
rect 270978 800 272006 856
rect 272174 800 273110 856
rect 273278 800 274214 856
rect 274382 800 275410 856
rect 275578 800 276514 856
rect 276682 800 277618 856
rect 277786 800 278814 856
rect 278982 800 279918 856
rect 280086 800 281022 856
rect 281190 800 282218 856
rect 282386 800 283322 856
rect 283490 800 284518 856
rect 284686 800 285622 856
rect 285790 800 286726 856
rect 286894 800 287922 856
rect 288090 800 289026 856
rect 289194 800 290130 856
rect 290298 800 291326 856
rect 291494 800 292430 856
rect 292598 800 293534 856
rect 293702 800 294730 856
rect 294898 800 295834 856
rect 296002 800 296938 856
rect 297106 800 298134 856
rect 298302 800 299238 856
rect 299406 800 300342 856
rect 300510 800 301538 856
rect 301706 800 302642 856
rect 302810 800 303746 856
rect 303914 800 304942 856
rect 305110 800 306046 856
rect 306214 800 307150 856
rect 307318 800 308346 856
rect 308514 800 309450 856
rect 309618 800 310646 856
rect 310814 800 311750 856
rect 311918 800 312854 856
rect 313022 800 314050 856
rect 314218 800 315154 856
rect 315322 800 316258 856
rect 316426 800 317454 856
rect 317622 800 318558 856
rect 318726 800 319662 856
rect 319830 800 320858 856
rect 321026 800 321962 856
rect 322130 800 323066 856
rect 323234 800 324262 856
rect 324430 800 325366 856
rect 325534 800 326470 856
rect 326638 800 327666 856
rect 327834 800 328770 856
rect 328938 800 329874 856
rect 330042 800 331070 856
rect 331238 800 332174 856
rect 332342 800 333278 856
rect 333446 800 334474 856
rect 334642 800 335578 856
rect 335746 800 336774 856
rect 336942 800 337878 856
rect 338046 800 338982 856
rect 339150 800 340178 856
rect 340346 800 341282 856
rect 341450 800 342386 856
rect 342554 800 343582 856
rect 343750 800 344686 856
rect 344854 800 345790 856
rect 345958 800 346986 856
rect 347154 800 348090 856
rect 348258 800 349194 856
rect 349362 800 350390 856
rect 350558 800 351494 856
rect 351662 800 352598 856
rect 352766 800 353794 856
rect 353962 800 354898 856
rect 355066 800 356002 856
rect 356170 800 357198 856
rect 357366 800 358302 856
rect 358470 800 359406 856
rect 359574 800 360602 856
rect 360770 800 361706 856
rect 361874 800 362902 856
rect 363070 800 364006 856
rect 364174 800 365110 856
rect 365278 800 366306 856
rect 366474 800 367410 856
rect 367578 800 368514 856
rect 368682 800 369710 856
rect 369878 800 370814 856
rect 370982 800 371918 856
rect 372086 800 373114 856
rect 373282 800 374218 856
rect 374386 800 375322 856
rect 375490 800 376518 856
rect 376686 800 377622 856
rect 377790 800 378726 856
rect 378894 800 379922 856
rect 380090 800 381026 856
rect 381194 800 382130 856
rect 382298 800 383326 856
rect 383494 800 384430 856
rect 384598 800 385534 856
rect 385702 800 386730 856
rect 386898 800 387834 856
rect 388002 800 389030 856
rect 389198 800 390134 856
rect 390302 800 391238 856
rect 391406 800 392434 856
rect 392602 800 393538 856
rect 393706 800 394642 856
rect 394810 800 395838 856
rect 396006 800 396942 856
rect 397110 800 398046 856
rect 398214 800 399242 856
rect 399410 800 400346 856
rect 400514 800 401450 856
rect 401618 800 402646 856
rect 402814 800 403750 856
rect 403918 800 404854 856
rect 405022 800 406050 856
rect 406218 800 407154 856
rect 407322 800 408258 856
rect 408426 800 409454 856
rect 409622 800 410558 856
rect 410726 800 411662 856
rect 411830 800 412858 856
rect 413026 800 413962 856
rect 414130 800 415158 856
rect 415326 800 416262 856
rect 416430 800 417366 856
rect 417534 800 418562 856
rect 418730 800 419666 856
rect 419834 800 420770 856
rect 420938 800 421966 856
rect 422134 800 423070 856
rect 423238 800 424174 856
rect 424342 800 425370 856
rect 425538 800 426474 856
rect 426642 800 427578 856
rect 427746 800 428774 856
rect 428942 800 429878 856
rect 430046 800 430982 856
rect 431150 800 432178 856
rect 432346 800 433282 856
rect 433450 800 434386 856
rect 434554 800 435582 856
rect 435750 800 436686 856
rect 436854 800 437790 856
rect 437958 800 438986 856
rect 439154 800 440090 856
rect 440258 800 441286 856
rect 441454 800 442390 856
rect 442558 800 443494 856
rect 443662 800 444690 856
rect 444858 800 445794 856
rect 445962 800 446898 856
rect 447066 800 448094 856
rect 448262 800 449198 856
rect 449366 800 450302 856
rect 450470 800 451498 856
rect 451666 800 452602 856
rect 452770 800 453706 856
rect 453874 800 454902 856
rect 455070 800 456006 856
rect 456174 800 457110 856
rect 457278 800 458306 856
rect 458474 800 459410 856
rect 459578 800 460514 856
rect 460682 800 461710 856
rect 461878 800 462814 856
rect 462982 800 463918 856
rect 464086 800 465114 856
rect 465282 800 466218 856
rect 466386 800 467414 856
rect 467582 800 468518 856
rect 468686 800 469622 856
rect 469790 800 470818 856
rect 470986 800 471922 856
rect 472090 800 473026 856
rect 473194 800 474222 856
rect 474390 800 475326 856
rect 475494 800 476430 856
rect 476598 800 477626 856
rect 477794 800 478730 856
rect 478898 800 479834 856
rect 480002 800 481030 856
rect 481198 800 482134 856
rect 482302 800 483238 856
rect 483406 800 484434 856
rect 484602 800 485538 856
rect 485706 800 486642 856
rect 486810 800 487838 856
rect 488006 800 488942 856
rect 489110 800 490046 856
rect 490214 800 491242 856
rect 491410 800 492346 856
rect 492514 800 493542 856
rect 493710 800 494646 856
rect 494814 800 495750 856
rect 495918 800 496946 856
rect 497114 800 498050 856
rect 498218 800 499154 856
rect 499322 800 500350 856
rect 500518 800 501454 856
rect 501622 800 502558 856
rect 502726 800 503754 856
rect 503922 800 504858 856
rect 505026 800 505962 856
rect 506130 800 507158 856
rect 507326 800 508262 856
rect 508430 800 509366 856
rect 509534 800 510562 856
rect 510730 800 511666 856
rect 511834 800 512770 856
rect 512938 800 513966 856
rect 514134 800 515070 856
rect 515238 800 516174 856
rect 516342 800 517370 856
rect 517538 800 518474 856
rect 518642 800 519670 856
rect 519838 800 520774 856
rect 520942 800 521878 856
rect 522046 800 523074 856
rect 523242 800 524178 856
rect 524346 800 525282 856
rect 525450 800 526478 856
rect 526646 800 527582 856
rect 527750 800 528686 856
rect 528854 800 529882 856
rect 530050 800 530986 856
rect 531154 800 532090 856
rect 532258 800 533286 856
rect 533454 800 534390 856
rect 534558 800 535494 856
rect 535662 800 536690 856
rect 536858 800 537794 856
rect 537962 800 538898 856
rect 539066 800 540094 856
rect 540262 800 541198 856
rect 541366 800 542302 856
rect 542470 800 543498 856
rect 543666 800 544602 856
rect 544770 800 545798 856
rect 545966 800 546902 856
rect 547070 800 548006 856
rect 548174 800 549202 856
rect 549370 800 550306 856
rect 550474 800 551410 856
rect 551578 800 552606 856
rect 552774 800 553710 856
rect 553878 800 554814 856
rect 554982 800 556010 856
rect 556178 800 557114 856
rect 557282 800 557476 856
<< metal3 >>
rect 0 619080 800 619200
rect 0 481448 800 481568
rect 0 343816 800 343936
rect 0 206184 800 206304
rect 0 68688 800 68808
rect 567200 644920 568000 645040
rect 567200 558968 568000 559088
rect 567200 472880 568000 473000
rect 567200 386928 568000 387048
rect 567200 300976 568000 301096
rect 567200 214888 568000 215008
rect 567200 128936 568000 129056
rect 567200 42984 568000 43104
<< obsm3 >>
rect 1669 2143 557488 685473
<< metal4 >>
rect 4208 2128 4528 685488
rect 19568 2128 19888 685488
rect 34928 2128 35248 685488
rect 50288 2128 50608 685488
rect 65648 2128 65968 685488
rect 81008 2128 81328 685488
rect 96368 2128 96688 685488
rect 111728 2128 112048 685488
rect 127088 2128 127408 685488
rect 142448 2128 142768 685488
rect 157808 2128 158128 685488
rect 173168 2128 173488 685488
rect 188528 2128 188848 685488
rect 203888 2128 204208 685488
rect 219248 2128 219568 685488
rect 234608 2128 234928 685488
rect 249968 2128 250288 685488
rect 265328 2128 265648 685488
rect 280688 2128 281008 685488
rect 296048 2128 296368 685488
rect 311408 2128 311728 685488
rect 326768 2128 327088 685488
rect 342128 2128 342448 685488
rect 357488 2128 357808 685488
rect 372848 2128 373168 685488
rect 388208 2128 388528 685488
rect 403568 2128 403888 685488
rect 418928 2128 419248 685488
rect 434288 2128 434608 685488
rect 449648 2128 449968 685488
rect 465008 2128 465328 685488
rect 480368 2128 480688 685488
rect 495728 2128 496048 685488
rect 511088 2128 511408 685488
rect 526448 2128 526768 685488
rect 541808 2128 542128 685488
rect 557168 2128 557488 685488
<< obsm4 >>
rect 3555 3435 4128 680645
rect 4608 3435 19488 680645
rect 19968 3435 34848 680645
rect 35328 3435 50208 680645
rect 50688 3435 65568 680645
rect 66048 3435 80928 680645
rect 81408 3435 96288 680645
rect 96768 3435 111648 680645
rect 112128 3435 127008 680645
rect 127488 3435 142368 680645
rect 142848 3435 157728 680645
rect 158208 3435 173088 680645
rect 173568 3435 188448 680645
rect 188928 3435 203808 680645
rect 204288 3435 219168 680645
rect 219648 3435 234528 680645
rect 235008 3435 249888 680645
rect 250368 3435 265248 680645
rect 265728 3435 280608 680645
rect 281088 3435 295968 680645
rect 296448 3435 311328 680645
rect 311808 3435 326688 680645
rect 327168 3435 342048 680645
rect 342528 3435 357408 680645
rect 357888 3435 372768 680645
rect 373248 3435 388128 680645
rect 388608 3435 403488 680645
rect 403968 3435 418848 680645
rect 419328 3435 434208 680645
rect 434688 3435 449568 680645
rect 450048 3435 464928 680645
rect 465408 3435 480288 680645
rect 480768 3435 495648 680645
rect 496128 3435 511008 680645
rect 511488 3435 526368 680645
rect 526848 3435 541728 680645
rect 542208 3435 550285 680645
<< labels >>
rlabel metal3 s 0 68688 800 68808 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal3 s 567200 128936 568000 129056 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 547234 687200 547290 688000 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 551834 687200 551890 688000 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal3 s 0 343816 800 343936 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 556434 687200 556490 688000 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 561678 0 561734 800 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal3 s 567200 214888 568000 215008 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s 0 481448 800 481568 6 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal2 s 562874 0 562930 800 6 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal2 s 561034 687200 561090 688000 6 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal2 s 558274 0 558330 800 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s 0 619080 800 619200 6 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s 567200 300976 568000 301096 6 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal2 s 565634 687200 565690 688000 6 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s 567200 386928 568000 387048 6 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal2 s 563978 0 564034 800 6 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal2 s 565082 0 565138 800 6 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal2 s 566278 0 566334 800 6 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s 567200 472880 568000 473000 6 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s 567200 558968 568000 559088 6 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 567200 644920 568000 645040 6 analog_io[29]
port 22 nsew signal bidirectional
rlabel metal2 s 528742 687200 528798 688000 6 analog_io[2]
port 23 nsew signal bidirectional
rlabel metal2 s 567382 0 567438 800 6 analog_io[30]
port 24 nsew signal bidirectional
rlabel metal2 s 533342 687200 533398 688000 6 analog_io[3]
port 25 nsew signal bidirectional
rlabel metal3 s 0 206184 800 206304 6 analog_io[4]
port 26 nsew signal bidirectional
rlabel metal2 s 537942 687200 537998 688000 6 analog_io[5]
port 27 nsew signal bidirectional
rlabel metal2 s 559470 0 559526 800 6 analog_io[6]
port 28 nsew signal bidirectional
rlabel metal2 s 542542 687200 542598 688000 6 analog_io[7]
port 29 nsew signal bidirectional
rlabel metal3 s 567200 42984 568000 43104 6 analog_io[8]
port 30 nsew signal bidirectional
rlabel metal2 s 560574 0 560630 800 6 analog_io[9]
port 31 nsew signal bidirectional
rlabel metal2 s 2318 687200 2374 688000 6 io_in[0]
port 32 nsew signal input
rlabel metal2 s 140778 687200 140834 688000 6 io_in[10]
port 33 nsew signal input
rlabel metal2 s 154670 687200 154726 688000 6 io_in[11]
port 34 nsew signal input
rlabel metal2 s 168562 687200 168618 688000 6 io_in[12]
port 35 nsew signal input
rlabel metal2 s 182362 687200 182418 688000 6 io_in[13]
port 36 nsew signal input
rlabel metal2 s 196254 687200 196310 688000 6 io_in[14]
port 37 nsew signal input
rlabel metal2 s 210054 687200 210110 688000 6 io_in[15]
port 38 nsew signal input
rlabel metal2 s 223946 687200 224002 688000 6 io_in[16]
port 39 nsew signal input
rlabel metal2 s 237746 687200 237802 688000 6 io_in[17]
port 40 nsew signal input
rlabel metal2 s 251638 687200 251694 688000 6 io_in[18]
port 41 nsew signal input
rlabel metal2 s 265530 687200 265586 688000 6 io_in[19]
port 42 nsew signal input
rlabel metal2 s 16118 687200 16174 688000 6 io_in[1]
port 43 nsew signal input
rlabel metal2 s 279330 687200 279386 688000 6 io_in[20]
port 44 nsew signal input
rlabel metal2 s 293222 687200 293278 688000 6 io_in[21]
port 45 nsew signal input
rlabel metal2 s 307022 687200 307078 688000 6 io_in[22]
port 46 nsew signal input
rlabel metal2 s 320914 687200 320970 688000 6 io_in[23]
port 47 nsew signal input
rlabel metal2 s 334806 687200 334862 688000 6 io_in[24]
port 48 nsew signal input
rlabel metal2 s 348606 687200 348662 688000 6 io_in[25]
port 49 nsew signal input
rlabel metal2 s 362498 687200 362554 688000 6 io_in[26]
port 50 nsew signal input
rlabel metal2 s 376298 687200 376354 688000 6 io_in[27]
port 51 nsew signal input
rlabel metal2 s 390190 687200 390246 688000 6 io_in[28]
port 52 nsew signal input
rlabel metal2 s 403990 687200 404046 688000 6 io_in[29]
port 53 nsew signal input
rlabel metal2 s 30010 687200 30066 688000 6 io_in[2]
port 54 nsew signal input
rlabel metal2 s 417882 687200 417938 688000 6 io_in[30]
port 55 nsew signal input
rlabel metal2 s 431774 687200 431830 688000 6 io_in[31]
port 56 nsew signal input
rlabel metal2 s 445574 687200 445630 688000 6 io_in[32]
port 57 nsew signal input
rlabel metal2 s 459466 687200 459522 688000 6 io_in[33]
port 58 nsew signal input
rlabel metal2 s 473266 687200 473322 688000 6 io_in[34]
port 59 nsew signal input
rlabel metal2 s 487158 687200 487214 688000 6 io_in[35]
port 60 nsew signal input
rlabel metal2 s 501050 687200 501106 688000 6 io_in[36]
port 61 nsew signal input
rlabel metal2 s 514850 687200 514906 688000 6 io_in[37]
port 62 nsew signal input
rlabel metal2 s 43810 687200 43866 688000 6 io_in[3]
port 63 nsew signal input
rlabel metal2 s 57702 687200 57758 688000 6 io_in[4]
port 64 nsew signal input
rlabel metal2 s 71502 687200 71558 688000 6 io_in[5]
port 65 nsew signal input
rlabel metal2 s 85394 687200 85450 688000 6 io_in[6]
port 66 nsew signal input
rlabel metal2 s 99286 687200 99342 688000 6 io_in[7]
port 67 nsew signal input
rlabel metal2 s 113086 687200 113142 688000 6 io_in[8]
port 68 nsew signal input
rlabel metal2 s 126978 687200 127034 688000 6 io_in[9]
port 69 nsew signal input
rlabel metal2 s 6918 687200 6974 688000 6 io_oeb[0]
port 70 nsew signal output
rlabel metal2 s 145470 687200 145526 688000 6 io_oeb[10]
port 71 nsew signal output
rlabel metal2 s 159270 687200 159326 688000 6 io_oeb[11]
port 72 nsew signal output
rlabel metal2 s 173162 687200 173218 688000 6 io_oeb[12]
port 73 nsew signal output
rlabel metal2 s 186962 687200 187018 688000 6 io_oeb[13]
port 74 nsew signal output
rlabel metal2 s 200854 687200 200910 688000 6 io_oeb[14]
port 75 nsew signal output
rlabel metal2 s 214654 687200 214710 688000 6 io_oeb[15]
port 76 nsew signal output
rlabel metal2 s 228546 687200 228602 688000 6 io_oeb[16]
port 77 nsew signal output
rlabel metal2 s 242438 687200 242494 688000 6 io_oeb[17]
port 78 nsew signal output
rlabel metal2 s 256238 687200 256294 688000 6 io_oeb[18]
port 79 nsew signal output
rlabel metal2 s 270130 687200 270186 688000 6 io_oeb[19]
port 80 nsew signal output
rlabel metal2 s 20718 687200 20774 688000 6 io_oeb[1]
port 81 nsew signal output
rlabel metal2 s 283930 687200 283986 688000 6 io_oeb[20]
port 82 nsew signal output
rlabel metal2 s 297822 687200 297878 688000 6 io_oeb[21]
port 83 nsew signal output
rlabel metal2 s 311714 687200 311770 688000 6 io_oeb[22]
port 84 nsew signal output
rlabel metal2 s 325514 687200 325570 688000 6 io_oeb[23]
port 85 nsew signal output
rlabel metal2 s 339406 687200 339462 688000 6 io_oeb[24]
port 86 nsew signal output
rlabel metal2 s 353206 687200 353262 688000 6 io_oeb[25]
port 87 nsew signal output
rlabel metal2 s 367098 687200 367154 688000 6 io_oeb[26]
port 88 nsew signal output
rlabel metal2 s 380990 687200 381046 688000 6 io_oeb[27]
port 89 nsew signal output
rlabel metal2 s 394790 687200 394846 688000 6 io_oeb[28]
port 90 nsew signal output
rlabel metal2 s 408682 687200 408738 688000 6 io_oeb[29]
port 91 nsew signal output
rlabel metal2 s 34610 687200 34666 688000 6 io_oeb[2]
port 92 nsew signal output
rlabel metal2 s 422482 687200 422538 688000 6 io_oeb[30]
port 93 nsew signal output
rlabel metal2 s 436374 687200 436430 688000 6 io_oeb[31]
port 94 nsew signal output
rlabel metal2 s 450174 687200 450230 688000 6 io_oeb[32]
port 95 nsew signal output
rlabel metal2 s 464066 687200 464122 688000 6 io_oeb[33]
port 96 nsew signal output
rlabel metal2 s 477958 687200 478014 688000 6 io_oeb[34]
port 97 nsew signal output
rlabel metal2 s 491758 687200 491814 688000 6 io_oeb[35]
port 98 nsew signal output
rlabel metal2 s 505650 687200 505706 688000 6 io_oeb[36]
port 99 nsew signal output
rlabel metal2 s 519450 687200 519506 688000 6 io_oeb[37]
port 100 nsew signal output
rlabel metal2 s 48410 687200 48466 688000 6 io_oeb[3]
port 101 nsew signal output
rlabel metal2 s 62302 687200 62358 688000 6 io_oeb[4]
port 102 nsew signal output
rlabel metal2 s 76194 687200 76250 688000 6 io_oeb[5]
port 103 nsew signal output
rlabel metal2 s 89994 687200 90050 688000 6 io_oeb[6]
port 104 nsew signal output
rlabel metal2 s 103886 687200 103942 688000 6 io_oeb[7]
port 105 nsew signal output
rlabel metal2 s 117686 687200 117742 688000 6 io_oeb[8]
port 106 nsew signal output
rlabel metal2 s 131578 687200 131634 688000 6 io_oeb[9]
port 107 nsew signal output
rlabel metal2 s 11518 687200 11574 688000 6 io_out[0]
port 108 nsew signal output
rlabel metal2 s 150070 687200 150126 688000 6 io_out[10]
port 109 nsew signal output
rlabel metal2 s 163870 687200 163926 688000 6 io_out[11]
port 110 nsew signal output
rlabel metal2 s 177762 687200 177818 688000 6 io_out[12]
port 111 nsew signal output
rlabel metal2 s 191654 687200 191710 688000 6 io_out[13]
port 112 nsew signal output
rlabel metal2 s 205454 687200 205510 688000 6 io_out[14]
port 113 nsew signal output
rlabel metal2 s 219346 687200 219402 688000 6 io_out[15]
port 114 nsew signal output
rlabel metal2 s 233146 687200 233202 688000 6 io_out[16]
port 115 nsew signal output
rlabel metal2 s 247038 687200 247094 688000 6 io_out[17]
port 116 nsew signal output
rlabel metal2 s 260838 687200 260894 688000 6 io_out[18]
port 117 nsew signal output
rlabel metal2 s 274730 687200 274786 688000 6 io_out[19]
port 118 nsew signal output
rlabel metal2 s 25318 687200 25374 688000 6 io_out[1]
port 119 nsew signal output
rlabel metal2 s 288622 687200 288678 688000 6 io_out[20]
port 120 nsew signal output
rlabel metal2 s 302422 687200 302478 688000 6 io_out[21]
port 121 nsew signal output
rlabel metal2 s 316314 687200 316370 688000 6 io_out[22]
port 122 nsew signal output
rlabel metal2 s 330114 687200 330170 688000 6 io_out[23]
port 123 nsew signal output
rlabel metal2 s 344006 687200 344062 688000 6 io_out[24]
port 124 nsew signal output
rlabel metal2 s 357898 687200 357954 688000 6 io_out[25]
port 125 nsew signal output
rlabel metal2 s 371698 687200 371754 688000 6 io_out[26]
port 126 nsew signal output
rlabel metal2 s 385590 687200 385646 688000 6 io_out[27]
port 127 nsew signal output
rlabel metal2 s 399390 687200 399446 688000 6 io_out[28]
port 128 nsew signal output
rlabel metal2 s 413282 687200 413338 688000 6 io_out[29]
port 129 nsew signal output
rlabel metal2 s 39210 687200 39266 688000 6 io_out[2]
port 130 nsew signal output
rlabel metal2 s 427082 687200 427138 688000 6 io_out[30]
port 131 nsew signal output
rlabel metal2 s 440974 687200 441030 688000 6 io_out[31]
port 132 nsew signal output
rlabel metal2 s 454866 687200 454922 688000 6 io_out[32]
port 133 nsew signal output
rlabel metal2 s 468666 687200 468722 688000 6 io_out[33]
port 134 nsew signal output
rlabel metal2 s 482558 687200 482614 688000 6 io_out[34]
port 135 nsew signal output
rlabel metal2 s 496358 687200 496414 688000 6 io_out[35]
port 136 nsew signal output
rlabel metal2 s 510250 687200 510306 688000 6 io_out[36]
port 137 nsew signal output
rlabel metal2 s 524142 687200 524198 688000 6 io_out[37]
port 138 nsew signal output
rlabel metal2 s 53102 687200 53158 688000 6 io_out[3]
port 139 nsew signal output
rlabel metal2 s 66902 687200 66958 688000 6 io_out[4]
port 140 nsew signal output
rlabel metal2 s 80794 687200 80850 688000 6 io_out[5]
port 141 nsew signal output
rlabel metal2 s 94594 687200 94650 688000 6 io_out[6]
port 142 nsew signal output
rlabel metal2 s 108486 687200 108542 688000 6 io_out[7]
port 143 nsew signal output
rlabel metal2 s 122378 687200 122434 688000 6 io_out[8]
port 144 nsew signal output
rlabel metal2 s 136178 687200 136234 688000 6 io_out[9]
port 145 nsew signal output
rlabel metal2 s 120906 0 120962 800 6 la_data_in[0]
port 146 nsew signal input
rlabel metal2 s 461766 0 461822 800 6 la_data_in[100]
port 147 nsew signal input
rlabel metal2 s 465170 0 465226 800 6 la_data_in[101]
port 148 nsew signal input
rlabel metal2 s 468574 0 468630 800 6 la_data_in[102]
port 149 nsew signal input
rlabel metal2 s 471978 0 472034 800 6 la_data_in[103]
port 150 nsew signal input
rlabel metal2 s 475382 0 475438 800 6 la_data_in[104]
port 151 nsew signal input
rlabel metal2 s 478786 0 478842 800 6 la_data_in[105]
port 152 nsew signal input
rlabel metal2 s 482190 0 482246 800 6 la_data_in[106]
port 153 nsew signal input
rlabel metal2 s 485594 0 485650 800 6 la_data_in[107]
port 154 nsew signal input
rlabel metal2 s 488998 0 489054 800 6 la_data_in[108]
port 155 nsew signal input
rlabel metal2 s 492402 0 492458 800 6 la_data_in[109]
port 156 nsew signal input
rlabel metal2 s 155038 0 155094 800 6 la_data_in[10]
port 157 nsew signal input
rlabel metal2 s 495806 0 495862 800 6 la_data_in[110]
port 158 nsew signal input
rlabel metal2 s 499210 0 499266 800 6 la_data_in[111]
port 159 nsew signal input
rlabel metal2 s 502614 0 502670 800 6 la_data_in[112]
port 160 nsew signal input
rlabel metal2 s 506018 0 506074 800 6 la_data_in[113]
port 161 nsew signal input
rlabel metal2 s 509422 0 509478 800 6 la_data_in[114]
port 162 nsew signal input
rlabel metal2 s 512826 0 512882 800 6 la_data_in[115]
port 163 nsew signal input
rlabel metal2 s 516230 0 516286 800 6 la_data_in[116]
port 164 nsew signal input
rlabel metal2 s 519726 0 519782 800 6 la_data_in[117]
port 165 nsew signal input
rlabel metal2 s 523130 0 523186 800 6 la_data_in[118]
port 166 nsew signal input
rlabel metal2 s 526534 0 526590 800 6 la_data_in[119]
port 167 nsew signal input
rlabel metal2 s 158442 0 158498 800 6 la_data_in[11]
port 168 nsew signal input
rlabel metal2 s 529938 0 529994 800 6 la_data_in[120]
port 169 nsew signal input
rlabel metal2 s 533342 0 533398 800 6 la_data_in[121]
port 170 nsew signal input
rlabel metal2 s 536746 0 536802 800 6 la_data_in[122]
port 171 nsew signal input
rlabel metal2 s 540150 0 540206 800 6 la_data_in[123]
port 172 nsew signal input
rlabel metal2 s 543554 0 543610 800 6 la_data_in[124]
port 173 nsew signal input
rlabel metal2 s 546958 0 547014 800 6 la_data_in[125]
port 174 nsew signal input
rlabel metal2 s 550362 0 550418 800 6 la_data_in[126]
port 175 nsew signal input
rlabel metal2 s 553766 0 553822 800 6 la_data_in[127]
port 176 nsew signal input
rlabel metal2 s 161846 0 161902 800 6 la_data_in[12]
port 177 nsew signal input
rlabel metal2 s 165250 0 165306 800 6 la_data_in[13]
port 178 nsew signal input
rlabel metal2 s 168654 0 168710 800 6 la_data_in[14]
port 179 nsew signal input
rlabel metal2 s 172058 0 172114 800 6 la_data_in[15]
port 180 nsew signal input
rlabel metal2 s 175462 0 175518 800 6 la_data_in[16]
port 181 nsew signal input
rlabel metal2 s 178866 0 178922 800 6 la_data_in[17]
port 182 nsew signal input
rlabel metal2 s 182270 0 182326 800 6 la_data_in[18]
port 183 nsew signal input
rlabel metal2 s 185674 0 185730 800 6 la_data_in[19]
port 184 nsew signal input
rlabel metal2 s 124310 0 124366 800 6 la_data_in[1]
port 185 nsew signal input
rlabel metal2 s 189078 0 189134 800 6 la_data_in[20]
port 186 nsew signal input
rlabel metal2 s 192482 0 192538 800 6 la_data_in[21]
port 187 nsew signal input
rlabel metal2 s 195886 0 195942 800 6 la_data_in[22]
port 188 nsew signal input
rlabel metal2 s 199290 0 199346 800 6 la_data_in[23]
port 189 nsew signal input
rlabel metal2 s 202694 0 202750 800 6 la_data_in[24]
port 190 nsew signal input
rlabel metal2 s 206098 0 206154 800 6 la_data_in[25]
port 191 nsew signal input
rlabel metal2 s 209594 0 209650 800 6 la_data_in[26]
port 192 nsew signal input
rlabel metal2 s 212998 0 213054 800 6 la_data_in[27]
port 193 nsew signal input
rlabel metal2 s 216402 0 216458 800 6 la_data_in[28]
port 194 nsew signal input
rlabel metal2 s 219806 0 219862 800 6 la_data_in[29]
port 195 nsew signal input
rlabel metal2 s 127714 0 127770 800 6 la_data_in[2]
port 196 nsew signal input
rlabel metal2 s 223210 0 223266 800 6 la_data_in[30]
port 197 nsew signal input
rlabel metal2 s 226614 0 226670 800 6 la_data_in[31]
port 198 nsew signal input
rlabel metal2 s 230018 0 230074 800 6 la_data_in[32]
port 199 nsew signal input
rlabel metal2 s 233422 0 233478 800 6 la_data_in[33]
port 200 nsew signal input
rlabel metal2 s 236826 0 236882 800 6 la_data_in[34]
port 201 nsew signal input
rlabel metal2 s 240230 0 240286 800 6 la_data_in[35]
port 202 nsew signal input
rlabel metal2 s 243634 0 243690 800 6 la_data_in[36]
port 203 nsew signal input
rlabel metal2 s 247038 0 247094 800 6 la_data_in[37]
port 204 nsew signal input
rlabel metal2 s 250442 0 250498 800 6 la_data_in[38]
port 205 nsew signal input
rlabel metal2 s 253846 0 253902 800 6 la_data_in[39]
port 206 nsew signal input
rlabel metal2 s 131210 0 131266 800 6 la_data_in[3]
port 207 nsew signal input
rlabel metal2 s 257250 0 257306 800 6 la_data_in[40]
port 208 nsew signal input
rlabel metal2 s 260654 0 260710 800 6 la_data_in[41]
port 209 nsew signal input
rlabel metal2 s 264058 0 264114 800 6 la_data_in[42]
port 210 nsew signal input
rlabel metal2 s 267462 0 267518 800 6 la_data_in[43]
port 211 nsew signal input
rlabel metal2 s 270866 0 270922 800 6 la_data_in[44]
port 212 nsew signal input
rlabel metal2 s 274270 0 274326 800 6 la_data_in[45]
port 213 nsew signal input
rlabel metal2 s 277674 0 277730 800 6 la_data_in[46]
port 214 nsew signal input
rlabel metal2 s 281078 0 281134 800 6 la_data_in[47]
port 215 nsew signal input
rlabel metal2 s 284574 0 284630 800 6 la_data_in[48]
port 216 nsew signal input
rlabel metal2 s 287978 0 288034 800 6 la_data_in[49]
port 217 nsew signal input
rlabel metal2 s 134614 0 134670 800 6 la_data_in[4]
port 218 nsew signal input
rlabel metal2 s 291382 0 291438 800 6 la_data_in[50]
port 219 nsew signal input
rlabel metal2 s 294786 0 294842 800 6 la_data_in[51]
port 220 nsew signal input
rlabel metal2 s 298190 0 298246 800 6 la_data_in[52]
port 221 nsew signal input
rlabel metal2 s 301594 0 301650 800 6 la_data_in[53]
port 222 nsew signal input
rlabel metal2 s 304998 0 305054 800 6 la_data_in[54]
port 223 nsew signal input
rlabel metal2 s 308402 0 308458 800 6 la_data_in[55]
port 224 nsew signal input
rlabel metal2 s 311806 0 311862 800 6 la_data_in[56]
port 225 nsew signal input
rlabel metal2 s 315210 0 315266 800 6 la_data_in[57]
port 226 nsew signal input
rlabel metal2 s 318614 0 318670 800 6 la_data_in[58]
port 227 nsew signal input
rlabel metal2 s 322018 0 322074 800 6 la_data_in[59]
port 228 nsew signal input
rlabel metal2 s 138018 0 138074 800 6 la_data_in[5]
port 229 nsew signal input
rlabel metal2 s 325422 0 325478 800 6 la_data_in[60]
port 230 nsew signal input
rlabel metal2 s 328826 0 328882 800 6 la_data_in[61]
port 231 nsew signal input
rlabel metal2 s 332230 0 332286 800 6 la_data_in[62]
port 232 nsew signal input
rlabel metal2 s 335634 0 335690 800 6 la_data_in[63]
port 233 nsew signal input
rlabel metal2 s 339038 0 339094 800 6 la_data_in[64]
port 234 nsew signal input
rlabel metal2 s 342442 0 342498 800 6 la_data_in[65]
port 235 nsew signal input
rlabel metal2 s 345846 0 345902 800 6 la_data_in[66]
port 236 nsew signal input
rlabel metal2 s 349250 0 349306 800 6 la_data_in[67]
port 237 nsew signal input
rlabel metal2 s 352654 0 352710 800 6 la_data_in[68]
port 238 nsew signal input
rlabel metal2 s 356058 0 356114 800 6 la_data_in[69]
port 239 nsew signal input
rlabel metal2 s 141422 0 141478 800 6 la_data_in[6]
port 240 nsew signal input
rlabel metal2 s 359462 0 359518 800 6 la_data_in[70]
port 241 nsew signal input
rlabel metal2 s 362958 0 363014 800 6 la_data_in[71]
port 242 nsew signal input
rlabel metal2 s 366362 0 366418 800 6 la_data_in[72]
port 243 nsew signal input
rlabel metal2 s 369766 0 369822 800 6 la_data_in[73]
port 244 nsew signal input
rlabel metal2 s 373170 0 373226 800 6 la_data_in[74]
port 245 nsew signal input
rlabel metal2 s 376574 0 376630 800 6 la_data_in[75]
port 246 nsew signal input
rlabel metal2 s 379978 0 380034 800 6 la_data_in[76]
port 247 nsew signal input
rlabel metal2 s 383382 0 383438 800 6 la_data_in[77]
port 248 nsew signal input
rlabel metal2 s 386786 0 386842 800 6 la_data_in[78]
port 249 nsew signal input
rlabel metal2 s 390190 0 390246 800 6 la_data_in[79]
port 250 nsew signal input
rlabel metal2 s 144826 0 144882 800 6 la_data_in[7]
port 251 nsew signal input
rlabel metal2 s 393594 0 393650 800 6 la_data_in[80]
port 252 nsew signal input
rlabel metal2 s 396998 0 397054 800 6 la_data_in[81]
port 253 nsew signal input
rlabel metal2 s 400402 0 400458 800 6 la_data_in[82]
port 254 nsew signal input
rlabel metal2 s 403806 0 403862 800 6 la_data_in[83]
port 255 nsew signal input
rlabel metal2 s 407210 0 407266 800 6 la_data_in[84]
port 256 nsew signal input
rlabel metal2 s 410614 0 410670 800 6 la_data_in[85]
port 257 nsew signal input
rlabel metal2 s 414018 0 414074 800 6 la_data_in[86]
port 258 nsew signal input
rlabel metal2 s 417422 0 417478 800 6 la_data_in[87]
port 259 nsew signal input
rlabel metal2 s 420826 0 420882 800 6 la_data_in[88]
port 260 nsew signal input
rlabel metal2 s 424230 0 424286 800 6 la_data_in[89]
port 261 nsew signal input
rlabel metal2 s 148230 0 148286 800 6 la_data_in[8]
port 262 nsew signal input
rlabel metal2 s 427634 0 427690 800 6 la_data_in[90]
port 263 nsew signal input
rlabel metal2 s 431038 0 431094 800 6 la_data_in[91]
port 264 nsew signal input
rlabel metal2 s 434442 0 434498 800 6 la_data_in[92]
port 265 nsew signal input
rlabel metal2 s 437846 0 437902 800 6 la_data_in[93]
port 266 nsew signal input
rlabel metal2 s 441342 0 441398 800 6 la_data_in[94]
port 267 nsew signal input
rlabel metal2 s 444746 0 444802 800 6 la_data_in[95]
port 268 nsew signal input
rlabel metal2 s 448150 0 448206 800 6 la_data_in[96]
port 269 nsew signal input
rlabel metal2 s 451554 0 451610 800 6 la_data_in[97]
port 270 nsew signal input
rlabel metal2 s 454958 0 455014 800 6 la_data_in[98]
port 271 nsew signal input
rlabel metal2 s 458362 0 458418 800 6 la_data_in[99]
port 272 nsew signal input
rlabel metal2 s 151634 0 151690 800 6 la_data_in[9]
port 273 nsew signal input
rlabel metal2 s 122102 0 122158 800 6 la_data_out[0]
port 274 nsew signal output
rlabel metal2 s 462870 0 462926 800 6 la_data_out[100]
port 275 nsew signal output
rlabel metal2 s 466274 0 466330 800 6 la_data_out[101]
port 276 nsew signal output
rlabel metal2 s 469678 0 469734 800 6 la_data_out[102]
port 277 nsew signal output
rlabel metal2 s 473082 0 473138 800 6 la_data_out[103]
port 278 nsew signal output
rlabel metal2 s 476486 0 476542 800 6 la_data_out[104]
port 279 nsew signal output
rlabel metal2 s 479890 0 479946 800 6 la_data_out[105]
port 280 nsew signal output
rlabel metal2 s 483294 0 483350 800 6 la_data_out[106]
port 281 nsew signal output
rlabel metal2 s 486698 0 486754 800 6 la_data_out[107]
port 282 nsew signal output
rlabel metal2 s 490102 0 490158 800 6 la_data_out[108]
port 283 nsew signal output
rlabel metal2 s 493598 0 493654 800 6 la_data_out[109]
port 284 nsew signal output
rlabel metal2 s 156142 0 156198 800 6 la_data_out[10]
port 285 nsew signal output
rlabel metal2 s 497002 0 497058 800 6 la_data_out[110]
port 286 nsew signal output
rlabel metal2 s 500406 0 500462 800 6 la_data_out[111]
port 287 nsew signal output
rlabel metal2 s 503810 0 503866 800 6 la_data_out[112]
port 288 nsew signal output
rlabel metal2 s 507214 0 507270 800 6 la_data_out[113]
port 289 nsew signal output
rlabel metal2 s 510618 0 510674 800 6 la_data_out[114]
port 290 nsew signal output
rlabel metal2 s 514022 0 514078 800 6 la_data_out[115]
port 291 nsew signal output
rlabel metal2 s 517426 0 517482 800 6 la_data_out[116]
port 292 nsew signal output
rlabel metal2 s 520830 0 520886 800 6 la_data_out[117]
port 293 nsew signal output
rlabel metal2 s 524234 0 524290 800 6 la_data_out[118]
port 294 nsew signal output
rlabel metal2 s 527638 0 527694 800 6 la_data_out[119]
port 295 nsew signal output
rlabel metal2 s 159546 0 159602 800 6 la_data_out[11]
port 296 nsew signal output
rlabel metal2 s 531042 0 531098 800 6 la_data_out[120]
port 297 nsew signal output
rlabel metal2 s 534446 0 534502 800 6 la_data_out[121]
port 298 nsew signal output
rlabel metal2 s 537850 0 537906 800 6 la_data_out[122]
port 299 nsew signal output
rlabel metal2 s 541254 0 541310 800 6 la_data_out[123]
port 300 nsew signal output
rlabel metal2 s 544658 0 544714 800 6 la_data_out[124]
port 301 nsew signal output
rlabel metal2 s 548062 0 548118 800 6 la_data_out[125]
port 302 nsew signal output
rlabel metal2 s 551466 0 551522 800 6 la_data_out[126]
port 303 nsew signal output
rlabel metal2 s 554870 0 554926 800 6 la_data_out[127]
port 304 nsew signal output
rlabel metal2 s 162950 0 163006 800 6 la_data_out[12]
port 305 nsew signal output
rlabel metal2 s 166354 0 166410 800 6 la_data_out[13]
port 306 nsew signal output
rlabel metal2 s 169758 0 169814 800 6 la_data_out[14]
port 307 nsew signal output
rlabel metal2 s 173162 0 173218 800 6 la_data_out[15]
port 308 nsew signal output
rlabel metal2 s 176566 0 176622 800 6 la_data_out[16]
port 309 nsew signal output
rlabel metal2 s 179970 0 180026 800 6 la_data_out[17]
port 310 nsew signal output
rlabel metal2 s 183466 0 183522 800 6 la_data_out[18]
port 311 nsew signal output
rlabel metal2 s 186870 0 186926 800 6 la_data_out[19]
port 312 nsew signal output
rlabel metal2 s 125506 0 125562 800 6 la_data_out[1]
port 313 nsew signal output
rlabel metal2 s 190274 0 190330 800 6 la_data_out[20]
port 314 nsew signal output
rlabel metal2 s 193678 0 193734 800 6 la_data_out[21]
port 315 nsew signal output
rlabel metal2 s 197082 0 197138 800 6 la_data_out[22]
port 316 nsew signal output
rlabel metal2 s 200486 0 200542 800 6 la_data_out[23]
port 317 nsew signal output
rlabel metal2 s 203890 0 203946 800 6 la_data_out[24]
port 318 nsew signal output
rlabel metal2 s 207294 0 207350 800 6 la_data_out[25]
port 319 nsew signal output
rlabel metal2 s 210698 0 210754 800 6 la_data_out[26]
port 320 nsew signal output
rlabel metal2 s 214102 0 214158 800 6 la_data_out[27]
port 321 nsew signal output
rlabel metal2 s 217506 0 217562 800 6 la_data_out[28]
port 322 nsew signal output
rlabel metal2 s 220910 0 220966 800 6 la_data_out[29]
port 323 nsew signal output
rlabel metal2 s 128910 0 128966 800 6 la_data_out[2]
port 324 nsew signal output
rlabel metal2 s 224314 0 224370 800 6 la_data_out[30]
port 325 nsew signal output
rlabel metal2 s 227718 0 227774 800 6 la_data_out[31]
port 326 nsew signal output
rlabel metal2 s 231122 0 231178 800 6 la_data_out[32]
port 327 nsew signal output
rlabel metal2 s 234526 0 234582 800 6 la_data_out[33]
port 328 nsew signal output
rlabel metal2 s 237930 0 237986 800 6 la_data_out[34]
port 329 nsew signal output
rlabel metal2 s 241334 0 241390 800 6 la_data_out[35]
port 330 nsew signal output
rlabel metal2 s 244738 0 244794 800 6 la_data_out[36]
port 331 nsew signal output
rlabel metal2 s 248142 0 248198 800 6 la_data_out[37]
port 332 nsew signal output
rlabel metal2 s 251546 0 251602 800 6 la_data_out[38]
port 333 nsew signal output
rlabel metal2 s 254950 0 255006 800 6 la_data_out[39]
port 334 nsew signal output
rlabel metal2 s 132314 0 132370 800 6 la_data_out[3]
port 335 nsew signal output
rlabel metal2 s 258354 0 258410 800 6 la_data_out[40]
port 336 nsew signal output
rlabel metal2 s 261850 0 261906 800 6 la_data_out[41]
port 337 nsew signal output
rlabel metal2 s 265254 0 265310 800 6 la_data_out[42]
port 338 nsew signal output
rlabel metal2 s 268658 0 268714 800 6 la_data_out[43]
port 339 nsew signal output
rlabel metal2 s 272062 0 272118 800 6 la_data_out[44]
port 340 nsew signal output
rlabel metal2 s 275466 0 275522 800 6 la_data_out[45]
port 341 nsew signal output
rlabel metal2 s 278870 0 278926 800 6 la_data_out[46]
port 342 nsew signal output
rlabel metal2 s 282274 0 282330 800 6 la_data_out[47]
port 343 nsew signal output
rlabel metal2 s 285678 0 285734 800 6 la_data_out[48]
port 344 nsew signal output
rlabel metal2 s 289082 0 289138 800 6 la_data_out[49]
port 345 nsew signal output
rlabel metal2 s 135718 0 135774 800 6 la_data_out[4]
port 346 nsew signal output
rlabel metal2 s 292486 0 292542 800 6 la_data_out[50]
port 347 nsew signal output
rlabel metal2 s 295890 0 295946 800 6 la_data_out[51]
port 348 nsew signal output
rlabel metal2 s 299294 0 299350 800 6 la_data_out[52]
port 349 nsew signal output
rlabel metal2 s 302698 0 302754 800 6 la_data_out[53]
port 350 nsew signal output
rlabel metal2 s 306102 0 306158 800 6 la_data_out[54]
port 351 nsew signal output
rlabel metal2 s 309506 0 309562 800 6 la_data_out[55]
port 352 nsew signal output
rlabel metal2 s 312910 0 312966 800 6 la_data_out[56]
port 353 nsew signal output
rlabel metal2 s 316314 0 316370 800 6 la_data_out[57]
port 354 nsew signal output
rlabel metal2 s 319718 0 319774 800 6 la_data_out[58]
port 355 nsew signal output
rlabel metal2 s 323122 0 323178 800 6 la_data_out[59]
port 356 nsew signal output
rlabel metal2 s 139122 0 139178 800 6 la_data_out[5]
port 357 nsew signal output
rlabel metal2 s 326526 0 326582 800 6 la_data_out[60]
port 358 nsew signal output
rlabel metal2 s 329930 0 329986 800 6 la_data_out[61]
port 359 nsew signal output
rlabel metal2 s 333334 0 333390 800 6 la_data_out[62]
port 360 nsew signal output
rlabel metal2 s 336830 0 336886 800 6 la_data_out[63]
port 361 nsew signal output
rlabel metal2 s 340234 0 340290 800 6 la_data_out[64]
port 362 nsew signal output
rlabel metal2 s 343638 0 343694 800 6 la_data_out[65]
port 363 nsew signal output
rlabel metal2 s 347042 0 347098 800 6 la_data_out[66]
port 364 nsew signal output
rlabel metal2 s 350446 0 350502 800 6 la_data_out[67]
port 365 nsew signal output
rlabel metal2 s 353850 0 353906 800 6 la_data_out[68]
port 366 nsew signal output
rlabel metal2 s 357254 0 357310 800 6 la_data_out[69]
port 367 nsew signal output
rlabel metal2 s 142526 0 142582 800 6 la_data_out[6]
port 368 nsew signal output
rlabel metal2 s 360658 0 360714 800 6 la_data_out[70]
port 369 nsew signal output
rlabel metal2 s 364062 0 364118 800 6 la_data_out[71]
port 370 nsew signal output
rlabel metal2 s 367466 0 367522 800 6 la_data_out[72]
port 371 nsew signal output
rlabel metal2 s 370870 0 370926 800 6 la_data_out[73]
port 372 nsew signal output
rlabel metal2 s 374274 0 374330 800 6 la_data_out[74]
port 373 nsew signal output
rlabel metal2 s 377678 0 377734 800 6 la_data_out[75]
port 374 nsew signal output
rlabel metal2 s 381082 0 381138 800 6 la_data_out[76]
port 375 nsew signal output
rlabel metal2 s 384486 0 384542 800 6 la_data_out[77]
port 376 nsew signal output
rlabel metal2 s 387890 0 387946 800 6 la_data_out[78]
port 377 nsew signal output
rlabel metal2 s 391294 0 391350 800 6 la_data_out[79]
port 378 nsew signal output
rlabel metal2 s 145930 0 145986 800 6 la_data_out[7]
port 379 nsew signal output
rlabel metal2 s 394698 0 394754 800 6 la_data_out[80]
port 380 nsew signal output
rlabel metal2 s 398102 0 398158 800 6 la_data_out[81]
port 381 nsew signal output
rlabel metal2 s 401506 0 401562 800 6 la_data_out[82]
port 382 nsew signal output
rlabel metal2 s 404910 0 404966 800 6 la_data_out[83]
port 383 nsew signal output
rlabel metal2 s 408314 0 408370 800 6 la_data_out[84]
port 384 nsew signal output
rlabel metal2 s 411718 0 411774 800 6 la_data_out[85]
port 385 nsew signal output
rlabel metal2 s 415214 0 415270 800 6 la_data_out[86]
port 386 nsew signal output
rlabel metal2 s 418618 0 418674 800 6 la_data_out[87]
port 387 nsew signal output
rlabel metal2 s 422022 0 422078 800 6 la_data_out[88]
port 388 nsew signal output
rlabel metal2 s 425426 0 425482 800 6 la_data_out[89]
port 389 nsew signal output
rlabel metal2 s 149334 0 149390 800 6 la_data_out[8]
port 390 nsew signal output
rlabel metal2 s 428830 0 428886 800 6 la_data_out[90]
port 391 nsew signal output
rlabel metal2 s 432234 0 432290 800 6 la_data_out[91]
port 392 nsew signal output
rlabel metal2 s 435638 0 435694 800 6 la_data_out[92]
port 393 nsew signal output
rlabel metal2 s 439042 0 439098 800 6 la_data_out[93]
port 394 nsew signal output
rlabel metal2 s 442446 0 442502 800 6 la_data_out[94]
port 395 nsew signal output
rlabel metal2 s 445850 0 445906 800 6 la_data_out[95]
port 396 nsew signal output
rlabel metal2 s 449254 0 449310 800 6 la_data_out[96]
port 397 nsew signal output
rlabel metal2 s 452658 0 452714 800 6 la_data_out[97]
port 398 nsew signal output
rlabel metal2 s 456062 0 456118 800 6 la_data_out[98]
port 399 nsew signal output
rlabel metal2 s 459466 0 459522 800 6 la_data_out[99]
port 400 nsew signal output
rlabel metal2 s 152738 0 152794 800 6 la_data_out[9]
port 401 nsew signal output
rlabel metal2 s 123206 0 123262 800 6 la_oen[0]
port 402 nsew signal input
rlabel metal2 s 463974 0 464030 800 6 la_oen[100]
port 403 nsew signal input
rlabel metal2 s 467470 0 467526 800 6 la_oen[101]
port 404 nsew signal input
rlabel metal2 s 470874 0 470930 800 6 la_oen[102]
port 405 nsew signal input
rlabel metal2 s 474278 0 474334 800 6 la_oen[103]
port 406 nsew signal input
rlabel metal2 s 477682 0 477738 800 6 la_oen[104]
port 407 nsew signal input
rlabel metal2 s 481086 0 481142 800 6 la_oen[105]
port 408 nsew signal input
rlabel metal2 s 484490 0 484546 800 6 la_oen[106]
port 409 nsew signal input
rlabel metal2 s 487894 0 487950 800 6 la_oen[107]
port 410 nsew signal input
rlabel metal2 s 491298 0 491354 800 6 la_oen[108]
port 411 nsew signal input
rlabel metal2 s 494702 0 494758 800 6 la_oen[109]
port 412 nsew signal input
rlabel metal2 s 157338 0 157394 800 6 la_oen[10]
port 413 nsew signal input
rlabel metal2 s 498106 0 498162 800 6 la_oen[110]
port 414 nsew signal input
rlabel metal2 s 501510 0 501566 800 6 la_oen[111]
port 415 nsew signal input
rlabel metal2 s 504914 0 504970 800 6 la_oen[112]
port 416 nsew signal input
rlabel metal2 s 508318 0 508374 800 6 la_oen[113]
port 417 nsew signal input
rlabel metal2 s 511722 0 511778 800 6 la_oen[114]
port 418 nsew signal input
rlabel metal2 s 515126 0 515182 800 6 la_oen[115]
port 419 nsew signal input
rlabel metal2 s 518530 0 518586 800 6 la_oen[116]
port 420 nsew signal input
rlabel metal2 s 521934 0 521990 800 6 la_oen[117]
port 421 nsew signal input
rlabel metal2 s 525338 0 525394 800 6 la_oen[118]
port 422 nsew signal input
rlabel metal2 s 528742 0 528798 800 6 la_oen[119]
port 423 nsew signal input
rlabel metal2 s 160742 0 160798 800 6 la_oen[11]
port 424 nsew signal input
rlabel metal2 s 532146 0 532202 800 6 la_oen[120]
port 425 nsew signal input
rlabel metal2 s 535550 0 535606 800 6 la_oen[121]
port 426 nsew signal input
rlabel metal2 s 538954 0 539010 800 6 la_oen[122]
port 427 nsew signal input
rlabel metal2 s 542358 0 542414 800 6 la_oen[123]
port 428 nsew signal input
rlabel metal2 s 545854 0 545910 800 6 la_oen[124]
port 429 nsew signal input
rlabel metal2 s 549258 0 549314 800 6 la_oen[125]
port 430 nsew signal input
rlabel metal2 s 552662 0 552718 800 6 la_oen[126]
port 431 nsew signal input
rlabel metal2 s 556066 0 556122 800 6 la_oen[127]
port 432 nsew signal input
rlabel metal2 s 164146 0 164202 800 6 la_oen[12]
port 433 nsew signal input
rlabel metal2 s 167550 0 167606 800 6 la_oen[13]
port 434 nsew signal input
rlabel metal2 s 170954 0 171010 800 6 la_oen[14]
port 435 nsew signal input
rlabel metal2 s 174358 0 174414 800 6 la_oen[15]
port 436 nsew signal input
rlabel metal2 s 177762 0 177818 800 6 la_oen[16]
port 437 nsew signal input
rlabel metal2 s 181166 0 181222 800 6 la_oen[17]
port 438 nsew signal input
rlabel metal2 s 184570 0 184626 800 6 la_oen[18]
port 439 nsew signal input
rlabel metal2 s 187974 0 188030 800 6 la_oen[19]
port 440 nsew signal input
rlabel metal2 s 126610 0 126666 800 6 la_oen[1]
port 441 nsew signal input
rlabel metal2 s 191378 0 191434 800 6 la_oen[20]
port 442 nsew signal input
rlabel metal2 s 194782 0 194838 800 6 la_oen[21]
port 443 nsew signal input
rlabel metal2 s 198186 0 198242 800 6 la_oen[22]
port 444 nsew signal input
rlabel metal2 s 201590 0 201646 800 6 la_oen[23]
port 445 nsew signal input
rlabel metal2 s 204994 0 205050 800 6 la_oen[24]
port 446 nsew signal input
rlabel metal2 s 208398 0 208454 800 6 la_oen[25]
port 447 nsew signal input
rlabel metal2 s 211802 0 211858 800 6 la_oen[26]
port 448 nsew signal input
rlabel metal2 s 215206 0 215262 800 6 la_oen[27]
port 449 nsew signal input
rlabel metal2 s 218610 0 218666 800 6 la_oen[28]
port 450 nsew signal input
rlabel metal2 s 222014 0 222070 800 6 la_oen[29]
port 451 nsew signal input
rlabel metal2 s 130014 0 130070 800 6 la_oen[2]
port 452 nsew signal input
rlabel metal2 s 225418 0 225474 800 6 la_oen[30]
port 453 nsew signal input
rlabel metal2 s 228822 0 228878 800 6 la_oen[31]
port 454 nsew signal input
rlabel metal2 s 232226 0 232282 800 6 la_oen[32]
port 455 nsew signal input
rlabel metal2 s 235722 0 235778 800 6 la_oen[33]
port 456 nsew signal input
rlabel metal2 s 239126 0 239182 800 6 la_oen[34]
port 457 nsew signal input
rlabel metal2 s 242530 0 242586 800 6 la_oen[35]
port 458 nsew signal input
rlabel metal2 s 245934 0 245990 800 6 la_oen[36]
port 459 nsew signal input
rlabel metal2 s 249338 0 249394 800 6 la_oen[37]
port 460 nsew signal input
rlabel metal2 s 252742 0 252798 800 6 la_oen[38]
port 461 nsew signal input
rlabel metal2 s 256146 0 256202 800 6 la_oen[39]
port 462 nsew signal input
rlabel metal2 s 133418 0 133474 800 6 la_oen[3]
port 463 nsew signal input
rlabel metal2 s 259550 0 259606 800 6 la_oen[40]
port 464 nsew signal input
rlabel metal2 s 262954 0 263010 800 6 la_oen[41]
port 465 nsew signal input
rlabel metal2 s 266358 0 266414 800 6 la_oen[42]
port 466 nsew signal input
rlabel metal2 s 269762 0 269818 800 6 la_oen[43]
port 467 nsew signal input
rlabel metal2 s 273166 0 273222 800 6 la_oen[44]
port 468 nsew signal input
rlabel metal2 s 276570 0 276626 800 6 la_oen[45]
port 469 nsew signal input
rlabel metal2 s 279974 0 280030 800 6 la_oen[46]
port 470 nsew signal input
rlabel metal2 s 283378 0 283434 800 6 la_oen[47]
port 471 nsew signal input
rlabel metal2 s 286782 0 286838 800 6 la_oen[48]
port 472 nsew signal input
rlabel metal2 s 290186 0 290242 800 6 la_oen[49]
port 473 nsew signal input
rlabel metal2 s 136822 0 136878 800 6 la_oen[4]
port 474 nsew signal input
rlabel metal2 s 293590 0 293646 800 6 la_oen[50]
port 475 nsew signal input
rlabel metal2 s 296994 0 297050 800 6 la_oen[51]
port 476 nsew signal input
rlabel metal2 s 300398 0 300454 800 6 la_oen[52]
port 477 nsew signal input
rlabel metal2 s 303802 0 303858 800 6 la_oen[53]
port 478 nsew signal input
rlabel metal2 s 307206 0 307262 800 6 la_oen[54]
port 479 nsew signal input
rlabel metal2 s 310702 0 310758 800 6 la_oen[55]
port 480 nsew signal input
rlabel metal2 s 314106 0 314162 800 6 la_oen[56]
port 481 nsew signal input
rlabel metal2 s 317510 0 317566 800 6 la_oen[57]
port 482 nsew signal input
rlabel metal2 s 320914 0 320970 800 6 la_oen[58]
port 483 nsew signal input
rlabel metal2 s 324318 0 324374 800 6 la_oen[59]
port 484 nsew signal input
rlabel metal2 s 140226 0 140282 800 6 la_oen[5]
port 485 nsew signal input
rlabel metal2 s 327722 0 327778 800 6 la_oen[60]
port 486 nsew signal input
rlabel metal2 s 331126 0 331182 800 6 la_oen[61]
port 487 nsew signal input
rlabel metal2 s 334530 0 334586 800 6 la_oen[62]
port 488 nsew signal input
rlabel metal2 s 337934 0 337990 800 6 la_oen[63]
port 489 nsew signal input
rlabel metal2 s 341338 0 341394 800 6 la_oen[64]
port 490 nsew signal input
rlabel metal2 s 344742 0 344798 800 6 la_oen[65]
port 491 nsew signal input
rlabel metal2 s 348146 0 348202 800 6 la_oen[66]
port 492 nsew signal input
rlabel metal2 s 351550 0 351606 800 6 la_oen[67]
port 493 nsew signal input
rlabel metal2 s 354954 0 355010 800 6 la_oen[68]
port 494 nsew signal input
rlabel metal2 s 358358 0 358414 800 6 la_oen[69]
port 495 nsew signal input
rlabel metal2 s 143630 0 143686 800 6 la_oen[6]
port 496 nsew signal input
rlabel metal2 s 361762 0 361818 800 6 la_oen[70]
port 497 nsew signal input
rlabel metal2 s 365166 0 365222 800 6 la_oen[71]
port 498 nsew signal input
rlabel metal2 s 368570 0 368626 800 6 la_oen[72]
port 499 nsew signal input
rlabel metal2 s 371974 0 372030 800 6 la_oen[73]
port 500 nsew signal input
rlabel metal2 s 375378 0 375434 800 6 la_oen[74]
port 501 nsew signal input
rlabel metal2 s 378782 0 378838 800 6 la_oen[75]
port 502 nsew signal input
rlabel metal2 s 382186 0 382242 800 6 la_oen[76]
port 503 nsew signal input
rlabel metal2 s 385590 0 385646 800 6 la_oen[77]
port 504 nsew signal input
rlabel metal2 s 389086 0 389142 800 6 la_oen[78]
port 505 nsew signal input
rlabel metal2 s 392490 0 392546 800 6 la_oen[79]
port 506 nsew signal input
rlabel metal2 s 147034 0 147090 800 6 la_oen[7]
port 507 nsew signal input
rlabel metal2 s 395894 0 395950 800 6 la_oen[80]
port 508 nsew signal input
rlabel metal2 s 399298 0 399354 800 6 la_oen[81]
port 509 nsew signal input
rlabel metal2 s 402702 0 402758 800 6 la_oen[82]
port 510 nsew signal input
rlabel metal2 s 406106 0 406162 800 6 la_oen[83]
port 511 nsew signal input
rlabel metal2 s 409510 0 409566 800 6 la_oen[84]
port 512 nsew signal input
rlabel metal2 s 412914 0 412970 800 6 la_oen[85]
port 513 nsew signal input
rlabel metal2 s 416318 0 416374 800 6 la_oen[86]
port 514 nsew signal input
rlabel metal2 s 419722 0 419778 800 6 la_oen[87]
port 515 nsew signal input
rlabel metal2 s 423126 0 423182 800 6 la_oen[88]
port 516 nsew signal input
rlabel metal2 s 426530 0 426586 800 6 la_oen[89]
port 517 nsew signal input
rlabel metal2 s 150438 0 150494 800 6 la_oen[8]
port 518 nsew signal input
rlabel metal2 s 429934 0 429990 800 6 la_oen[90]
port 519 nsew signal input
rlabel metal2 s 433338 0 433394 800 6 la_oen[91]
port 520 nsew signal input
rlabel metal2 s 436742 0 436798 800 6 la_oen[92]
port 521 nsew signal input
rlabel metal2 s 440146 0 440202 800 6 la_oen[93]
port 522 nsew signal input
rlabel metal2 s 443550 0 443606 800 6 la_oen[94]
port 523 nsew signal input
rlabel metal2 s 446954 0 447010 800 6 la_oen[95]
port 524 nsew signal input
rlabel metal2 s 450358 0 450414 800 6 la_oen[96]
port 525 nsew signal input
rlabel metal2 s 453762 0 453818 800 6 la_oen[97]
port 526 nsew signal input
rlabel metal2 s 457166 0 457222 800 6 la_oen[98]
port 527 nsew signal input
rlabel metal2 s 460570 0 460626 800 6 la_oen[99]
port 528 nsew signal input
rlabel metal2 s 153842 0 153898 800 6 la_oen[9]
port 529 nsew signal input
rlabel metal2 s 557170 0 557226 800 6 user_clock2
port 530 nsew signal input
rlabel metal2 s 570 0 626 800 6 wb_clk_i
port 531 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wb_rst_i
port 532 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 wbs_ack_o
port 533 nsew signal output
rlabel metal2 s 7378 0 7434 800 6 wbs_adr_i[0]
port 534 nsew signal input
rlabel metal2 s 45926 0 45982 800 6 wbs_adr_i[10]
port 535 nsew signal input
rlabel metal2 s 49330 0 49386 800 6 wbs_adr_i[11]
port 536 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 wbs_adr_i[12]
port 537 nsew signal input
rlabel metal2 s 56230 0 56286 800 6 wbs_adr_i[13]
port 538 nsew signal input
rlabel metal2 s 59634 0 59690 800 6 wbs_adr_i[14]
port 539 nsew signal input
rlabel metal2 s 63038 0 63094 800 6 wbs_adr_i[15]
port 540 nsew signal input
rlabel metal2 s 66442 0 66498 800 6 wbs_adr_i[16]
port 541 nsew signal input
rlabel metal2 s 69846 0 69902 800 6 wbs_adr_i[17]
port 542 nsew signal input
rlabel metal2 s 73250 0 73306 800 6 wbs_adr_i[18]
port 543 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 wbs_adr_i[19]
port 544 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 wbs_adr_i[1]
port 545 nsew signal input
rlabel metal2 s 80058 0 80114 800 6 wbs_adr_i[20]
port 546 nsew signal input
rlabel metal2 s 83462 0 83518 800 6 wbs_adr_i[21]
port 547 nsew signal input
rlabel metal2 s 86866 0 86922 800 6 wbs_adr_i[22]
port 548 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 wbs_adr_i[23]
port 549 nsew signal input
rlabel metal2 s 93674 0 93730 800 6 wbs_adr_i[24]
port 550 nsew signal input
rlabel metal2 s 97078 0 97134 800 6 wbs_adr_i[25]
port 551 nsew signal input
rlabel metal2 s 100482 0 100538 800 6 wbs_adr_i[26]
port 552 nsew signal input
rlabel metal2 s 103886 0 103942 800 6 wbs_adr_i[27]
port 553 nsew signal input
rlabel metal2 s 107290 0 107346 800 6 wbs_adr_i[28]
port 554 nsew signal input
rlabel metal2 s 110694 0 110750 800 6 wbs_adr_i[29]
port 555 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 wbs_adr_i[2]
port 556 nsew signal input
rlabel metal2 s 114098 0 114154 800 6 wbs_adr_i[30]
port 557 nsew signal input
rlabel metal2 s 117502 0 117558 800 6 wbs_adr_i[31]
port 558 nsew signal input
rlabel metal2 s 20994 0 21050 800 6 wbs_adr_i[3]
port 559 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 wbs_adr_i[4]
port 560 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 wbs_adr_i[5]
port 561 nsew signal input
rlabel metal2 s 32310 0 32366 800 6 wbs_adr_i[6]
port 562 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 wbs_adr_i[7]
port 563 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 wbs_adr_i[8]
port 564 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 wbs_adr_i[9]
port 565 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 wbs_cyc_i
port 566 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_dat_i[0]
port 567 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 wbs_dat_i[10]
port 568 nsew signal input
rlabel metal2 s 50526 0 50582 800 6 wbs_dat_i[11]
port 569 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 wbs_dat_i[12]
port 570 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 wbs_dat_i[13]
port 571 nsew signal input
rlabel metal2 s 60738 0 60794 800 6 wbs_dat_i[14]
port 572 nsew signal input
rlabel metal2 s 64142 0 64198 800 6 wbs_dat_i[15]
port 573 nsew signal input
rlabel metal2 s 67546 0 67602 800 6 wbs_dat_i[16]
port 574 nsew signal input
rlabel metal2 s 70950 0 71006 800 6 wbs_dat_i[17]
port 575 nsew signal input
rlabel metal2 s 74354 0 74410 800 6 wbs_dat_i[18]
port 576 nsew signal input
rlabel metal2 s 77758 0 77814 800 6 wbs_dat_i[19]
port 577 nsew signal input
rlabel metal2 s 12990 0 13046 800 6 wbs_dat_i[1]
port 578 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 wbs_dat_i[20]
port 579 nsew signal input
rlabel metal2 s 84566 0 84622 800 6 wbs_dat_i[21]
port 580 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 wbs_dat_i[22]
port 581 nsew signal input
rlabel metal2 s 91374 0 91430 800 6 wbs_dat_i[23]
port 582 nsew signal input
rlabel metal2 s 94778 0 94834 800 6 wbs_dat_i[24]
port 583 nsew signal input
rlabel metal2 s 98182 0 98238 800 6 wbs_dat_i[25]
port 584 nsew signal input
rlabel metal2 s 101586 0 101642 800 6 wbs_dat_i[26]
port 585 nsew signal input
rlabel metal2 s 105082 0 105138 800 6 wbs_dat_i[27]
port 586 nsew signal input
rlabel metal2 s 108486 0 108542 800 6 wbs_dat_i[28]
port 587 nsew signal input
rlabel metal2 s 111890 0 111946 800 6 wbs_dat_i[29]
port 588 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 wbs_dat_i[2]
port 589 nsew signal input
rlabel metal2 s 115294 0 115350 800 6 wbs_dat_i[30]
port 590 nsew signal input
rlabel metal2 s 118698 0 118754 800 6 wbs_dat_i[31]
port 591 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 wbs_dat_i[3]
port 592 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 wbs_dat_i[4]
port 593 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 wbs_dat_i[5]
port 594 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 wbs_dat_i[6]
port 595 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 wbs_dat_i[7]
port 596 nsew signal input
rlabel metal2 s 40314 0 40370 800 6 wbs_dat_i[8]
port 597 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 wbs_dat_i[9]
port 598 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_dat_o[0]
port 599 nsew signal output
rlabel metal2 s 48226 0 48282 800 6 wbs_dat_o[10]
port 600 nsew signal output
rlabel metal2 s 51630 0 51686 800 6 wbs_dat_o[11]
port 601 nsew signal output
rlabel metal2 s 55034 0 55090 800 6 wbs_dat_o[12]
port 602 nsew signal output
rlabel metal2 s 58438 0 58494 800 6 wbs_dat_o[13]
port 603 nsew signal output
rlabel metal2 s 61842 0 61898 800 6 wbs_dat_o[14]
port 604 nsew signal output
rlabel metal2 s 65246 0 65302 800 6 wbs_dat_o[15]
port 605 nsew signal output
rlabel metal2 s 68650 0 68706 800 6 wbs_dat_o[16]
port 606 nsew signal output
rlabel metal2 s 72054 0 72110 800 6 wbs_dat_o[17]
port 607 nsew signal output
rlabel metal2 s 75458 0 75514 800 6 wbs_dat_o[18]
port 608 nsew signal output
rlabel metal2 s 78954 0 79010 800 6 wbs_dat_o[19]
port 609 nsew signal output
rlabel metal2 s 14186 0 14242 800 6 wbs_dat_o[1]
port 610 nsew signal output
rlabel metal2 s 82358 0 82414 800 6 wbs_dat_o[20]
port 611 nsew signal output
rlabel metal2 s 85762 0 85818 800 6 wbs_dat_o[21]
port 612 nsew signal output
rlabel metal2 s 89166 0 89222 800 6 wbs_dat_o[22]
port 613 nsew signal output
rlabel metal2 s 92570 0 92626 800 6 wbs_dat_o[23]
port 614 nsew signal output
rlabel metal2 s 95974 0 96030 800 6 wbs_dat_o[24]
port 615 nsew signal output
rlabel metal2 s 99378 0 99434 800 6 wbs_dat_o[25]
port 616 nsew signal output
rlabel metal2 s 102782 0 102838 800 6 wbs_dat_o[26]
port 617 nsew signal output
rlabel metal2 s 106186 0 106242 800 6 wbs_dat_o[27]
port 618 nsew signal output
rlabel metal2 s 109590 0 109646 800 6 wbs_dat_o[28]
port 619 nsew signal output
rlabel metal2 s 112994 0 113050 800 6 wbs_dat_o[29]
port 620 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 wbs_dat_o[2]
port 621 nsew signal output
rlabel metal2 s 116398 0 116454 800 6 wbs_dat_o[30]
port 622 nsew signal output
rlabel metal2 s 119802 0 119858 800 6 wbs_dat_o[31]
port 623 nsew signal output
rlabel metal2 s 23202 0 23258 800 6 wbs_dat_o[3]
port 624 nsew signal output
rlabel metal2 s 27802 0 27858 800 6 wbs_dat_o[4]
port 625 nsew signal output
rlabel metal2 s 31206 0 31262 800 6 wbs_dat_o[5]
port 626 nsew signal output
rlabel metal2 s 34610 0 34666 800 6 wbs_dat_o[6]
port 627 nsew signal output
rlabel metal2 s 38014 0 38070 800 6 wbs_dat_o[7]
port 628 nsew signal output
rlabel metal2 s 41418 0 41474 800 6 wbs_dat_o[8]
port 629 nsew signal output
rlabel metal2 s 44822 0 44878 800 6 wbs_dat_o[9]
port 630 nsew signal output
rlabel metal2 s 10782 0 10838 800 6 wbs_sel_i[0]
port 631 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 wbs_sel_i[1]
port 632 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 wbs_sel_i[2]
port 633 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 wbs_sel_i[3]
port 634 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 wbs_stb_i
port 635 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wbs_we_i
port 636 nsew signal input
rlabel metal4 s 557168 2128 557488 685488 6 VPWR
port 637 nsew power bidirectional
rlabel metal4 s 526448 2128 526768 685488 6 VPWR
port 638 nsew power bidirectional
rlabel metal4 s 495728 2128 496048 685488 6 VPWR
port 639 nsew power bidirectional
rlabel metal4 s 465008 2128 465328 685488 6 VPWR
port 640 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 685488 6 VPWR
port 641 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 685488 6 VPWR
port 642 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 685488 6 VPWR
port 643 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 685488 6 VPWR
port 644 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 685488 6 VPWR
port 645 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 685488 6 VPWR
port 646 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 685488 6 VPWR
port 647 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 685488 6 VPWR
port 648 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 685488 6 VPWR
port 649 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 685488 6 VPWR
port 650 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 685488 6 VPWR
port 651 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 685488 6 VPWR
port 652 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 685488 6 VPWR
port 653 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 685488 6 VPWR
port 654 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 685488 6 VPWR
port 655 nsew power bidirectional
rlabel metal4 s 541808 2128 542128 685488 6 VGND
port 656 nsew ground bidirectional
rlabel metal4 s 511088 2128 511408 685488 6 VGND
port 657 nsew ground bidirectional
rlabel metal4 s 480368 2128 480688 685488 6 VGND
port 658 nsew ground bidirectional
rlabel metal4 s 449648 2128 449968 685488 6 VGND
port 659 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 685488 6 VGND
port 660 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 685488 6 VGND
port 661 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 685488 6 VGND
port 662 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 685488 6 VGND
port 663 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 685488 6 VGND
port 664 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 685488 6 VGND
port 665 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 685488 6 VGND
port 666 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 685488 6 VGND
port 667 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 685488 6 VGND
port 668 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 685488 6 VGND
port 669 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 685488 6 VGND
port 670 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 685488 6 VGND
port 671 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 685488 6 VGND
port 672 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 685488 6 VGND
port 673 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 568000 688000
string LEFview TRUE
<< end >>

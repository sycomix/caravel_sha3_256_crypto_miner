magic
tech sky130A
magscale 1 2
timestamp 1608118574
<< obsli1 >>
rect 1104 2159 562856 681649
<< obsm1 >>
rect 566 1096 562856 681680
<< metal2 >>
rect 2318 683200 2374 684000
rect 6918 683200 6974 684000
rect 11518 683200 11574 684000
rect 16118 683200 16174 684000
rect 20718 683200 20774 684000
rect 25410 683200 25466 684000
rect 30010 683200 30066 684000
rect 34610 683200 34666 684000
rect 39210 683200 39266 684000
rect 43902 683200 43958 684000
rect 48502 683200 48558 684000
rect 53102 683200 53158 684000
rect 57702 683200 57758 684000
rect 62394 683200 62450 684000
rect 66994 683200 67050 684000
rect 71594 683200 71650 684000
rect 76194 683200 76250 684000
rect 80886 683200 80942 684000
rect 85486 683200 85542 684000
rect 90086 683200 90142 684000
rect 94686 683200 94742 684000
rect 99378 683200 99434 684000
rect 103978 683200 104034 684000
rect 108578 683200 108634 684000
rect 113178 683200 113234 684000
rect 117870 683200 117926 684000
rect 122470 683200 122526 684000
rect 127070 683200 127126 684000
rect 131670 683200 131726 684000
rect 136362 683200 136418 684000
rect 140962 683200 141018 684000
rect 145562 683200 145618 684000
rect 150162 683200 150218 684000
rect 154854 683200 154910 684000
rect 159454 683200 159510 684000
rect 164054 683200 164110 684000
rect 168654 683200 168710 684000
rect 173346 683200 173402 684000
rect 177946 683200 178002 684000
rect 182546 683200 182602 684000
rect 187146 683200 187202 684000
rect 191838 683200 191894 684000
rect 196438 683200 196494 684000
rect 201038 683200 201094 684000
rect 205638 683200 205694 684000
rect 210330 683200 210386 684000
rect 214930 683200 214986 684000
rect 219530 683200 219586 684000
rect 224130 683200 224186 684000
rect 228822 683200 228878 684000
rect 233422 683200 233478 684000
rect 238022 683200 238078 684000
rect 242622 683200 242678 684000
rect 247314 683200 247370 684000
rect 251914 683200 251970 684000
rect 256514 683200 256570 684000
rect 261114 683200 261170 684000
rect 265806 683200 265862 684000
rect 270406 683200 270462 684000
rect 275006 683200 275062 684000
rect 279606 683200 279662 684000
rect 284298 683200 284354 684000
rect 288898 683200 288954 684000
rect 293498 683200 293554 684000
rect 298098 683200 298154 684000
rect 302698 683200 302754 684000
rect 307390 683200 307446 684000
rect 311990 683200 312046 684000
rect 316590 683200 316646 684000
rect 321190 683200 321246 684000
rect 325882 683200 325938 684000
rect 330482 683200 330538 684000
rect 335082 683200 335138 684000
rect 339682 683200 339738 684000
rect 344374 683200 344430 684000
rect 348974 683200 349030 684000
rect 353574 683200 353630 684000
rect 358174 683200 358230 684000
rect 362866 683200 362922 684000
rect 367466 683200 367522 684000
rect 372066 683200 372122 684000
rect 376666 683200 376722 684000
rect 381358 683200 381414 684000
rect 385958 683200 386014 684000
rect 390558 683200 390614 684000
rect 395158 683200 395214 684000
rect 399850 683200 399906 684000
rect 404450 683200 404506 684000
rect 409050 683200 409106 684000
rect 413650 683200 413706 684000
rect 418342 683200 418398 684000
rect 422942 683200 422998 684000
rect 427542 683200 427598 684000
rect 432142 683200 432198 684000
rect 436834 683200 436890 684000
rect 441434 683200 441490 684000
rect 446034 683200 446090 684000
rect 450634 683200 450690 684000
rect 455326 683200 455382 684000
rect 459926 683200 459982 684000
rect 464526 683200 464582 684000
rect 469126 683200 469182 684000
rect 473818 683200 473874 684000
rect 478418 683200 478474 684000
rect 483018 683200 483074 684000
rect 487618 683200 487674 684000
rect 492310 683200 492366 684000
rect 496910 683200 496966 684000
rect 501510 683200 501566 684000
rect 506110 683200 506166 684000
rect 510802 683200 510858 684000
rect 515402 683200 515458 684000
rect 520002 683200 520058 684000
rect 524602 683200 524658 684000
rect 529294 683200 529350 684000
rect 533894 683200 533950 684000
rect 538494 683200 538550 684000
rect 543094 683200 543150 684000
rect 547786 683200 547842 684000
rect 552386 683200 552442 684000
rect 556986 683200 557042 684000
rect 561586 683200 561642 684000
rect 570 0 626 800
rect 1674 0 1730 800
rect 2778 0 2834 800
rect 3974 0 4030 800
rect 5078 0 5134 800
rect 6182 0 6238 800
rect 7378 0 7434 800
rect 8482 0 8538 800
rect 9586 0 9642 800
rect 10782 0 10838 800
rect 11886 0 11942 800
rect 12990 0 13046 800
rect 14186 0 14242 800
rect 15290 0 15346 800
rect 16486 0 16542 800
rect 17590 0 17646 800
rect 18694 0 18750 800
rect 19890 0 19946 800
rect 20994 0 21050 800
rect 22098 0 22154 800
rect 23294 0 23350 800
rect 24398 0 24454 800
rect 25502 0 25558 800
rect 26698 0 26754 800
rect 27802 0 27858 800
rect 28906 0 28962 800
rect 30102 0 30158 800
rect 31206 0 31262 800
rect 32402 0 32458 800
rect 33506 0 33562 800
rect 34610 0 34666 800
rect 35806 0 35862 800
rect 36910 0 36966 800
rect 38014 0 38070 800
rect 39210 0 39266 800
rect 40314 0 40370 800
rect 41418 0 41474 800
rect 42614 0 42670 800
rect 43718 0 43774 800
rect 44822 0 44878 800
rect 46018 0 46074 800
rect 47122 0 47178 800
rect 48318 0 48374 800
rect 49422 0 49478 800
rect 50526 0 50582 800
rect 51722 0 51778 800
rect 52826 0 52882 800
rect 53930 0 53986 800
rect 55126 0 55182 800
rect 56230 0 56286 800
rect 57334 0 57390 800
rect 58530 0 58586 800
rect 59634 0 59690 800
rect 60830 0 60886 800
rect 61934 0 61990 800
rect 63038 0 63094 800
rect 64234 0 64290 800
rect 65338 0 65394 800
rect 66442 0 66498 800
rect 67638 0 67694 800
rect 68742 0 68798 800
rect 69846 0 69902 800
rect 71042 0 71098 800
rect 72146 0 72202 800
rect 73250 0 73306 800
rect 74446 0 74502 800
rect 75550 0 75606 800
rect 76746 0 76802 800
rect 77850 0 77906 800
rect 78954 0 79010 800
rect 80150 0 80206 800
rect 81254 0 81310 800
rect 82358 0 82414 800
rect 83554 0 83610 800
rect 84658 0 84714 800
rect 85762 0 85818 800
rect 86958 0 87014 800
rect 88062 0 88118 800
rect 89166 0 89222 800
rect 90362 0 90418 800
rect 91466 0 91522 800
rect 92662 0 92718 800
rect 93766 0 93822 800
rect 94870 0 94926 800
rect 96066 0 96122 800
rect 97170 0 97226 800
rect 98274 0 98330 800
rect 99470 0 99526 800
rect 100574 0 100630 800
rect 101678 0 101734 800
rect 102874 0 102930 800
rect 103978 0 104034 800
rect 105174 0 105230 800
rect 106278 0 106334 800
rect 107382 0 107438 800
rect 108578 0 108634 800
rect 109682 0 109738 800
rect 110786 0 110842 800
rect 111982 0 112038 800
rect 113086 0 113142 800
rect 114190 0 114246 800
rect 115386 0 115442 800
rect 116490 0 116546 800
rect 117594 0 117650 800
rect 118790 0 118846 800
rect 119894 0 119950 800
rect 121090 0 121146 800
rect 122194 0 122250 800
rect 123298 0 123354 800
rect 124494 0 124550 800
rect 125598 0 125654 800
rect 126702 0 126758 800
rect 127898 0 127954 800
rect 129002 0 129058 800
rect 130106 0 130162 800
rect 131302 0 131358 800
rect 132406 0 132462 800
rect 133510 0 133566 800
rect 134706 0 134762 800
rect 135810 0 135866 800
rect 137006 0 137062 800
rect 138110 0 138166 800
rect 139214 0 139270 800
rect 140410 0 140466 800
rect 141514 0 141570 800
rect 142618 0 142674 800
rect 143814 0 143870 800
rect 144918 0 144974 800
rect 146022 0 146078 800
rect 147218 0 147274 800
rect 148322 0 148378 800
rect 149518 0 149574 800
rect 150622 0 150678 800
rect 151726 0 151782 800
rect 152922 0 152978 800
rect 154026 0 154082 800
rect 155130 0 155186 800
rect 156326 0 156382 800
rect 157430 0 157486 800
rect 158534 0 158590 800
rect 159730 0 159786 800
rect 160834 0 160890 800
rect 161938 0 161994 800
rect 163134 0 163190 800
rect 164238 0 164294 800
rect 165434 0 165490 800
rect 166538 0 166594 800
rect 167642 0 167698 800
rect 168838 0 168894 800
rect 169942 0 169998 800
rect 171046 0 171102 800
rect 172242 0 172298 800
rect 173346 0 173402 800
rect 174450 0 174506 800
rect 175646 0 175702 800
rect 176750 0 176806 800
rect 177854 0 177910 800
rect 179050 0 179106 800
rect 180154 0 180210 800
rect 181350 0 181406 800
rect 182454 0 182510 800
rect 183558 0 183614 800
rect 184754 0 184810 800
rect 185858 0 185914 800
rect 186962 0 187018 800
rect 188158 0 188214 800
rect 189262 0 189318 800
rect 190366 0 190422 800
rect 191562 0 191618 800
rect 192666 0 192722 800
rect 193862 0 193918 800
rect 194966 0 195022 800
rect 196070 0 196126 800
rect 197266 0 197322 800
rect 198370 0 198426 800
rect 199474 0 199530 800
rect 200670 0 200726 800
rect 201774 0 201830 800
rect 202878 0 202934 800
rect 204074 0 204130 800
rect 205178 0 205234 800
rect 206282 0 206338 800
rect 207478 0 207534 800
rect 208582 0 208638 800
rect 209778 0 209834 800
rect 210882 0 210938 800
rect 211986 0 212042 800
rect 213182 0 213238 800
rect 214286 0 214342 800
rect 215390 0 215446 800
rect 216586 0 216642 800
rect 217690 0 217746 800
rect 218794 0 218850 800
rect 219990 0 220046 800
rect 221094 0 221150 800
rect 222198 0 222254 800
rect 223394 0 223450 800
rect 224498 0 224554 800
rect 225694 0 225750 800
rect 226798 0 226854 800
rect 227902 0 227958 800
rect 229098 0 229154 800
rect 230202 0 230258 800
rect 231306 0 231362 800
rect 232502 0 232558 800
rect 233606 0 233662 800
rect 234710 0 234766 800
rect 235906 0 235962 800
rect 237010 0 237066 800
rect 238206 0 238262 800
rect 239310 0 239366 800
rect 240414 0 240470 800
rect 241610 0 241666 800
rect 242714 0 242770 800
rect 243818 0 243874 800
rect 245014 0 245070 800
rect 246118 0 246174 800
rect 247222 0 247278 800
rect 248418 0 248474 800
rect 249522 0 249578 800
rect 250626 0 250682 800
rect 251822 0 251878 800
rect 252926 0 252982 800
rect 254122 0 254178 800
rect 255226 0 255282 800
rect 256330 0 256386 800
rect 257526 0 257582 800
rect 258630 0 258686 800
rect 259734 0 259790 800
rect 260930 0 260986 800
rect 262034 0 262090 800
rect 263138 0 263194 800
rect 264334 0 264390 800
rect 265438 0 265494 800
rect 266542 0 266598 800
rect 267738 0 267794 800
rect 268842 0 268898 800
rect 270038 0 270094 800
rect 271142 0 271198 800
rect 272246 0 272302 800
rect 273442 0 273498 800
rect 274546 0 274602 800
rect 275650 0 275706 800
rect 276846 0 276902 800
rect 277950 0 278006 800
rect 279054 0 279110 800
rect 280250 0 280306 800
rect 281354 0 281410 800
rect 282550 0 282606 800
rect 283654 0 283710 800
rect 284758 0 284814 800
rect 285954 0 286010 800
rect 287058 0 287114 800
rect 288162 0 288218 800
rect 289358 0 289414 800
rect 290462 0 290518 800
rect 291566 0 291622 800
rect 292762 0 292818 800
rect 293866 0 293922 800
rect 294970 0 295026 800
rect 296166 0 296222 800
rect 297270 0 297326 800
rect 298466 0 298522 800
rect 299570 0 299626 800
rect 300674 0 300730 800
rect 301870 0 301926 800
rect 302974 0 303030 800
rect 304078 0 304134 800
rect 305274 0 305330 800
rect 306378 0 306434 800
rect 307482 0 307538 800
rect 308678 0 308734 800
rect 309782 0 309838 800
rect 310886 0 310942 800
rect 312082 0 312138 800
rect 313186 0 313242 800
rect 314382 0 314438 800
rect 315486 0 315542 800
rect 316590 0 316646 800
rect 317786 0 317842 800
rect 318890 0 318946 800
rect 319994 0 320050 800
rect 321190 0 321246 800
rect 322294 0 322350 800
rect 323398 0 323454 800
rect 324594 0 324650 800
rect 325698 0 325754 800
rect 326802 0 326858 800
rect 327998 0 328054 800
rect 329102 0 329158 800
rect 330298 0 330354 800
rect 331402 0 331458 800
rect 332506 0 332562 800
rect 333702 0 333758 800
rect 334806 0 334862 800
rect 335910 0 335966 800
rect 337106 0 337162 800
rect 338210 0 338266 800
rect 339314 0 339370 800
rect 340510 0 340566 800
rect 341614 0 341670 800
rect 342810 0 342866 800
rect 343914 0 343970 800
rect 345018 0 345074 800
rect 346214 0 346270 800
rect 347318 0 347374 800
rect 348422 0 348478 800
rect 349618 0 349674 800
rect 350722 0 350778 800
rect 351826 0 351882 800
rect 353022 0 353078 800
rect 354126 0 354182 800
rect 355230 0 355286 800
rect 356426 0 356482 800
rect 357530 0 357586 800
rect 358726 0 358782 800
rect 359830 0 359886 800
rect 360934 0 360990 800
rect 362130 0 362186 800
rect 363234 0 363290 800
rect 364338 0 364394 800
rect 365534 0 365590 800
rect 366638 0 366694 800
rect 367742 0 367798 800
rect 368938 0 368994 800
rect 370042 0 370098 800
rect 371146 0 371202 800
rect 372342 0 372398 800
rect 373446 0 373502 800
rect 374642 0 374698 800
rect 375746 0 375802 800
rect 376850 0 376906 800
rect 378046 0 378102 800
rect 379150 0 379206 800
rect 380254 0 380310 800
rect 381450 0 381506 800
rect 382554 0 382610 800
rect 383658 0 383714 800
rect 384854 0 384910 800
rect 385958 0 386014 800
rect 387154 0 387210 800
rect 388258 0 388314 800
rect 389362 0 389418 800
rect 390558 0 390614 800
rect 391662 0 391718 800
rect 392766 0 392822 800
rect 393962 0 394018 800
rect 395066 0 395122 800
rect 396170 0 396226 800
rect 397366 0 397422 800
rect 398470 0 398526 800
rect 399574 0 399630 800
rect 400770 0 400826 800
rect 401874 0 401930 800
rect 403070 0 403126 800
rect 404174 0 404230 800
rect 405278 0 405334 800
rect 406474 0 406530 800
rect 407578 0 407634 800
rect 408682 0 408738 800
rect 409878 0 409934 800
rect 410982 0 411038 800
rect 412086 0 412142 800
rect 413282 0 413338 800
rect 414386 0 414442 800
rect 415490 0 415546 800
rect 416686 0 416742 800
rect 417790 0 417846 800
rect 418986 0 419042 800
rect 420090 0 420146 800
rect 421194 0 421250 800
rect 422390 0 422446 800
rect 423494 0 423550 800
rect 424598 0 424654 800
rect 425794 0 425850 800
rect 426898 0 426954 800
rect 428002 0 428058 800
rect 429198 0 429254 800
rect 430302 0 430358 800
rect 431498 0 431554 800
rect 432602 0 432658 800
rect 433706 0 433762 800
rect 434902 0 434958 800
rect 436006 0 436062 800
rect 437110 0 437166 800
rect 438306 0 438362 800
rect 439410 0 439466 800
rect 440514 0 440570 800
rect 441710 0 441766 800
rect 442814 0 442870 800
rect 443918 0 443974 800
rect 445114 0 445170 800
rect 446218 0 446274 800
rect 447414 0 447470 800
rect 448518 0 448574 800
rect 449622 0 449678 800
rect 450818 0 450874 800
rect 451922 0 451978 800
rect 453026 0 453082 800
rect 454222 0 454278 800
rect 455326 0 455382 800
rect 456430 0 456486 800
rect 457626 0 457682 800
rect 458730 0 458786 800
rect 459834 0 459890 800
rect 461030 0 461086 800
rect 462134 0 462190 800
rect 463330 0 463386 800
rect 464434 0 464490 800
rect 465538 0 465594 800
rect 466734 0 466790 800
rect 467838 0 467894 800
rect 468942 0 468998 800
rect 470138 0 470194 800
rect 471242 0 471298 800
rect 472346 0 472402 800
rect 473542 0 473598 800
rect 474646 0 474702 800
rect 475842 0 475898 800
rect 476946 0 477002 800
rect 478050 0 478106 800
rect 479246 0 479302 800
rect 480350 0 480406 800
rect 481454 0 481510 800
rect 482650 0 482706 800
rect 483754 0 483810 800
rect 484858 0 484914 800
rect 486054 0 486110 800
rect 487158 0 487214 800
rect 488262 0 488318 800
rect 489458 0 489514 800
rect 490562 0 490618 800
rect 491758 0 491814 800
rect 492862 0 492918 800
rect 493966 0 494022 800
rect 495162 0 495218 800
rect 496266 0 496322 800
rect 497370 0 497426 800
rect 498566 0 498622 800
rect 499670 0 499726 800
rect 500774 0 500830 800
rect 501970 0 502026 800
rect 503074 0 503130 800
rect 504178 0 504234 800
rect 505374 0 505430 800
rect 506478 0 506534 800
rect 507674 0 507730 800
rect 508778 0 508834 800
rect 509882 0 509938 800
rect 511078 0 511134 800
rect 512182 0 512238 800
rect 513286 0 513342 800
rect 514482 0 514538 800
rect 515586 0 515642 800
rect 516690 0 516746 800
rect 517886 0 517942 800
rect 518990 0 519046 800
rect 520186 0 520242 800
rect 521290 0 521346 800
rect 522394 0 522450 800
rect 523590 0 523646 800
rect 524694 0 524750 800
rect 525798 0 525854 800
rect 526994 0 527050 800
rect 528098 0 528154 800
rect 529202 0 529258 800
rect 530398 0 530454 800
rect 531502 0 531558 800
rect 532606 0 532662 800
rect 533802 0 533858 800
rect 534906 0 534962 800
rect 536102 0 536158 800
rect 537206 0 537262 800
rect 538310 0 538366 800
rect 539506 0 539562 800
rect 540610 0 540666 800
rect 541714 0 541770 800
rect 542910 0 542966 800
rect 544014 0 544070 800
rect 545118 0 545174 800
rect 546314 0 546370 800
rect 547418 0 547474 800
rect 548522 0 548578 800
rect 549718 0 549774 800
rect 550822 0 550878 800
rect 552018 0 552074 800
rect 553122 0 553178 800
rect 554226 0 554282 800
rect 555422 0 555478 800
rect 556526 0 556582 800
rect 557630 0 557686 800
rect 558826 0 558882 800
rect 559930 0 559986 800
rect 561034 0 561090 800
rect 562230 0 562286 800
rect 563334 0 563390 800
<< obsm2 >>
rect 572 683144 2262 683200
rect 2430 683144 6862 683200
rect 7030 683144 11462 683200
rect 11630 683144 16062 683200
rect 16230 683144 20662 683200
rect 20830 683144 25354 683200
rect 25522 683144 29954 683200
rect 30122 683144 34554 683200
rect 34722 683144 39154 683200
rect 39322 683144 43846 683200
rect 44014 683144 48446 683200
rect 48614 683144 53046 683200
rect 53214 683144 57646 683200
rect 57814 683144 62338 683200
rect 62506 683144 66938 683200
rect 67106 683144 71538 683200
rect 71706 683144 76138 683200
rect 76306 683144 80830 683200
rect 80998 683144 85430 683200
rect 85598 683144 90030 683200
rect 90198 683144 94630 683200
rect 94798 683144 99322 683200
rect 99490 683144 103922 683200
rect 104090 683144 108522 683200
rect 108690 683144 113122 683200
rect 113290 683144 117814 683200
rect 117982 683144 122414 683200
rect 122582 683144 127014 683200
rect 127182 683144 131614 683200
rect 131782 683144 136306 683200
rect 136474 683144 140906 683200
rect 141074 683144 145506 683200
rect 145674 683144 150106 683200
rect 150274 683144 154798 683200
rect 154966 683144 159398 683200
rect 159566 683144 163998 683200
rect 164166 683144 168598 683200
rect 168766 683144 173290 683200
rect 173458 683144 177890 683200
rect 178058 683144 182490 683200
rect 182658 683144 187090 683200
rect 187258 683144 191782 683200
rect 191950 683144 196382 683200
rect 196550 683144 200982 683200
rect 201150 683144 205582 683200
rect 205750 683144 210274 683200
rect 210442 683144 214874 683200
rect 215042 683144 219474 683200
rect 219642 683144 224074 683200
rect 224242 683144 228766 683200
rect 228934 683144 233366 683200
rect 233534 683144 237966 683200
rect 238134 683144 242566 683200
rect 242734 683144 247258 683200
rect 247426 683144 251858 683200
rect 252026 683144 256458 683200
rect 256626 683144 261058 683200
rect 261226 683144 265750 683200
rect 265918 683144 270350 683200
rect 270518 683144 274950 683200
rect 275118 683144 279550 683200
rect 279718 683144 284242 683200
rect 284410 683144 288842 683200
rect 289010 683144 293442 683200
rect 293610 683144 298042 683200
rect 298210 683144 302642 683200
rect 302810 683144 307334 683200
rect 307502 683144 311934 683200
rect 312102 683144 316534 683200
rect 316702 683144 321134 683200
rect 321302 683144 325826 683200
rect 325994 683144 330426 683200
rect 330594 683144 335026 683200
rect 335194 683144 339626 683200
rect 339794 683144 344318 683200
rect 344486 683144 348918 683200
rect 349086 683144 353518 683200
rect 353686 683144 358118 683200
rect 358286 683144 362810 683200
rect 362978 683144 367410 683200
rect 367578 683144 372010 683200
rect 372178 683144 376610 683200
rect 376778 683144 381302 683200
rect 381470 683144 385902 683200
rect 386070 683144 390502 683200
rect 390670 683144 395102 683200
rect 395270 683144 399794 683200
rect 399962 683144 404394 683200
rect 404562 683144 408994 683200
rect 409162 683144 413594 683200
rect 413762 683144 418286 683200
rect 418454 683144 422886 683200
rect 423054 683144 427486 683200
rect 427654 683144 432086 683200
rect 432254 683144 436778 683200
rect 436946 683144 441378 683200
rect 441546 683144 445978 683200
rect 446146 683144 450578 683200
rect 450746 683144 455270 683200
rect 455438 683144 459870 683200
rect 460038 683144 464470 683200
rect 464638 683144 469070 683200
rect 469238 683144 473762 683200
rect 473930 683144 478362 683200
rect 478530 683144 482962 683200
rect 483130 683144 487562 683200
rect 487730 683144 492254 683200
rect 492422 683144 496854 683200
rect 497022 683144 501454 683200
rect 501622 683144 506054 683200
rect 506222 683144 510746 683200
rect 510914 683144 515346 683200
rect 515514 683144 519946 683200
rect 520114 683144 524546 683200
rect 524714 683144 529238 683200
rect 529406 683144 533838 683200
rect 534006 683144 538438 683200
rect 538606 683144 543038 683200
rect 543206 683144 547730 683200
rect 547898 683144 552330 683200
rect 552498 683144 556930 683200
rect 557098 683144 557672 683200
rect 572 856 557672 683144
rect 682 800 1618 856
rect 1786 800 2722 856
rect 2890 800 3918 856
rect 4086 800 5022 856
rect 5190 800 6126 856
rect 6294 800 7322 856
rect 7490 800 8426 856
rect 8594 800 9530 856
rect 9698 800 10726 856
rect 10894 800 11830 856
rect 11998 800 12934 856
rect 13102 800 14130 856
rect 14298 800 15234 856
rect 15402 800 16430 856
rect 16598 800 17534 856
rect 17702 800 18638 856
rect 18806 800 19834 856
rect 20002 800 20938 856
rect 21106 800 22042 856
rect 22210 800 23238 856
rect 23406 800 24342 856
rect 24510 800 25446 856
rect 25614 800 26642 856
rect 26810 800 27746 856
rect 27914 800 28850 856
rect 29018 800 30046 856
rect 30214 800 31150 856
rect 31318 800 32346 856
rect 32514 800 33450 856
rect 33618 800 34554 856
rect 34722 800 35750 856
rect 35918 800 36854 856
rect 37022 800 37958 856
rect 38126 800 39154 856
rect 39322 800 40258 856
rect 40426 800 41362 856
rect 41530 800 42558 856
rect 42726 800 43662 856
rect 43830 800 44766 856
rect 44934 800 45962 856
rect 46130 800 47066 856
rect 47234 800 48262 856
rect 48430 800 49366 856
rect 49534 800 50470 856
rect 50638 800 51666 856
rect 51834 800 52770 856
rect 52938 800 53874 856
rect 54042 800 55070 856
rect 55238 800 56174 856
rect 56342 800 57278 856
rect 57446 800 58474 856
rect 58642 800 59578 856
rect 59746 800 60774 856
rect 60942 800 61878 856
rect 62046 800 62982 856
rect 63150 800 64178 856
rect 64346 800 65282 856
rect 65450 800 66386 856
rect 66554 800 67582 856
rect 67750 800 68686 856
rect 68854 800 69790 856
rect 69958 800 70986 856
rect 71154 800 72090 856
rect 72258 800 73194 856
rect 73362 800 74390 856
rect 74558 800 75494 856
rect 75662 800 76690 856
rect 76858 800 77794 856
rect 77962 800 78898 856
rect 79066 800 80094 856
rect 80262 800 81198 856
rect 81366 800 82302 856
rect 82470 800 83498 856
rect 83666 800 84602 856
rect 84770 800 85706 856
rect 85874 800 86902 856
rect 87070 800 88006 856
rect 88174 800 89110 856
rect 89278 800 90306 856
rect 90474 800 91410 856
rect 91578 800 92606 856
rect 92774 800 93710 856
rect 93878 800 94814 856
rect 94982 800 96010 856
rect 96178 800 97114 856
rect 97282 800 98218 856
rect 98386 800 99414 856
rect 99582 800 100518 856
rect 100686 800 101622 856
rect 101790 800 102818 856
rect 102986 800 103922 856
rect 104090 800 105118 856
rect 105286 800 106222 856
rect 106390 800 107326 856
rect 107494 800 108522 856
rect 108690 800 109626 856
rect 109794 800 110730 856
rect 110898 800 111926 856
rect 112094 800 113030 856
rect 113198 800 114134 856
rect 114302 800 115330 856
rect 115498 800 116434 856
rect 116602 800 117538 856
rect 117706 800 118734 856
rect 118902 800 119838 856
rect 120006 800 121034 856
rect 121202 800 122138 856
rect 122306 800 123242 856
rect 123410 800 124438 856
rect 124606 800 125542 856
rect 125710 800 126646 856
rect 126814 800 127842 856
rect 128010 800 128946 856
rect 129114 800 130050 856
rect 130218 800 131246 856
rect 131414 800 132350 856
rect 132518 800 133454 856
rect 133622 800 134650 856
rect 134818 800 135754 856
rect 135922 800 136950 856
rect 137118 800 138054 856
rect 138222 800 139158 856
rect 139326 800 140354 856
rect 140522 800 141458 856
rect 141626 800 142562 856
rect 142730 800 143758 856
rect 143926 800 144862 856
rect 145030 800 145966 856
rect 146134 800 147162 856
rect 147330 800 148266 856
rect 148434 800 149462 856
rect 149630 800 150566 856
rect 150734 800 151670 856
rect 151838 800 152866 856
rect 153034 800 153970 856
rect 154138 800 155074 856
rect 155242 800 156270 856
rect 156438 800 157374 856
rect 157542 800 158478 856
rect 158646 800 159674 856
rect 159842 800 160778 856
rect 160946 800 161882 856
rect 162050 800 163078 856
rect 163246 800 164182 856
rect 164350 800 165378 856
rect 165546 800 166482 856
rect 166650 800 167586 856
rect 167754 800 168782 856
rect 168950 800 169886 856
rect 170054 800 170990 856
rect 171158 800 172186 856
rect 172354 800 173290 856
rect 173458 800 174394 856
rect 174562 800 175590 856
rect 175758 800 176694 856
rect 176862 800 177798 856
rect 177966 800 178994 856
rect 179162 800 180098 856
rect 180266 800 181294 856
rect 181462 800 182398 856
rect 182566 800 183502 856
rect 183670 800 184698 856
rect 184866 800 185802 856
rect 185970 800 186906 856
rect 187074 800 188102 856
rect 188270 800 189206 856
rect 189374 800 190310 856
rect 190478 800 191506 856
rect 191674 800 192610 856
rect 192778 800 193806 856
rect 193974 800 194910 856
rect 195078 800 196014 856
rect 196182 800 197210 856
rect 197378 800 198314 856
rect 198482 800 199418 856
rect 199586 800 200614 856
rect 200782 800 201718 856
rect 201886 800 202822 856
rect 202990 800 204018 856
rect 204186 800 205122 856
rect 205290 800 206226 856
rect 206394 800 207422 856
rect 207590 800 208526 856
rect 208694 800 209722 856
rect 209890 800 210826 856
rect 210994 800 211930 856
rect 212098 800 213126 856
rect 213294 800 214230 856
rect 214398 800 215334 856
rect 215502 800 216530 856
rect 216698 800 217634 856
rect 217802 800 218738 856
rect 218906 800 219934 856
rect 220102 800 221038 856
rect 221206 800 222142 856
rect 222310 800 223338 856
rect 223506 800 224442 856
rect 224610 800 225638 856
rect 225806 800 226742 856
rect 226910 800 227846 856
rect 228014 800 229042 856
rect 229210 800 230146 856
rect 230314 800 231250 856
rect 231418 800 232446 856
rect 232614 800 233550 856
rect 233718 800 234654 856
rect 234822 800 235850 856
rect 236018 800 236954 856
rect 237122 800 238150 856
rect 238318 800 239254 856
rect 239422 800 240358 856
rect 240526 800 241554 856
rect 241722 800 242658 856
rect 242826 800 243762 856
rect 243930 800 244958 856
rect 245126 800 246062 856
rect 246230 800 247166 856
rect 247334 800 248362 856
rect 248530 800 249466 856
rect 249634 800 250570 856
rect 250738 800 251766 856
rect 251934 800 252870 856
rect 253038 800 254066 856
rect 254234 800 255170 856
rect 255338 800 256274 856
rect 256442 800 257470 856
rect 257638 800 258574 856
rect 258742 800 259678 856
rect 259846 800 260874 856
rect 261042 800 261978 856
rect 262146 800 263082 856
rect 263250 800 264278 856
rect 264446 800 265382 856
rect 265550 800 266486 856
rect 266654 800 267682 856
rect 267850 800 268786 856
rect 268954 800 269982 856
rect 270150 800 271086 856
rect 271254 800 272190 856
rect 272358 800 273386 856
rect 273554 800 274490 856
rect 274658 800 275594 856
rect 275762 800 276790 856
rect 276958 800 277894 856
rect 278062 800 278998 856
rect 279166 800 280194 856
rect 280362 800 281298 856
rect 281466 800 282494 856
rect 282662 800 283598 856
rect 283766 800 284702 856
rect 284870 800 285898 856
rect 286066 800 287002 856
rect 287170 800 288106 856
rect 288274 800 289302 856
rect 289470 800 290406 856
rect 290574 800 291510 856
rect 291678 800 292706 856
rect 292874 800 293810 856
rect 293978 800 294914 856
rect 295082 800 296110 856
rect 296278 800 297214 856
rect 297382 800 298410 856
rect 298578 800 299514 856
rect 299682 800 300618 856
rect 300786 800 301814 856
rect 301982 800 302918 856
rect 303086 800 304022 856
rect 304190 800 305218 856
rect 305386 800 306322 856
rect 306490 800 307426 856
rect 307594 800 308622 856
rect 308790 800 309726 856
rect 309894 800 310830 856
rect 310998 800 312026 856
rect 312194 800 313130 856
rect 313298 800 314326 856
rect 314494 800 315430 856
rect 315598 800 316534 856
rect 316702 800 317730 856
rect 317898 800 318834 856
rect 319002 800 319938 856
rect 320106 800 321134 856
rect 321302 800 322238 856
rect 322406 800 323342 856
rect 323510 800 324538 856
rect 324706 800 325642 856
rect 325810 800 326746 856
rect 326914 800 327942 856
rect 328110 800 329046 856
rect 329214 800 330242 856
rect 330410 800 331346 856
rect 331514 800 332450 856
rect 332618 800 333646 856
rect 333814 800 334750 856
rect 334918 800 335854 856
rect 336022 800 337050 856
rect 337218 800 338154 856
rect 338322 800 339258 856
rect 339426 800 340454 856
rect 340622 800 341558 856
rect 341726 800 342754 856
rect 342922 800 343858 856
rect 344026 800 344962 856
rect 345130 800 346158 856
rect 346326 800 347262 856
rect 347430 800 348366 856
rect 348534 800 349562 856
rect 349730 800 350666 856
rect 350834 800 351770 856
rect 351938 800 352966 856
rect 353134 800 354070 856
rect 354238 800 355174 856
rect 355342 800 356370 856
rect 356538 800 357474 856
rect 357642 800 358670 856
rect 358838 800 359774 856
rect 359942 800 360878 856
rect 361046 800 362074 856
rect 362242 800 363178 856
rect 363346 800 364282 856
rect 364450 800 365478 856
rect 365646 800 366582 856
rect 366750 800 367686 856
rect 367854 800 368882 856
rect 369050 800 369986 856
rect 370154 800 371090 856
rect 371258 800 372286 856
rect 372454 800 373390 856
rect 373558 800 374586 856
rect 374754 800 375690 856
rect 375858 800 376794 856
rect 376962 800 377990 856
rect 378158 800 379094 856
rect 379262 800 380198 856
rect 380366 800 381394 856
rect 381562 800 382498 856
rect 382666 800 383602 856
rect 383770 800 384798 856
rect 384966 800 385902 856
rect 386070 800 387098 856
rect 387266 800 388202 856
rect 388370 800 389306 856
rect 389474 800 390502 856
rect 390670 800 391606 856
rect 391774 800 392710 856
rect 392878 800 393906 856
rect 394074 800 395010 856
rect 395178 800 396114 856
rect 396282 800 397310 856
rect 397478 800 398414 856
rect 398582 800 399518 856
rect 399686 800 400714 856
rect 400882 800 401818 856
rect 401986 800 403014 856
rect 403182 800 404118 856
rect 404286 800 405222 856
rect 405390 800 406418 856
rect 406586 800 407522 856
rect 407690 800 408626 856
rect 408794 800 409822 856
rect 409990 800 410926 856
rect 411094 800 412030 856
rect 412198 800 413226 856
rect 413394 800 414330 856
rect 414498 800 415434 856
rect 415602 800 416630 856
rect 416798 800 417734 856
rect 417902 800 418930 856
rect 419098 800 420034 856
rect 420202 800 421138 856
rect 421306 800 422334 856
rect 422502 800 423438 856
rect 423606 800 424542 856
rect 424710 800 425738 856
rect 425906 800 426842 856
rect 427010 800 427946 856
rect 428114 800 429142 856
rect 429310 800 430246 856
rect 430414 800 431442 856
rect 431610 800 432546 856
rect 432714 800 433650 856
rect 433818 800 434846 856
rect 435014 800 435950 856
rect 436118 800 437054 856
rect 437222 800 438250 856
rect 438418 800 439354 856
rect 439522 800 440458 856
rect 440626 800 441654 856
rect 441822 800 442758 856
rect 442926 800 443862 856
rect 444030 800 445058 856
rect 445226 800 446162 856
rect 446330 800 447358 856
rect 447526 800 448462 856
rect 448630 800 449566 856
rect 449734 800 450762 856
rect 450930 800 451866 856
rect 452034 800 452970 856
rect 453138 800 454166 856
rect 454334 800 455270 856
rect 455438 800 456374 856
rect 456542 800 457570 856
rect 457738 800 458674 856
rect 458842 800 459778 856
rect 459946 800 460974 856
rect 461142 800 462078 856
rect 462246 800 463274 856
rect 463442 800 464378 856
rect 464546 800 465482 856
rect 465650 800 466678 856
rect 466846 800 467782 856
rect 467950 800 468886 856
rect 469054 800 470082 856
rect 470250 800 471186 856
rect 471354 800 472290 856
rect 472458 800 473486 856
rect 473654 800 474590 856
rect 474758 800 475786 856
rect 475954 800 476890 856
rect 477058 800 477994 856
rect 478162 800 479190 856
rect 479358 800 480294 856
rect 480462 800 481398 856
rect 481566 800 482594 856
rect 482762 800 483698 856
rect 483866 800 484802 856
rect 484970 800 485998 856
rect 486166 800 487102 856
rect 487270 800 488206 856
rect 488374 800 489402 856
rect 489570 800 490506 856
rect 490674 800 491702 856
rect 491870 800 492806 856
rect 492974 800 493910 856
rect 494078 800 495106 856
rect 495274 800 496210 856
rect 496378 800 497314 856
rect 497482 800 498510 856
rect 498678 800 499614 856
rect 499782 800 500718 856
rect 500886 800 501914 856
rect 502082 800 503018 856
rect 503186 800 504122 856
rect 504290 800 505318 856
rect 505486 800 506422 856
rect 506590 800 507618 856
rect 507786 800 508722 856
rect 508890 800 509826 856
rect 509994 800 511022 856
rect 511190 800 512126 856
rect 512294 800 513230 856
rect 513398 800 514426 856
rect 514594 800 515530 856
rect 515698 800 516634 856
rect 516802 800 517830 856
rect 517998 800 518934 856
rect 519102 800 520130 856
rect 520298 800 521234 856
rect 521402 800 522338 856
rect 522506 800 523534 856
rect 523702 800 524638 856
rect 524806 800 525742 856
rect 525910 800 526938 856
rect 527106 800 528042 856
rect 528210 800 529146 856
rect 529314 800 530342 856
rect 530510 800 531446 856
rect 531614 800 532550 856
rect 532718 800 533746 856
rect 533914 800 534850 856
rect 535018 800 536046 856
rect 536214 800 537150 856
rect 537318 800 538254 856
rect 538422 800 539450 856
rect 539618 800 540554 856
rect 540722 800 541658 856
rect 541826 800 542854 856
rect 543022 800 543958 856
rect 544126 800 545062 856
rect 545230 800 546258 856
rect 546426 800 547362 856
rect 547530 800 548466 856
rect 548634 800 549662 856
rect 549830 800 550766 856
rect 550934 800 551962 856
rect 552130 800 553066 856
rect 553234 800 554170 856
rect 554338 800 555366 856
rect 555534 800 556470 856
rect 556638 800 557574 856
<< metal3 >>
rect 0 652672 800 652792
rect 0 590520 800 590640
rect 0 528368 800 528488
rect 0 466216 800 466336
rect 0 404064 800 404184
rect 0 341776 800 341896
rect 0 279624 800 279744
rect 0 217472 800 217592
rect 0 155320 800 155440
rect 0 93168 800 93288
rect 0 31016 800 31136
rect 563200 634992 564000 635112
rect 563200 537344 564000 537464
rect 563200 439560 564000 439680
rect 563200 341912 564000 342032
rect 563200 244128 564000 244248
rect 563200 146480 564000 146600
rect 563200 48832 564000 48952
<< obsm3 >>
rect 4208 851 557599 681665
<< metal4 >>
rect 4208 2128 4528 681680
rect 19568 2128 19888 681680
rect 34928 2128 35248 681680
rect 50288 2128 50608 681680
rect 65648 2128 65968 681680
rect 81008 2128 81328 681680
rect 96368 2128 96688 681680
rect 111728 2128 112048 681680
rect 127088 2128 127408 681680
rect 142448 2128 142768 681680
rect 157808 2128 158128 681680
rect 173168 2128 173488 681680
rect 188528 2128 188848 681680
rect 203888 2128 204208 681680
rect 219248 2128 219568 681680
rect 234608 2128 234928 681680
rect 249968 2128 250288 681680
rect 265328 2128 265648 681680
rect 280688 2128 281008 681680
rect 296048 2128 296368 681680
rect 311408 2128 311728 681680
rect 326768 2128 327088 681680
rect 342128 2128 342448 681680
rect 357488 2128 357808 681680
rect 372848 2128 373168 681680
rect 388208 2128 388528 681680
rect 403568 2128 403888 681680
rect 418928 2128 419248 681680
rect 434288 2128 434608 681680
rect 449648 2128 449968 681680
rect 465008 2128 465328 681680
rect 480368 2128 480688 681680
rect 495728 2128 496048 681680
rect 511088 2128 511408 681680
rect 526448 2128 526768 681680
rect 541808 2128 542128 681680
rect 557168 2128 557488 681680
<< obsm4 >>
rect 45875 33355 50208 679693
rect 50688 33355 65568 679693
rect 66048 33355 80928 679693
rect 81408 33355 96288 679693
rect 96768 33355 111648 679693
rect 112128 33355 127008 679693
rect 127488 33355 142368 679693
rect 142848 33355 157728 679693
rect 158208 33355 173088 679693
rect 173568 33355 188448 679693
rect 188928 33355 203808 679693
rect 204288 33355 219168 679693
rect 219648 33355 234528 679693
rect 235008 33355 249888 679693
rect 250368 33355 265248 679693
rect 265728 33355 280608 679693
rect 281088 33355 295968 679693
rect 296448 33355 311328 679693
rect 311808 33355 326688 679693
rect 327168 33355 342048 679693
rect 342528 33355 357408 679693
rect 357888 33355 372768 679693
rect 373248 33355 388128 679693
rect 388608 33355 400141 679693
<< labels >>
rlabel metal2 s 558826 0 558882 800 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal3 s 563200 146480 564000 146600 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal3 s 0 279624 800 279744 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal3 s 563200 244128 564000 244248 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 543094 683200 543150 684000 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal3 s 0 341776 800 341896 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal3 s 563200 341912 564000 342032 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal3 s 0 404064 800 404184 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s 0 466216 800 466336 6 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal2 s 547786 683200 547842 684000 6 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s 0 528368 800 528488 6 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal2 s 529294 683200 529350 684000 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal2 s 561034 0 561090 800 6 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s 0 590520 800 590640 6 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s 563200 439560 564000 439680 6 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal2 s 562230 0 562286 800 6 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal2 s 552386 683200 552442 684000 6 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal2 s 556986 683200 557042 684000 6 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s 563200 537344 564000 537464 6 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s 563200 634992 564000 635112 6 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal2 s 563334 0 563390 800 6 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal2 s 561586 683200 561642 684000 6 analog_io[29]
port 22 nsew signal bidirectional
rlabel metal3 s 0 31016 800 31136 6 analog_io[2]
port 23 nsew signal bidirectional
rlabel metal3 s 0 652672 800 652792 6 analog_io[30]
port 24 nsew signal bidirectional
rlabel metal3 s 0 93168 800 93288 6 analog_io[3]
port 25 nsew signal bidirectional
rlabel metal2 s 559930 0 559986 800 6 analog_io[4]
port 26 nsew signal bidirectional
rlabel metal2 s 533894 683200 533950 684000 6 analog_io[5]
port 27 nsew signal bidirectional
rlabel metal3 s 563200 48832 564000 48952 6 analog_io[6]
port 28 nsew signal bidirectional
rlabel metal2 s 538494 683200 538550 684000 6 analog_io[7]
port 29 nsew signal bidirectional
rlabel metal3 s 0 155320 800 155440 6 analog_io[8]
port 30 nsew signal bidirectional
rlabel metal3 s 0 217472 800 217592 6 analog_io[9]
port 31 nsew signal bidirectional
rlabel metal2 s 2318 683200 2374 684000 6 io_in[0]
port 32 nsew signal input
rlabel metal2 s 140962 683200 141018 684000 6 io_in[10]
port 33 nsew signal input
rlabel metal2 s 154854 683200 154910 684000 6 io_in[11]
port 34 nsew signal input
rlabel metal2 s 168654 683200 168710 684000 6 io_in[12]
port 35 nsew signal input
rlabel metal2 s 182546 683200 182602 684000 6 io_in[13]
port 36 nsew signal input
rlabel metal2 s 196438 683200 196494 684000 6 io_in[14]
port 37 nsew signal input
rlabel metal2 s 210330 683200 210386 684000 6 io_in[15]
port 38 nsew signal input
rlabel metal2 s 224130 683200 224186 684000 6 io_in[16]
port 39 nsew signal input
rlabel metal2 s 238022 683200 238078 684000 6 io_in[17]
port 40 nsew signal input
rlabel metal2 s 251914 683200 251970 684000 6 io_in[18]
port 41 nsew signal input
rlabel metal2 s 265806 683200 265862 684000 6 io_in[19]
port 42 nsew signal input
rlabel metal2 s 16118 683200 16174 684000 6 io_in[1]
port 43 nsew signal input
rlabel metal2 s 279606 683200 279662 684000 6 io_in[20]
port 44 nsew signal input
rlabel metal2 s 293498 683200 293554 684000 6 io_in[21]
port 45 nsew signal input
rlabel metal2 s 307390 683200 307446 684000 6 io_in[22]
port 46 nsew signal input
rlabel metal2 s 321190 683200 321246 684000 6 io_in[23]
port 47 nsew signal input
rlabel metal2 s 335082 683200 335138 684000 6 io_in[24]
port 48 nsew signal input
rlabel metal2 s 348974 683200 349030 684000 6 io_in[25]
port 49 nsew signal input
rlabel metal2 s 362866 683200 362922 684000 6 io_in[26]
port 50 nsew signal input
rlabel metal2 s 376666 683200 376722 684000 6 io_in[27]
port 51 nsew signal input
rlabel metal2 s 390558 683200 390614 684000 6 io_in[28]
port 52 nsew signal input
rlabel metal2 s 404450 683200 404506 684000 6 io_in[29]
port 53 nsew signal input
rlabel metal2 s 30010 683200 30066 684000 6 io_in[2]
port 54 nsew signal input
rlabel metal2 s 418342 683200 418398 684000 6 io_in[30]
port 55 nsew signal input
rlabel metal2 s 432142 683200 432198 684000 6 io_in[31]
port 56 nsew signal input
rlabel metal2 s 446034 683200 446090 684000 6 io_in[32]
port 57 nsew signal input
rlabel metal2 s 459926 683200 459982 684000 6 io_in[33]
port 58 nsew signal input
rlabel metal2 s 473818 683200 473874 684000 6 io_in[34]
port 59 nsew signal input
rlabel metal2 s 487618 683200 487674 684000 6 io_in[35]
port 60 nsew signal input
rlabel metal2 s 501510 683200 501566 684000 6 io_in[36]
port 61 nsew signal input
rlabel metal2 s 515402 683200 515458 684000 6 io_in[37]
port 62 nsew signal input
rlabel metal2 s 43902 683200 43958 684000 6 io_in[3]
port 63 nsew signal input
rlabel metal2 s 57702 683200 57758 684000 6 io_in[4]
port 64 nsew signal input
rlabel metal2 s 71594 683200 71650 684000 6 io_in[5]
port 65 nsew signal input
rlabel metal2 s 85486 683200 85542 684000 6 io_in[6]
port 66 nsew signal input
rlabel metal2 s 99378 683200 99434 684000 6 io_in[7]
port 67 nsew signal input
rlabel metal2 s 113178 683200 113234 684000 6 io_in[8]
port 68 nsew signal input
rlabel metal2 s 127070 683200 127126 684000 6 io_in[9]
port 69 nsew signal input
rlabel metal2 s 6918 683200 6974 684000 6 io_oeb[0]
port 70 nsew signal output
rlabel metal2 s 145562 683200 145618 684000 6 io_oeb[10]
port 71 nsew signal output
rlabel metal2 s 159454 683200 159510 684000 6 io_oeb[11]
port 72 nsew signal output
rlabel metal2 s 173346 683200 173402 684000 6 io_oeb[12]
port 73 nsew signal output
rlabel metal2 s 187146 683200 187202 684000 6 io_oeb[13]
port 74 nsew signal output
rlabel metal2 s 201038 683200 201094 684000 6 io_oeb[14]
port 75 nsew signal output
rlabel metal2 s 214930 683200 214986 684000 6 io_oeb[15]
port 76 nsew signal output
rlabel metal2 s 228822 683200 228878 684000 6 io_oeb[16]
port 77 nsew signal output
rlabel metal2 s 242622 683200 242678 684000 6 io_oeb[17]
port 78 nsew signal output
rlabel metal2 s 256514 683200 256570 684000 6 io_oeb[18]
port 79 nsew signal output
rlabel metal2 s 270406 683200 270462 684000 6 io_oeb[19]
port 80 nsew signal output
rlabel metal2 s 20718 683200 20774 684000 6 io_oeb[1]
port 81 nsew signal output
rlabel metal2 s 284298 683200 284354 684000 6 io_oeb[20]
port 82 nsew signal output
rlabel metal2 s 298098 683200 298154 684000 6 io_oeb[21]
port 83 nsew signal output
rlabel metal2 s 311990 683200 312046 684000 6 io_oeb[22]
port 84 nsew signal output
rlabel metal2 s 325882 683200 325938 684000 6 io_oeb[23]
port 85 nsew signal output
rlabel metal2 s 339682 683200 339738 684000 6 io_oeb[24]
port 86 nsew signal output
rlabel metal2 s 353574 683200 353630 684000 6 io_oeb[25]
port 87 nsew signal output
rlabel metal2 s 367466 683200 367522 684000 6 io_oeb[26]
port 88 nsew signal output
rlabel metal2 s 381358 683200 381414 684000 6 io_oeb[27]
port 89 nsew signal output
rlabel metal2 s 395158 683200 395214 684000 6 io_oeb[28]
port 90 nsew signal output
rlabel metal2 s 409050 683200 409106 684000 6 io_oeb[29]
port 91 nsew signal output
rlabel metal2 s 34610 683200 34666 684000 6 io_oeb[2]
port 92 nsew signal output
rlabel metal2 s 422942 683200 422998 684000 6 io_oeb[30]
port 93 nsew signal output
rlabel metal2 s 436834 683200 436890 684000 6 io_oeb[31]
port 94 nsew signal output
rlabel metal2 s 450634 683200 450690 684000 6 io_oeb[32]
port 95 nsew signal output
rlabel metal2 s 464526 683200 464582 684000 6 io_oeb[33]
port 96 nsew signal output
rlabel metal2 s 478418 683200 478474 684000 6 io_oeb[34]
port 97 nsew signal output
rlabel metal2 s 492310 683200 492366 684000 6 io_oeb[35]
port 98 nsew signal output
rlabel metal2 s 506110 683200 506166 684000 6 io_oeb[36]
port 99 nsew signal output
rlabel metal2 s 520002 683200 520058 684000 6 io_oeb[37]
port 100 nsew signal output
rlabel metal2 s 48502 683200 48558 684000 6 io_oeb[3]
port 101 nsew signal output
rlabel metal2 s 62394 683200 62450 684000 6 io_oeb[4]
port 102 nsew signal output
rlabel metal2 s 76194 683200 76250 684000 6 io_oeb[5]
port 103 nsew signal output
rlabel metal2 s 90086 683200 90142 684000 6 io_oeb[6]
port 104 nsew signal output
rlabel metal2 s 103978 683200 104034 684000 6 io_oeb[7]
port 105 nsew signal output
rlabel metal2 s 117870 683200 117926 684000 6 io_oeb[8]
port 106 nsew signal output
rlabel metal2 s 131670 683200 131726 684000 6 io_oeb[9]
port 107 nsew signal output
rlabel metal2 s 11518 683200 11574 684000 6 io_out[0]
port 108 nsew signal output
rlabel metal2 s 150162 683200 150218 684000 6 io_out[10]
port 109 nsew signal output
rlabel metal2 s 164054 683200 164110 684000 6 io_out[11]
port 110 nsew signal output
rlabel metal2 s 177946 683200 178002 684000 6 io_out[12]
port 111 nsew signal output
rlabel metal2 s 191838 683200 191894 684000 6 io_out[13]
port 112 nsew signal output
rlabel metal2 s 205638 683200 205694 684000 6 io_out[14]
port 113 nsew signal output
rlabel metal2 s 219530 683200 219586 684000 6 io_out[15]
port 114 nsew signal output
rlabel metal2 s 233422 683200 233478 684000 6 io_out[16]
port 115 nsew signal output
rlabel metal2 s 247314 683200 247370 684000 6 io_out[17]
port 116 nsew signal output
rlabel metal2 s 261114 683200 261170 684000 6 io_out[18]
port 117 nsew signal output
rlabel metal2 s 275006 683200 275062 684000 6 io_out[19]
port 118 nsew signal output
rlabel metal2 s 25410 683200 25466 684000 6 io_out[1]
port 119 nsew signal output
rlabel metal2 s 288898 683200 288954 684000 6 io_out[20]
port 120 nsew signal output
rlabel metal2 s 302698 683200 302754 684000 6 io_out[21]
port 121 nsew signal output
rlabel metal2 s 316590 683200 316646 684000 6 io_out[22]
port 122 nsew signal output
rlabel metal2 s 330482 683200 330538 684000 6 io_out[23]
port 123 nsew signal output
rlabel metal2 s 344374 683200 344430 684000 6 io_out[24]
port 124 nsew signal output
rlabel metal2 s 358174 683200 358230 684000 6 io_out[25]
port 125 nsew signal output
rlabel metal2 s 372066 683200 372122 684000 6 io_out[26]
port 126 nsew signal output
rlabel metal2 s 385958 683200 386014 684000 6 io_out[27]
port 127 nsew signal output
rlabel metal2 s 399850 683200 399906 684000 6 io_out[28]
port 128 nsew signal output
rlabel metal2 s 413650 683200 413706 684000 6 io_out[29]
port 129 nsew signal output
rlabel metal2 s 39210 683200 39266 684000 6 io_out[2]
port 130 nsew signal output
rlabel metal2 s 427542 683200 427598 684000 6 io_out[30]
port 131 nsew signal output
rlabel metal2 s 441434 683200 441490 684000 6 io_out[31]
port 132 nsew signal output
rlabel metal2 s 455326 683200 455382 684000 6 io_out[32]
port 133 nsew signal output
rlabel metal2 s 469126 683200 469182 684000 6 io_out[33]
port 134 nsew signal output
rlabel metal2 s 483018 683200 483074 684000 6 io_out[34]
port 135 nsew signal output
rlabel metal2 s 496910 683200 496966 684000 6 io_out[35]
port 136 nsew signal output
rlabel metal2 s 510802 683200 510858 684000 6 io_out[36]
port 137 nsew signal output
rlabel metal2 s 524602 683200 524658 684000 6 io_out[37]
port 138 nsew signal output
rlabel metal2 s 53102 683200 53158 684000 6 io_out[3]
port 139 nsew signal output
rlabel metal2 s 66994 683200 67050 684000 6 io_out[4]
port 140 nsew signal output
rlabel metal2 s 80886 683200 80942 684000 6 io_out[5]
port 141 nsew signal output
rlabel metal2 s 94686 683200 94742 684000 6 io_out[6]
port 142 nsew signal output
rlabel metal2 s 108578 683200 108634 684000 6 io_out[7]
port 143 nsew signal output
rlabel metal2 s 122470 683200 122526 684000 6 io_out[8]
port 144 nsew signal output
rlabel metal2 s 136362 683200 136418 684000 6 io_out[9]
port 145 nsew signal output
rlabel metal2 s 121090 0 121146 800 6 la_data_in[0]
port 146 nsew signal input
rlabel metal2 s 462134 0 462190 800 6 la_data_in[100]
port 147 nsew signal input
rlabel metal2 s 465538 0 465594 800 6 la_data_in[101]
port 148 nsew signal input
rlabel metal2 s 468942 0 468998 800 6 la_data_in[102]
port 149 nsew signal input
rlabel metal2 s 472346 0 472402 800 6 la_data_in[103]
port 150 nsew signal input
rlabel metal2 s 475842 0 475898 800 6 la_data_in[104]
port 151 nsew signal input
rlabel metal2 s 479246 0 479302 800 6 la_data_in[105]
port 152 nsew signal input
rlabel metal2 s 482650 0 482706 800 6 la_data_in[106]
port 153 nsew signal input
rlabel metal2 s 486054 0 486110 800 6 la_data_in[107]
port 154 nsew signal input
rlabel metal2 s 489458 0 489514 800 6 la_data_in[108]
port 155 nsew signal input
rlabel metal2 s 492862 0 492918 800 6 la_data_in[109]
port 156 nsew signal input
rlabel metal2 s 155130 0 155186 800 6 la_data_in[10]
port 157 nsew signal input
rlabel metal2 s 496266 0 496322 800 6 la_data_in[110]
port 158 nsew signal input
rlabel metal2 s 499670 0 499726 800 6 la_data_in[111]
port 159 nsew signal input
rlabel metal2 s 503074 0 503130 800 6 la_data_in[112]
port 160 nsew signal input
rlabel metal2 s 506478 0 506534 800 6 la_data_in[113]
port 161 nsew signal input
rlabel metal2 s 509882 0 509938 800 6 la_data_in[114]
port 162 nsew signal input
rlabel metal2 s 513286 0 513342 800 6 la_data_in[115]
port 163 nsew signal input
rlabel metal2 s 516690 0 516746 800 6 la_data_in[116]
port 164 nsew signal input
rlabel metal2 s 520186 0 520242 800 6 la_data_in[117]
port 165 nsew signal input
rlabel metal2 s 523590 0 523646 800 6 la_data_in[118]
port 166 nsew signal input
rlabel metal2 s 526994 0 527050 800 6 la_data_in[119]
port 167 nsew signal input
rlabel metal2 s 158534 0 158590 800 6 la_data_in[11]
port 168 nsew signal input
rlabel metal2 s 530398 0 530454 800 6 la_data_in[120]
port 169 nsew signal input
rlabel metal2 s 533802 0 533858 800 6 la_data_in[121]
port 170 nsew signal input
rlabel metal2 s 537206 0 537262 800 6 la_data_in[122]
port 171 nsew signal input
rlabel metal2 s 540610 0 540666 800 6 la_data_in[123]
port 172 nsew signal input
rlabel metal2 s 544014 0 544070 800 6 la_data_in[124]
port 173 nsew signal input
rlabel metal2 s 547418 0 547474 800 6 la_data_in[125]
port 174 nsew signal input
rlabel metal2 s 550822 0 550878 800 6 la_data_in[126]
port 175 nsew signal input
rlabel metal2 s 554226 0 554282 800 6 la_data_in[127]
port 176 nsew signal input
rlabel metal2 s 161938 0 161994 800 6 la_data_in[12]
port 177 nsew signal input
rlabel metal2 s 165434 0 165490 800 6 la_data_in[13]
port 178 nsew signal input
rlabel metal2 s 168838 0 168894 800 6 la_data_in[14]
port 179 nsew signal input
rlabel metal2 s 172242 0 172298 800 6 la_data_in[15]
port 180 nsew signal input
rlabel metal2 s 175646 0 175702 800 6 la_data_in[16]
port 181 nsew signal input
rlabel metal2 s 179050 0 179106 800 6 la_data_in[17]
port 182 nsew signal input
rlabel metal2 s 182454 0 182510 800 6 la_data_in[18]
port 183 nsew signal input
rlabel metal2 s 185858 0 185914 800 6 la_data_in[19]
port 184 nsew signal input
rlabel metal2 s 124494 0 124550 800 6 la_data_in[1]
port 185 nsew signal input
rlabel metal2 s 189262 0 189318 800 6 la_data_in[20]
port 186 nsew signal input
rlabel metal2 s 192666 0 192722 800 6 la_data_in[21]
port 187 nsew signal input
rlabel metal2 s 196070 0 196126 800 6 la_data_in[22]
port 188 nsew signal input
rlabel metal2 s 199474 0 199530 800 6 la_data_in[23]
port 189 nsew signal input
rlabel metal2 s 202878 0 202934 800 6 la_data_in[24]
port 190 nsew signal input
rlabel metal2 s 206282 0 206338 800 6 la_data_in[25]
port 191 nsew signal input
rlabel metal2 s 209778 0 209834 800 6 la_data_in[26]
port 192 nsew signal input
rlabel metal2 s 213182 0 213238 800 6 la_data_in[27]
port 193 nsew signal input
rlabel metal2 s 216586 0 216642 800 6 la_data_in[28]
port 194 nsew signal input
rlabel metal2 s 219990 0 220046 800 6 la_data_in[29]
port 195 nsew signal input
rlabel metal2 s 127898 0 127954 800 6 la_data_in[2]
port 196 nsew signal input
rlabel metal2 s 223394 0 223450 800 6 la_data_in[30]
port 197 nsew signal input
rlabel metal2 s 226798 0 226854 800 6 la_data_in[31]
port 198 nsew signal input
rlabel metal2 s 230202 0 230258 800 6 la_data_in[32]
port 199 nsew signal input
rlabel metal2 s 233606 0 233662 800 6 la_data_in[33]
port 200 nsew signal input
rlabel metal2 s 237010 0 237066 800 6 la_data_in[34]
port 201 nsew signal input
rlabel metal2 s 240414 0 240470 800 6 la_data_in[35]
port 202 nsew signal input
rlabel metal2 s 243818 0 243874 800 6 la_data_in[36]
port 203 nsew signal input
rlabel metal2 s 247222 0 247278 800 6 la_data_in[37]
port 204 nsew signal input
rlabel metal2 s 250626 0 250682 800 6 la_data_in[38]
port 205 nsew signal input
rlabel metal2 s 254122 0 254178 800 6 la_data_in[39]
port 206 nsew signal input
rlabel metal2 s 131302 0 131358 800 6 la_data_in[3]
port 207 nsew signal input
rlabel metal2 s 257526 0 257582 800 6 la_data_in[40]
port 208 nsew signal input
rlabel metal2 s 260930 0 260986 800 6 la_data_in[41]
port 209 nsew signal input
rlabel metal2 s 264334 0 264390 800 6 la_data_in[42]
port 210 nsew signal input
rlabel metal2 s 267738 0 267794 800 6 la_data_in[43]
port 211 nsew signal input
rlabel metal2 s 271142 0 271198 800 6 la_data_in[44]
port 212 nsew signal input
rlabel metal2 s 274546 0 274602 800 6 la_data_in[45]
port 213 nsew signal input
rlabel metal2 s 277950 0 278006 800 6 la_data_in[46]
port 214 nsew signal input
rlabel metal2 s 281354 0 281410 800 6 la_data_in[47]
port 215 nsew signal input
rlabel metal2 s 284758 0 284814 800 6 la_data_in[48]
port 216 nsew signal input
rlabel metal2 s 288162 0 288218 800 6 la_data_in[49]
port 217 nsew signal input
rlabel metal2 s 134706 0 134762 800 6 la_data_in[4]
port 218 nsew signal input
rlabel metal2 s 291566 0 291622 800 6 la_data_in[50]
port 219 nsew signal input
rlabel metal2 s 294970 0 295026 800 6 la_data_in[51]
port 220 nsew signal input
rlabel metal2 s 298466 0 298522 800 6 la_data_in[52]
port 221 nsew signal input
rlabel metal2 s 301870 0 301926 800 6 la_data_in[53]
port 222 nsew signal input
rlabel metal2 s 305274 0 305330 800 6 la_data_in[54]
port 223 nsew signal input
rlabel metal2 s 308678 0 308734 800 6 la_data_in[55]
port 224 nsew signal input
rlabel metal2 s 312082 0 312138 800 6 la_data_in[56]
port 225 nsew signal input
rlabel metal2 s 315486 0 315542 800 6 la_data_in[57]
port 226 nsew signal input
rlabel metal2 s 318890 0 318946 800 6 la_data_in[58]
port 227 nsew signal input
rlabel metal2 s 322294 0 322350 800 6 la_data_in[59]
port 228 nsew signal input
rlabel metal2 s 138110 0 138166 800 6 la_data_in[5]
port 229 nsew signal input
rlabel metal2 s 325698 0 325754 800 6 la_data_in[60]
port 230 nsew signal input
rlabel metal2 s 329102 0 329158 800 6 la_data_in[61]
port 231 nsew signal input
rlabel metal2 s 332506 0 332562 800 6 la_data_in[62]
port 232 nsew signal input
rlabel metal2 s 335910 0 335966 800 6 la_data_in[63]
port 233 nsew signal input
rlabel metal2 s 339314 0 339370 800 6 la_data_in[64]
port 234 nsew signal input
rlabel metal2 s 342810 0 342866 800 6 la_data_in[65]
port 235 nsew signal input
rlabel metal2 s 346214 0 346270 800 6 la_data_in[66]
port 236 nsew signal input
rlabel metal2 s 349618 0 349674 800 6 la_data_in[67]
port 237 nsew signal input
rlabel metal2 s 353022 0 353078 800 6 la_data_in[68]
port 238 nsew signal input
rlabel metal2 s 356426 0 356482 800 6 la_data_in[69]
port 239 nsew signal input
rlabel metal2 s 141514 0 141570 800 6 la_data_in[6]
port 240 nsew signal input
rlabel metal2 s 359830 0 359886 800 6 la_data_in[70]
port 241 nsew signal input
rlabel metal2 s 363234 0 363290 800 6 la_data_in[71]
port 242 nsew signal input
rlabel metal2 s 366638 0 366694 800 6 la_data_in[72]
port 243 nsew signal input
rlabel metal2 s 370042 0 370098 800 6 la_data_in[73]
port 244 nsew signal input
rlabel metal2 s 373446 0 373502 800 6 la_data_in[74]
port 245 nsew signal input
rlabel metal2 s 376850 0 376906 800 6 la_data_in[75]
port 246 nsew signal input
rlabel metal2 s 380254 0 380310 800 6 la_data_in[76]
port 247 nsew signal input
rlabel metal2 s 383658 0 383714 800 6 la_data_in[77]
port 248 nsew signal input
rlabel metal2 s 387154 0 387210 800 6 la_data_in[78]
port 249 nsew signal input
rlabel metal2 s 390558 0 390614 800 6 la_data_in[79]
port 250 nsew signal input
rlabel metal2 s 144918 0 144974 800 6 la_data_in[7]
port 251 nsew signal input
rlabel metal2 s 393962 0 394018 800 6 la_data_in[80]
port 252 nsew signal input
rlabel metal2 s 397366 0 397422 800 6 la_data_in[81]
port 253 nsew signal input
rlabel metal2 s 400770 0 400826 800 6 la_data_in[82]
port 254 nsew signal input
rlabel metal2 s 404174 0 404230 800 6 la_data_in[83]
port 255 nsew signal input
rlabel metal2 s 407578 0 407634 800 6 la_data_in[84]
port 256 nsew signal input
rlabel metal2 s 410982 0 411038 800 6 la_data_in[85]
port 257 nsew signal input
rlabel metal2 s 414386 0 414442 800 6 la_data_in[86]
port 258 nsew signal input
rlabel metal2 s 417790 0 417846 800 6 la_data_in[87]
port 259 nsew signal input
rlabel metal2 s 421194 0 421250 800 6 la_data_in[88]
port 260 nsew signal input
rlabel metal2 s 424598 0 424654 800 6 la_data_in[89]
port 261 nsew signal input
rlabel metal2 s 148322 0 148378 800 6 la_data_in[8]
port 262 nsew signal input
rlabel metal2 s 428002 0 428058 800 6 la_data_in[90]
port 263 nsew signal input
rlabel metal2 s 431498 0 431554 800 6 la_data_in[91]
port 264 nsew signal input
rlabel metal2 s 434902 0 434958 800 6 la_data_in[92]
port 265 nsew signal input
rlabel metal2 s 438306 0 438362 800 6 la_data_in[93]
port 266 nsew signal input
rlabel metal2 s 441710 0 441766 800 6 la_data_in[94]
port 267 nsew signal input
rlabel metal2 s 445114 0 445170 800 6 la_data_in[95]
port 268 nsew signal input
rlabel metal2 s 448518 0 448574 800 6 la_data_in[96]
port 269 nsew signal input
rlabel metal2 s 451922 0 451978 800 6 la_data_in[97]
port 270 nsew signal input
rlabel metal2 s 455326 0 455382 800 6 la_data_in[98]
port 271 nsew signal input
rlabel metal2 s 458730 0 458786 800 6 la_data_in[99]
port 272 nsew signal input
rlabel metal2 s 151726 0 151782 800 6 la_data_in[9]
port 273 nsew signal input
rlabel metal2 s 122194 0 122250 800 6 la_data_out[0]
port 274 nsew signal output
rlabel metal2 s 463330 0 463386 800 6 la_data_out[100]
port 275 nsew signal output
rlabel metal2 s 466734 0 466790 800 6 la_data_out[101]
port 276 nsew signal output
rlabel metal2 s 470138 0 470194 800 6 la_data_out[102]
port 277 nsew signal output
rlabel metal2 s 473542 0 473598 800 6 la_data_out[103]
port 278 nsew signal output
rlabel metal2 s 476946 0 477002 800 6 la_data_out[104]
port 279 nsew signal output
rlabel metal2 s 480350 0 480406 800 6 la_data_out[105]
port 280 nsew signal output
rlabel metal2 s 483754 0 483810 800 6 la_data_out[106]
port 281 nsew signal output
rlabel metal2 s 487158 0 487214 800 6 la_data_out[107]
port 282 nsew signal output
rlabel metal2 s 490562 0 490618 800 6 la_data_out[108]
port 283 nsew signal output
rlabel metal2 s 493966 0 494022 800 6 la_data_out[109]
port 284 nsew signal output
rlabel metal2 s 156326 0 156382 800 6 la_data_out[10]
port 285 nsew signal output
rlabel metal2 s 497370 0 497426 800 6 la_data_out[110]
port 286 nsew signal output
rlabel metal2 s 500774 0 500830 800 6 la_data_out[111]
port 287 nsew signal output
rlabel metal2 s 504178 0 504234 800 6 la_data_out[112]
port 288 nsew signal output
rlabel metal2 s 507674 0 507730 800 6 la_data_out[113]
port 289 nsew signal output
rlabel metal2 s 511078 0 511134 800 6 la_data_out[114]
port 290 nsew signal output
rlabel metal2 s 514482 0 514538 800 6 la_data_out[115]
port 291 nsew signal output
rlabel metal2 s 517886 0 517942 800 6 la_data_out[116]
port 292 nsew signal output
rlabel metal2 s 521290 0 521346 800 6 la_data_out[117]
port 293 nsew signal output
rlabel metal2 s 524694 0 524750 800 6 la_data_out[118]
port 294 nsew signal output
rlabel metal2 s 528098 0 528154 800 6 la_data_out[119]
port 295 nsew signal output
rlabel metal2 s 159730 0 159786 800 6 la_data_out[11]
port 296 nsew signal output
rlabel metal2 s 531502 0 531558 800 6 la_data_out[120]
port 297 nsew signal output
rlabel metal2 s 534906 0 534962 800 6 la_data_out[121]
port 298 nsew signal output
rlabel metal2 s 538310 0 538366 800 6 la_data_out[122]
port 299 nsew signal output
rlabel metal2 s 541714 0 541770 800 6 la_data_out[123]
port 300 nsew signal output
rlabel metal2 s 545118 0 545174 800 6 la_data_out[124]
port 301 nsew signal output
rlabel metal2 s 548522 0 548578 800 6 la_data_out[125]
port 302 nsew signal output
rlabel metal2 s 552018 0 552074 800 6 la_data_out[126]
port 303 nsew signal output
rlabel metal2 s 555422 0 555478 800 6 la_data_out[127]
port 304 nsew signal output
rlabel metal2 s 163134 0 163190 800 6 la_data_out[12]
port 305 nsew signal output
rlabel metal2 s 166538 0 166594 800 6 la_data_out[13]
port 306 nsew signal output
rlabel metal2 s 169942 0 169998 800 6 la_data_out[14]
port 307 nsew signal output
rlabel metal2 s 173346 0 173402 800 6 la_data_out[15]
port 308 nsew signal output
rlabel metal2 s 176750 0 176806 800 6 la_data_out[16]
port 309 nsew signal output
rlabel metal2 s 180154 0 180210 800 6 la_data_out[17]
port 310 nsew signal output
rlabel metal2 s 183558 0 183614 800 6 la_data_out[18]
port 311 nsew signal output
rlabel metal2 s 186962 0 187018 800 6 la_data_out[19]
port 312 nsew signal output
rlabel metal2 s 125598 0 125654 800 6 la_data_out[1]
port 313 nsew signal output
rlabel metal2 s 190366 0 190422 800 6 la_data_out[20]
port 314 nsew signal output
rlabel metal2 s 193862 0 193918 800 6 la_data_out[21]
port 315 nsew signal output
rlabel metal2 s 197266 0 197322 800 6 la_data_out[22]
port 316 nsew signal output
rlabel metal2 s 200670 0 200726 800 6 la_data_out[23]
port 317 nsew signal output
rlabel metal2 s 204074 0 204130 800 6 la_data_out[24]
port 318 nsew signal output
rlabel metal2 s 207478 0 207534 800 6 la_data_out[25]
port 319 nsew signal output
rlabel metal2 s 210882 0 210938 800 6 la_data_out[26]
port 320 nsew signal output
rlabel metal2 s 214286 0 214342 800 6 la_data_out[27]
port 321 nsew signal output
rlabel metal2 s 217690 0 217746 800 6 la_data_out[28]
port 322 nsew signal output
rlabel metal2 s 221094 0 221150 800 6 la_data_out[29]
port 323 nsew signal output
rlabel metal2 s 129002 0 129058 800 6 la_data_out[2]
port 324 nsew signal output
rlabel metal2 s 224498 0 224554 800 6 la_data_out[30]
port 325 nsew signal output
rlabel metal2 s 227902 0 227958 800 6 la_data_out[31]
port 326 nsew signal output
rlabel metal2 s 231306 0 231362 800 6 la_data_out[32]
port 327 nsew signal output
rlabel metal2 s 234710 0 234766 800 6 la_data_out[33]
port 328 nsew signal output
rlabel metal2 s 238206 0 238262 800 6 la_data_out[34]
port 329 nsew signal output
rlabel metal2 s 241610 0 241666 800 6 la_data_out[35]
port 330 nsew signal output
rlabel metal2 s 245014 0 245070 800 6 la_data_out[36]
port 331 nsew signal output
rlabel metal2 s 248418 0 248474 800 6 la_data_out[37]
port 332 nsew signal output
rlabel metal2 s 251822 0 251878 800 6 la_data_out[38]
port 333 nsew signal output
rlabel metal2 s 255226 0 255282 800 6 la_data_out[39]
port 334 nsew signal output
rlabel metal2 s 132406 0 132462 800 6 la_data_out[3]
port 335 nsew signal output
rlabel metal2 s 258630 0 258686 800 6 la_data_out[40]
port 336 nsew signal output
rlabel metal2 s 262034 0 262090 800 6 la_data_out[41]
port 337 nsew signal output
rlabel metal2 s 265438 0 265494 800 6 la_data_out[42]
port 338 nsew signal output
rlabel metal2 s 268842 0 268898 800 6 la_data_out[43]
port 339 nsew signal output
rlabel metal2 s 272246 0 272302 800 6 la_data_out[44]
port 340 nsew signal output
rlabel metal2 s 275650 0 275706 800 6 la_data_out[45]
port 341 nsew signal output
rlabel metal2 s 279054 0 279110 800 6 la_data_out[46]
port 342 nsew signal output
rlabel metal2 s 282550 0 282606 800 6 la_data_out[47]
port 343 nsew signal output
rlabel metal2 s 285954 0 286010 800 6 la_data_out[48]
port 344 nsew signal output
rlabel metal2 s 289358 0 289414 800 6 la_data_out[49]
port 345 nsew signal output
rlabel metal2 s 135810 0 135866 800 6 la_data_out[4]
port 346 nsew signal output
rlabel metal2 s 292762 0 292818 800 6 la_data_out[50]
port 347 nsew signal output
rlabel metal2 s 296166 0 296222 800 6 la_data_out[51]
port 348 nsew signal output
rlabel metal2 s 299570 0 299626 800 6 la_data_out[52]
port 349 nsew signal output
rlabel metal2 s 302974 0 303030 800 6 la_data_out[53]
port 350 nsew signal output
rlabel metal2 s 306378 0 306434 800 6 la_data_out[54]
port 351 nsew signal output
rlabel metal2 s 309782 0 309838 800 6 la_data_out[55]
port 352 nsew signal output
rlabel metal2 s 313186 0 313242 800 6 la_data_out[56]
port 353 nsew signal output
rlabel metal2 s 316590 0 316646 800 6 la_data_out[57]
port 354 nsew signal output
rlabel metal2 s 319994 0 320050 800 6 la_data_out[58]
port 355 nsew signal output
rlabel metal2 s 323398 0 323454 800 6 la_data_out[59]
port 356 nsew signal output
rlabel metal2 s 139214 0 139270 800 6 la_data_out[5]
port 357 nsew signal output
rlabel metal2 s 326802 0 326858 800 6 la_data_out[60]
port 358 nsew signal output
rlabel metal2 s 330298 0 330354 800 6 la_data_out[61]
port 359 nsew signal output
rlabel metal2 s 333702 0 333758 800 6 la_data_out[62]
port 360 nsew signal output
rlabel metal2 s 337106 0 337162 800 6 la_data_out[63]
port 361 nsew signal output
rlabel metal2 s 340510 0 340566 800 6 la_data_out[64]
port 362 nsew signal output
rlabel metal2 s 343914 0 343970 800 6 la_data_out[65]
port 363 nsew signal output
rlabel metal2 s 347318 0 347374 800 6 la_data_out[66]
port 364 nsew signal output
rlabel metal2 s 350722 0 350778 800 6 la_data_out[67]
port 365 nsew signal output
rlabel metal2 s 354126 0 354182 800 6 la_data_out[68]
port 366 nsew signal output
rlabel metal2 s 357530 0 357586 800 6 la_data_out[69]
port 367 nsew signal output
rlabel metal2 s 142618 0 142674 800 6 la_data_out[6]
port 368 nsew signal output
rlabel metal2 s 360934 0 360990 800 6 la_data_out[70]
port 369 nsew signal output
rlabel metal2 s 364338 0 364394 800 6 la_data_out[71]
port 370 nsew signal output
rlabel metal2 s 367742 0 367798 800 6 la_data_out[72]
port 371 nsew signal output
rlabel metal2 s 371146 0 371202 800 6 la_data_out[73]
port 372 nsew signal output
rlabel metal2 s 374642 0 374698 800 6 la_data_out[74]
port 373 nsew signal output
rlabel metal2 s 378046 0 378102 800 6 la_data_out[75]
port 374 nsew signal output
rlabel metal2 s 381450 0 381506 800 6 la_data_out[76]
port 375 nsew signal output
rlabel metal2 s 384854 0 384910 800 6 la_data_out[77]
port 376 nsew signal output
rlabel metal2 s 388258 0 388314 800 6 la_data_out[78]
port 377 nsew signal output
rlabel metal2 s 391662 0 391718 800 6 la_data_out[79]
port 378 nsew signal output
rlabel metal2 s 146022 0 146078 800 6 la_data_out[7]
port 379 nsew signal output
rlabel metal2 s 395066 0 395122 800 6 la_data_out[80]
port 380 nsew signal output
rlabel metal2 s 398470 0 398526 800 6 la_data_out[81]
port 381 nsew signal output
rlabel metal2 s 401874 0 401930 800 6 la_data_out[82]
port 382 nsew signal output
rlabel metal2 s 405278 0 405334 800 6 la_data_out[83]
port 383 nsew signal output
rlabel metal2 s 408682 0 408738 800 6 la_data_out[84]
port 384 nsew signal output
rlabel metal2 s 412086 0 412142 800 6 la_data_out[85]
port 385 nsew signal output
rlabel metal2 s 415490 0 415546 800 6 la_data_out[86]
port 386 nsew signal output
rlabel metal2 s 418986 0 419042 800 6 la_data_out[87]
port 387 nsew signal output
rlabel metal2 s 422390 0 422446 800 6 la_data_out[88]
port 388 nsew signal output
rlabel metal2 s 425794 0 425850 800 6 la_data_out[89]
port 389 nsew signal output
rlabel metal2 s 149518 0 149574 800 6 la_data_out[8]
port 390 nsew signal output
rlabel metal2 s 429198 0 429254 800 6 la_data_out[90]
port 391 nsew signal output
rlabel metal2 s 432602 0 432658 800 6 la_data_out[91]
port 392 nsew signal output
rlabel metal2 s 436006 0 436062 800 6 la_data_out[92]
port 393 nsew signal output
rlabel metal2 s 439410 0 439466 800 6 la_data_out[93]
port 394 nsew signal output
rlabel metal2 s 442814 0 442870 800 6 la_data_out[94]
port 395 nsew signal output
rlabel metal2 s 446218 0 446274 800 6 la_data_out[95]
port 396 nsew signal output
rlabel metal2 s 449622 0 449678 800 6 la_data_out[96]
port 397 nsew signal output
rlabel metal2 s 453026 0 453082 800 6 la_data_out[97]
port 398 nsew signal output
rlabel metal2 s 456430 0 456486 800 6 la_data_out[98]
port 399 nsew signal output
rlabel metal2 s 459834 0 459890 800 6 la_data_out[99]
port 400 nsew signal output
rlabel metal2 s 152922 0 152978 800 6 la_data_out[9]
port 401 nsew signal output
rlabel metal2 s 123298 0 123354 800 6 la_oen[0]
port 402 nsew signal input
rlabel metal2 s 464434 0 464490 800 6 la_oen[100]
port 403 nsew signal input
rlabel metal2 s 467838 0 467894 800 6 la_oen[101]
port 404 nsew signal input
rlabel metal2 s 471242 0 471298 800 6 la_oen[102]
port 405 nsew signal input
rlabel metal2 s 474646 0 474702 800 6 la_oen[103]
port 406 nsew signal input
rlabel metal2 s 478050 0 478106 800 6 la_oen[104]
port 407 nsew signal input
rlabel metal2 s 481454 0 481510 800 6 la_oen[105]
port 408 nsew signal input
rlabel metal2 s 484858 0 484914 800 6 la_oen[106]
port 409 nsew signal input
rlabel metal2 s 488262 0 488318 800 6 la_oen[107]
port 410 nsew signal input
rlabel metal2 s 491758 0 491814 800 6 la_oen[108]
port 411 nsew signal input
rlabel metal2 s 495162 0 495218 800 6 la_oen[109]
port 412 nsew signal input
rlabel metal2 s 157430 0 157486 800 6 la_oen[10]
port 413 nsew signal input
rlabel metal2 s 498566 0 498622 800 6 la_oen[110]
port 414 nsew signal input
rlabel metal2 s 501970 0 502026 800 6 la_oen[111]
port 415 nsew signal input
rlabel metal2 s 505374 0 505430 800 6 la_oen[112]
port 416 nsew signal input
rlabel metal2 s 508778 0 508834 800 6 la_oen[113]
port 417 nsew signal input
rlabel metal2 s 512182 0 512238 800 6 la_oen[114]
port 418 nsew signal input
rlabel metal2 s 515586 0 515642 800 6 la_oen[115]
port 419 nsew signal input
rlabel metal2 s 518990 0 519046 800 6 la_oen[116]
port 420 nsew signal input
rlabel metal2 s 522394 0 522450 800 6 la_oen[117]
port 421 nsew signal input
rlabel metal2 s 525798 0 525854 800 6 la_oen[118]
port 422 nsew signal input
rlabel metal2 s 529202 0 529258 800 6 la_oen[119]
port 423 nsew signal input
rlabel metal2 s 160834 0 160890 800 6 la_oen[11]
port 424 nsew signal input
rlabel metal2 s 532606 0 532662 800 6 la_oen[120]
port 425 nsew signal input
rlabel metal2 s 536102 0 536158 800 6 la_oen[121]
port 426 nsew signal input
rlabel metal2 s 539506 0 539562 800 6 la_oen[122]
port 427 nsew signal input
rlabel metal2 s 542910 0 542966 800 6 la_oen[123]
port 428 nsew signal input
rlabel metal2 s 546314 0 546370 800 6 la_oen[124]
port 429 nsew signal input
rlabel metal2 s 549718 0 549774 800 6 la_oen[125]
port 430 nsew signal input
rlabel metal2 s 553122 0 553178 800 6 la_oen[126]
port 431 nsew signal input
rlabel metal2 s 556526 0 556582 800 6 la_oen[127]
port 432 nsew signal input
rlabel metal2 s 164238 0 164294 800 6 la_oen[12]
port 433 nsew signal input
rlabel metal2 s 167642 0 167698 800 6 la_oen[13]
port 434 nsew signal input
rlabel metal2 s 171046 0 171102 800 6 la_oen[14]
port 435 nsew signal input
rlabel metal2 s 174450 0 174506 800 6 la_oen[15]
port 436 nsew signal input
rlabel metal2 s 177854 0 177910 800 6 la_oen[16]
port 437 nsew signal input
rlabel metal2 s 181350 0 181406 800 6 la_oen[17]
port 438 nsew signal input
rlabel metal2 s 184754 0 184810 800 6 la_oen[18]
port 439 nsew signal input
rlabel metal2 s 188158 0 188214 800 6 la_oen[19]
port 440 nsew signal input
rlabel metal2 s 126702 0 126758 800 6 la_oen[1]
port 441 nsew signal input
rlabel metal2 s 191562 0 191618 800 6 la_oen[20]
port 442 nsew signal input
rlabel metal2 s 194966 0 195022 800 6 la_oen[21]
port 443 nsew signal input
rlabel metal2 s 198370 0 198426 800 6 la_oen[22]
port 444 nsew signal input
rlabel metal2 s 201774 0 201830 800 6 la_oen[23]
port 445 nsew signal input
rlabel metal2 s 205178 0 205234 800 6 la_oen[24]
port 446 nsew signal input
rlabel metal2 s 208582 0 208638 800 6 la_oen[25]
port 447 nsew signal input
rlabel metal2 s 211986 0 212042 800 6 la_oen[26]
port 448 nsew signal input
rlabel metal2 s 215390 0 215446 800 6 la_oen[27]
port 449 nsew signal input
rlabel metal2 s 218794 0 218850 800 6 la_oen[28]
port 450 nsew signal input
rlabel metal2 s 222198 0 222254 800 6 la_oen[29]
port 451 nsew signal input
rlabel metal2 s 130106 0 130162 800 6 la_oen[2]
port 452 nsew signal input
rlabel metal2 s 225694 0 225750 800 6 la_oen[30]
port 453 nsew signal input
rlabel metal2 s 229098 0 229154 800 6 la_oen[31]
port 454 nsew signal input
rlabel metal2 s 232502 0 232558 800 6 la_oen[32]
port 455 nsew signal input
rlabel metal2 s 235906 0 235962 800 6 la_oen[33]
port 456 nsew signal input
rlabel metal2 s 239310 0 239366 800 6 la_oen[34]
port 457 nsew signal input
rlabel metal2 s 242714 0 242770 800 6 la_oen[35]
port 458 nsew signal input
rlabel metal2 s 246118 0 246174 800 6 la_oen[36]
port 459 nsew signal input
rlabel metal2 s 249522 0 249578 800 6 la_oen[37]
port 460 nsew signal input
rlabel metal2 s 252926 0 252982 800 6 la_oen[38]
port 461 nsew signal input
rlabel metal2 s 256330 0 256386 800 6 la_oen[39]
port 462 nsew signal input
rlabel metal2 s 133510 0 133566 800 6 la_oen[3]
port 463 nsew signal input
rlabel metal2 s 259734 0 259790 800 6 la_oen[40]
port 464 nsew signal input
rlabel metal2 s 263138 0 263194 800 6 la_oen[41]
port 465 nsew signal input
rlabel metal2 s 266542 0 266598 800 6 la_oen[42]
port 466 nsew signal input
rlabel metal2 s 270038 0 270094 800 6 la_oen[43]
port 467 nsew signal input
rlabel metal2 s 273442 0 273498 800 6 la_oen[44]
port 468 nsew signal input
rlabel metal2 s 276846 0 276902 800 6 la_oen[45]
port 469 nsew signal input
rlabel metal2 s 280250 0 280306 800 6 la_oen[46]
port 470 nsew signal input
rlabel metal2 s 283654 0 283710 800 6 la_oen[47]
port 471 nsew signal input
rlabel metal2 s 287058 0 287114 800 6 la_oen[48]
port 472 nsew signal input
rlabel metal2 s 290462 0 290518 800 6 la_oen[49]
port 473 nsew signal input
rlabel metal2 s 137006 0 137062 800 6 la_oen[4]
port 474 nsew signal input
rlabel metal2 s 293866 0 293922 800 6 la_oen[50]
port 475 nsew signal input
rlabel metal2 s 297270 0 297326 800 6 la_oen[51]
port 476 nsew signal input
rlabel metal2 s 300674 0 300730 800 6 la_oen[52]
port 477 nsew signal input
rlabel metal2 s 304078 0 304134 800 6 la_oen[53]
port 478 nsew signal input
rlabel metal2 s 307482 0 307538 800 6 la_oen[54]
port 479 nsew signal input
rlabel metal2 s 310886 0 310942 800 6 la_oen[55]
port 480 nsew signal input
rlabel metal2 s 314382 0 314438 800 6 la_oen[56]
port 481 nsew signal input
rlabel metal2 s 317786 0 317842 800 6 la_oen[57]
port 482 nsew signal input
rlabel metal2 s 321190 0 321246 800 6 la_oen[58]
port 483 nsew signal input
rlabel metal2 s 324594 0 324650 800 6 la_oen[59]
port 484 nsew signal input
rlabel metal2 s 140410 0 140466 800 6 la_oen[5]
port 485 nsew signal input
rlabel metal2 s 327998 0 328054 800 6 la_oen[60]
port 486 nsew signal input
rlabel metal2 s 331402 0 331458 800 6 la_oen[61]
port 487 nsew signal input
rlabel metal2 s 334806 0 334862 800 6 la_oen[62]
port 488 nsew signal input
rlabel metal2 s 338210 0 338266 800 6 la_oen[63]
port 489 nsew signal input
rlabel metal2 s 341614 0 341670 800 6 la_oen[64]
port 490 nsew signal input
rlabel metal2 s 345018 0 345074 800 6 la_oen[65]
port 491 nsew signal input
rlabel metal2 s 348422 0 348478 800 6 la_oen[66]
port 492 nsew signal input
rlabel metal2 s 351826 0 351882 800 6 la_oen[67]
port 493 nsew signal input
rlabel metal2 s 355230 0 355286 800 6 la_oen[68]
port 494 nsew signal input
rlabel metal2 s 358726 0 358782 800 6 la_oen[69]
port 495 nsew signal input
rlabel metal2 s 143814 0 143870 800 6 la_oen[6]
port 496 nsew signal input
rlabel metal2 s 362130 0 362186 800 6 la_oen[70]
port 497 nsew signal input
rlabel metal2 s 365534 0 365590 800 6 la_oen[71]
port 498 nsew signal input
rlabel metal2 s 368938 0 368994 800 6 la_oen[72]
port 499 nsew signal input
rlabel metal2 s 372342 0 372398 800 6 la_oen[73]
port 500 nsew signal input
rlabel metal2 s 375746 0 375802 800 6 la_oen[74]
port 501 nsew signal input
rlabel metal2 s 379150 0 379206 800 6 la_oen[75]
port 502 nsew signal input
rlabel metal2 s 382554 0 382610 800 6 la_oen[76]
port 503 nsew signal input
rlabel metal2 s 385958 0 386014 800 6 la_oen[77]
port 504 nsew signal input
rlabel metal2 s 389362 0 389418 800 6 la_oen[78]
port 505 nsew signal input
rlabel metal2 s 392766 0 392822 800 6 la_oen[79]
port 506 nsew signal input
rlabel metal2 s 147218 0 147274 800 6 la_oen[7]
port 507 nsew signal input
rlabel metal2 s 396170 0 396226 800 6 la_oen[80]
port 508 nsew signal input
rlabel metal2 s 399574 0 399630 800 6 la_oen[81]
port 509 nsew signal input
rlabel metal2 s 403070 0 403126 800 6 la_oen[82]
port 510 nsew signal input
rlabel metal2 s 406474 0 406530 800 6 la_oen[83]
port 511 nsew signal input
rlabel metal2 s 409878 0 409934 800 6 la_oen[84]
port 512 nsew signal input
rlabel metal2 s 413282 0 413338 800 6 la_oen[85]
port 513 nsew signal input
rlabel metal2 s 416686 0 416742 800 6 la_oen[86]
port 514 nsew signal input
rlabel metal2 s 420090 0 420146 800 6 la_oen[87]
port 515 nsew signal input
rlabel metal2 s 423494 0 423550 800 6 la_oen[88]
port 516 nsew signal input
rlabel metal2 s 426898 0 426954 800 6 la_oen[89]
port 517 nsew signal input
rlabel metal2 s 150622 0 150678 800 6 la_oen[8]
port 518 nsew signal input
rlabel metal2 s 430302 0 430358 800 6 la_oen[90]
port 519 nsew signal input
rlabel metal2 s 433706 0 433762 800 6 la_oen[91]
port 520 nsew signal input
rlabel metal2 s 437110 0 437166 800 6 la_oen[92]
port 521 nsew signal input
rlabel metal2 s 440514 0 440570 800 6 la_oen[93]
port 522 nsew signal input
rlabel metal2 s 443918 0 443974 800 6 la_oen[94]
port 523 nsew signal input
rlabel metal2 s 447414 0 447470 800 6 la_oen[95]
port 524 nsew signal input
rlabel metal2 s 450818 0 450874 800 6 la_oen[96]
port 525 nsew signal input
rlabel metal2 s 454222 0 454278 800 6 la_oen[97]
port 526 nsew signal input
rlabel metal2 s 457626 0 457682 800 6 la_oen[98]
port 527 nsew signal input
rlabel metal2 s 461030 0 461086 800 6 la_oen[99]
port 528 nsew signal input
rlabel metal2 s 154026 0 154082 800 6 la_oen[9]
port 529 nsew signal input
rlabel metal2 s 557630 0 557686 800 6 user_clock2
port 530 nsew signal input
rlabel metal2 s 570 0 626 800 6 wb_clk_i
port 531 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wb_rst_i
port 532 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 wbs_ack_o
port 533 nsew signal output
rlabel metal2 s 7378 0 7434 800 6 wbs_adr_i[0]
port 534 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 wbs_adr_i[10]
port 535 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 wbs_adr_i[11]
port 536 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 wbs_adr_i[12]
port 537 nsew signal input
rlabel metal2 s 56230 0 56286 800 6 wbs_adr_i[13]
port 538 nsew signal input
rlabel metal2 s 59634 0 59690 800 6 wbs_adr_i[14]
port 539 nsew signal input
rlabel metal2 s 63038 0 63094 800 6 wbs_adr_i[15]
port 540 nsew signal input
rlabel metal2 s 66442 0 66498 800 6 wbs_adr_i[16]
port 541 nsew signal input
rlabel metal2 s 69846 0 69902 800 6 wbs_adr_i[17]
port 542 nsew signal input
rlabel metal2 s 73250 0 73306 800 6 wbs_adr_i[18]
port 543 nsew signal input
rlabel metal2 s 76746 0 76802 800 6 wbs_adr_i[19]
port 544 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 wbs_adr_i[1]
port 545 nsew signal input
rlabel metal2 s 80150 0 80206 800 6 wbs_adr_i[20]
port 546 nsew signal input
rlabel metal2 s 83554 0 83610 800 6 wbs_adr_i[21]
port 547 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 wbs_adr_i[22]
port 548 nsew signal input
rlabel metal2 s 90362 0 90418 800 6 wbs_adr_i[23]
port 549 nsew signal input
rlabel metal2 s 93766 0 93822 800 6 wbs_adr_i[24]
port 550 nsew signal input
rlabel metal2 s 97170 0 97226 800 6 wbs_adr_i[25]
port 551 nsew signal input
rlabel metal2 s 100574 0 100630 800 6 wbs_adr_i[26]
port 552 nsew signal input
rlabel metal2 s 103978 0 104034 800 6 wbs_adr_i[27]
port 553 nsew signal input
rlabel metal2 s 107382 0 107438 800 6 wbs_adr_i[28]
port 554 nsew signal input
rlabel metal2 s 110786 0 110842 800 6 wbs_adr_i[29]
port 555 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 wbs_adr_i[2]
port 556 nsew signal input
rlabel metal2 s 114190 0 114246 800 6 wbs_adr_i[30]
port 557 nsew signal input
rlabel metal2 s 117594 0 117650 800 6 wbs_adr_i[31]
port 558 nsew signal input
rlabel metal2 s 20994 0 21050 800 6 wbs_adr_i[3]
port 559 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 wbs_adr_i[4]
port 560 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 wbs_adr_i[5]
port 561 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 wbs_adr_i[6]
port 562 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 wbs_adr_i[7]
port 563 nsew signal input
rlabel metal2 s 39210 0 39266 800 6 wbs_adr_i[8]
port 564 nsew signal input
rlabel metal2 s 42614 0 42670 800 6 wbs_adr_i[9]
port 565 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 wbs_cyc_i
port 566 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_dat_i[0]
port 567 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 wbs_dat_i[10]
port 568 nsew signal input
rlabel metal2 s 50526 0 50582 800 6 wbs_dat_i[11]
port 569 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 wbs_dat_i[12]
port 570 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 wbs_dat_i[13]
port 571 nsew signal input
rlabel metal2 s 60830 0 60886 800 6 wbs_dat_i[14]
port 572 nsew signal input
rlabel metal2 s 64234 0 64290 800 6 wbs_dat_i[15]
port 573 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 wbs_dat_i[16]
port 574 nsew signal input
rlabel metal2 s 71042 0 71098 800 6 wbs_dat_i[17]
port 575 nsew signal input
rlabel metal2 s 74446 0 74502 800 6 wbs_dat_i[18]
port 576 nsew signal input
rlabel metal2 s 77850 0 77906 800 6 wbs_dat_i[19]
port 577 nsew signal input
rlabel metal2 s 12990 0 13046 800 6 wbs_dat_i[1]
port 578 nsew signal input
rlabel metal2 s 81254 0 81310 800 6 wbs_dat_i[20]
port 579 nsew signal input
rlabel metal2 s 84658 0 84714 800 6 wbs_dat_i[21]
port 580 nsew signal input
rlabel metal2 s 88062 0 88118 800 6 wbs_dat_i[22]
port 581 nsew signal input
rlabel metal2 s 91466 0 91522 800 6 wbs_dat_i[23]
port 582 nsew signal input
rlabel metal2 s 94870 0 94926 800 6 wbs_dat_i[24]
port 583 nsew signal input
rlabel metal2 s 98274 0 98330 800 6 wbs_dat_i[25]
port 584 nsew signal input
rlabel metal2 s 101678 0 101734 800 6 wbs_dat_i[26]
port 585 nsew signal input
rlabel metal2 s 105174 0 105230 800 6 wbs_dat_i[27]
port 586 nsew signal input
rlabel metal2 s 108578 0 108634 800 6 wbs_dat_i[28]
port 587 nsew signal input
rlabel metal2 s 111982 0 112038 800 6 wbs_dat_i[29]
port 588 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 wbs_dat_i[2]
port 589 nsew signal input
rlabel metal2 s 115386 0 115442 800 6 wbs_dat_i[30]
port 590 nsew signal input
rlabel metal2 s 118790 0 118846 800 6 wbs_dat_i[31]
port 591 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 wbs_dat_i[3]
port 592 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 wbs_dat_i[4]
port 593 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 wbs_dat_i[5]
port 594 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 wbs_dat_i[6]
port 595 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 wbs_dat_i[7]
port 596 nsew signal input
rlabel metal2 s 40314 0 40370 800 6 wbs_dat_i[8]
port 597 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 wbs_dat_i[9]
port 598 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_dat_o[0]
port 599 nsew signal output
rlabel metal2 s 48318 0 48374 800 6 wbs_dat_o[10]
port 600 nsew signal output
rlabel metal2 s 51722 0 51778 800 6 wbs_dat_o[11]
port 601 nsew signal output
rlabel metal2 s 55126 0 55182 800 6 wbs_dat_o[12]
port 602 nsew signal output
rlabel metal2 s 58530 0 58586 800 6 wbs_dat_o[13]
port 603 nsew signal output
rlabel metal2 s 61934 0 61990 800 6 wbs_dat_o[14]
port 604 nsew signal output
rlabel metal2 s 65338 0 65394 800 6 wbs_dat_o[15]
port 605 nsew signal output
rlabel metal2 s 68742 0 68798 800 6 wbs_dat_o[16]
port 606 nsew signal output
rlabel metal2 s 72146 0 72202 800 6 wbs_dat_o[17]
port 607 nsew signal output
rlabel metal2 s 75550 0 75606 800 6 wbs_dat_o[18]
port 608 nsew signal output
rlabel metal2 s 78954 0 79010 800 6 wbs_dat_o[19]
port 609 nsew signal output
rlabel metal2 s 14186 0 14242 800 6 wbs_dat_o[1]
port 610 nsew signal output
rlabel metal2 s 82358 0 82414 800 6 wbs_dat_o[20]
port 611 nsew signal output
rlabel metal2 s 85762 0 85818 800 6 wbs_dat_o[21]
port 612 nsew signal output
rlabel metal2 s 89166 0 89222 800 6 wbs_dat_o[22]
port 613 nsew signal output
rlabel metal2 s 92662 0 92718 800 6 wbs_dat_o[23]
port 614 nsew signal output
rlabel metal2 s 96066 0 96122 800 6 wbs_dat_o[24]
port 615 nsew signal output
rlabel metal2 s 99470 0 99526 800 6 wbs_dat_o[25]
port 616 nsew signal output
rlabel metal2 s 102874 0 102930 800 6 wbs_dat_o[26]
port 617 nsew signal output
rlabel metal2 s 106278 0 106334 800 6 wbs_dat_o[27]
port 618 nsew signal output
rlabel metal2 s 109682 0 109738 800 6 wbs_dat_o[28]
port 619 nsew signal output
rlabel metal2 s 113086 0 113142 800 6 wbs_dat_o[29]
port 620 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 wbs_dat_o[2]
port 621 nsew signal output
rlabel metal2 s 116490 0 116546 800 6 wbs_dat_o[30]
port 622 nsew signal output
rlabel metal2 s 119894 0 119950 800 6 wbs_dat_o[31]
port 623 nsew signal output
rlabel metal2 s 23294 0 23350 800 6 wbs_dat_o[3]
port 624 nsew signal output
rlabel metal2 s 27802 0 27858 800 6 wbs_dat_o[4]
port 625 nsew signal output
rlabel metal2 s 31206 0 31262 800 6 wbs_dat_o[5]
port 626 nsew signal output
rlabel metal2 s 34610 0 34666 800 6 wbs_dat_o[6]
port 627 nsew signal output
rlabel metal2 s 38014 0 38070 800 6 wbs_dat_o[7]
port 628 nsew signal output
rlabel metal2 s 41418 0 41474 800 6 wbs_dat_o[8]
port 629 nsew signal output
rlabel metal2 s 44822 0 44878 800 6 wbs_dat_o[9]
port 630 nsew signal output
rlabel metal2 s 10782 0 10838 800 6 wbs_sel_i[0]
port 631 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 wbs_sel_i[1]
port 632 nsew signal input
rlabel metal2 s 19890 0 19946 800 6 wbs_sel_i[2]
port 633 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 wbs_sel_i[3]
port 634 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 wbs_stb_i
port 635 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wbs_we_i
port 636 nsew signal input
rlabel metal4 s 557168 2128 557488 681680 6 VPWR
port 637 nsew power bidirectional
rlabel metal4 s 526448 2128 526768 681680 6 VPWR
port 638 nsew power bidirectional
rlabel metal4 s 495728 2128 496048 681680 6 VPWR
port 639 nsew power bidirectional
rlabel metal4 s 465008 2128 465328 681680 6 VPWR
port 640 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 681680 6 VPWR
port 641 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 681680 6 VPWR
port 642 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 681680 6 VPWR
port 643 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 681680 6 VPWR
port 644 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 681680 6 VPWR
port 645 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 681680 6 VPWR
port 646 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 681680 6 VPWR
port 647 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 681680 6 VPWR
port 648 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 681680 6 VPWR
port 649 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 681680 6 VPWR
port 650 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 681680 6 VPWR
port 651 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 681680 6 VPWR
port 652 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 681680 6 VPWR
port 653 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 681680 6 VPWR
port 654 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 681680 6 VPWR
port 655 nsew power bidirectional
rlabel metal4 s 541808 2128 542128 681680 6 VGND
port 656 nsew ground bidirectional
rlabel metal4 s 511088 2128 511408 681680 6 VGND
port 657 nsew ground bidirectional
rlabel metal4 s 480368 2128 480688 681680 6 VGND
port 658 nsew ground bidirectional
rlabel metal4 s 449648 2128 449968 681680 6 VGND
port 659 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 681680 6 VGND
port 660 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 681680 6 VGND
port 661 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 681680 6 VGND
port 662 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 681680 6 VGND
port 663 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 681680 6 VGND
port 664 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 681680 6 VGND
port 665 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 681680 6 VGND
port 666 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 681680 6 VGND
port 667 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 681680 6 VGND
port 668 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 681680 6 VGND
port 669 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 681680 6 VGND
port 670 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 681680 6 VGND
port 671 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 681680 6 VGND
port 672 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 681680 6 VGND
port 673 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 564000 684000
string LEFview TRUE
<< end >>
